* NGSPICE file created from Motor_Top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

.subckt Motor_Top clock io_ba_match io_motor_irq io_pwm_high io_pwm_low io_qei_ch_a
+ io_qei_ch_b io_wbs_ack_o io_wbs_data_o[0] io_wbs_data_o[10] io_wbs_data_o[11] io_wbs_data_o[12]
+ io_wbs_data_o[13] io_wbs_data_o[14] io_wbs_data_o[15] io_wbs_data_o[16] io_wbs_data_o[17]
+ io_wbs_data_o[18] io_wbs_data_o[19] io_wbs_data_o[1] io_wbs_data_o[20] io_wbs_data_o[21]
+ io_wbs_data_o[22] io_wbs_data_o[23] io_wbs_data_o[24] io_wbs_data_o[25] io_wbs_data_o[26]
+ io_wbs_data_o[27] io_wbs_data_o[28] io_wbs_data_o[29] io_wbs_data_o[2] io_wbs_data_o[30]
+ io_wbs_data_o[31] io_wbs_data_o[3] io_wbs_data_o[4] io_wbs_data_o[5] io_wbs_data_o[6]
+ io_wbs_data_o[7] io_wbs_data_o[8] io_wbs_data_o[9] io_wbs_m2s_addr[0] io_wbs_m2s_addr[10]
+ io_wbs_m2s_addr[11] io_wbs_m2s_addr[12] io_wbs_m2s_addr[13] io_wbs_m2s_addr[14]
+ io_wbs_m2s_addr[15] io_wbs_m2s_addr[1] io_wbs_m2s_addr[2] io_wbs_m2s_addr[3] io_wbs_m2s_addr[4]
+ io_wbs_m2s_addr[5] io_wbs_m2s_addr[6] io_wbs_m2s_addr[7] io_wbs_m2s_addr[8] io_wbs_m2s_addr[9]
+ io_wbs_m2s_data[0] io_wbs_m2s_data[10] io_wbs_m2s_data[11] io_wbs_m2s_data[12] io_wbs_m2s_data[13]
+ io_wbs_m2s_data[14] io_wbs_m2s_data[15] io_wbs_m2s_data[16] io_wbs_m2s_data[17]
+ io_wbs_m2s_data[18] io_wbs_m2s_data[19] io_wbs_m2s_data[1] io_wbs_m2s_data[20] io_wbs_m2s_data[21]
+ io_wbs_m2s_data[22] io_wbs_m2s_data[23] io_wbs_m2s_data[24] io_wbs_m2s_data[25]
+ io_wbs_m2s_data[26] io_wbs_m2s_data[27] io_wbs_m2s_data[28] io_wbs_m2s_data[29]
+ io_wbs_m2s_data[2] io_wbs_m2s_data[30] io_wbs_m2s_data[31] io_wbs_m2s_data[3] io_wbs_m2s_data[4]
+ io_wbs_m2s_data[5] io_wbs_m2s_data[6] io_wbs_m2s_data[7] io_wbs_m2s_data[8] io_wbs_m2s_data[9]
+ io_wbs_m2s_sel[0] io_wbs_m2s_sel[1] io_wbs_m2s_sel[2] io_wbs_m2s_sel[3] io_wbs_m2s_stb
+ io_wbs_m2s_we reset vccd1 vssd1
X_05903_ _06038_/A _05906_/A vssd1 vssd1 vccd1 vccd1 _05904_/B sky130_fd_sc_hd__and2_1
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08731__B1 _08676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__nand2_1
X_06883_ _06883_/A _06883_/B vssd1 vssd1 vccd1 vccd1 _06884_/B sky130_fd_sc_hd__nor2_1
X_05834_ _05834_/A _05844_/C vssd1 vssd1 vccd1 vccd1 _05838_/B sky130_fd_sc_hd__or2_1
XFILLER_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08622_ _10790_/Q _08617_/X _08621_/Y vssd1 vssd1 vccd1 vccd1 _10790_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05765_ _05750_/X _05765_/B _05765_/C _05765_/D vssd1 vssd1 vccd1 vccd1 _05787_/A
+ sky130_fd_sc_hd__and4b_1
X_08553_ _10771_/Q _08553_/B vssd1 vssd1 vccd1 vccd1 _08554_/B sky130_fd_sc_hd__xor2_1
XFILLER_70_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08484_ _08484_/A vssd1 vssd1 vccd1 vccd1 _10744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07504_ _07504_/A _07504_/B _07535_/A vssd1 vssd1 vccd1 vccd1 _07505_/B sky130_fd_sc_hd__or3_1
X_05696_ _08173_/A _10552_/Q _05694_/Y _08160_/A vssd1 vssd1 vccd1 vccd1 _05798_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07435_ _07727_/A _07713_/A _07728_/B _07729_/B vssd1 vssd1 vccd1 vccd1 _07714_/S
+ sky130_fd_sc_hd__nand4_1
XFILLER_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07366_ _07366_/A _07366_/B _07366_/C vssd1 vssd1 vccd1 vccd1 _07367_/B sky130_fd_sc_hd__and3_1
X_09105_ _05462_/A _09148_/A _07969_/A _09104_/Y vssd1 vssd1 vccd1 vccd1 _09105_/X
+ sky130_fd_sc_hd__o211a_1
X_06317_ _06317_/A _06317_/B vssd1 vssd1 vccd1 vccd1 _06729_/A sky130_fd_sc_hd__nand2_1
X_07297_ _07310_/A _07297_/B vssd1 vssd1 vccd1 vccd1 _07298_/C sky130_fd_sc_hd__xnor2_1
X_06248_ input36/X _06238_/X _06246_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10612_/D
+ sky130_fd_sc_hd__o211a_1
X_09036_ _09209_/B vssd1 vssd1 vccd1 vccd1 _09036_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06179_ _10593_/Q vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__inv_2
XANTENNA__10357__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09275__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09938_ _10482_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _09940_/B sky130_fd_sc_hd__nand2_1
XFILLER_131_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05308__A _10671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09869_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__o21ai_2
XFILLER_46_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09214__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _10737_/CLK _10713_/D vssd1 vssd1 vccd1 vccd1 _10713_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08238__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10644_ _10646_/CLK _10644_/D vssd1 vssd1 vccd1 vccd1 _10644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10575_ _10833_/CLK _10575_/D vssd1 vssd1 vccd1 vccd1 _10575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_23_clock_A _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10009_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__and3_1
XANTENNA__10520__B1 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05550_ _10548_/Q _05629_/B vssd1 vssd1 vccd1 vccd1 _05630_/A sky130_fd_sc_hd__or2_1
XFILLER_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05481_ _05912_/B _05470_/B _05495_/A _08994_/A _05480_/Y vssd1 vssd1 vccd1 vccd1
+ _10542_/D sky130_fd_sc_hd__a221o_1
XFILLER_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05888__A _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07220_ _07102_/A _07215_/B _07249_/B _07248_/A vssd1 vssd1 vccd1 vccd1 _07242_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07151_ _07151_/A _07394_/A _07151_/C vssd1 vssd1 vccd1 vccd1 _07322_/A sky130_fd_sc_hd__and3_1
X_06102_ _10695_/Q _08208_/B vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__or2_1
X_07082_ _09356_/A _07060_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _07083_/B sky130_fd_sc_hd__o21ai_1
X_06033_ _08096_/A vssd1 vssd1 vccd1 vccd1 _06033_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_126_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10339__B1 _07539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07984_ _08015_/A vssd1 vssd1 vccd1 vccd1 _07985_/B sky130_fd_sc_hd__buf_4
XFILLER_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09723_ _09723_/A _09723_/B _09723_/C vssd1 vssd1 vccd1 vccd1 _09723_/Y sky130_fd_sc_hd__nand3_1
X_06935_ _06935_/A _06935_/B vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__xnor2_4
XFILLER_83_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06866_ _06867_/B _06866_/B vssd1 vssd1 vccd1 vccd1 _06868_/A sky130_fd_sc_hd__and2b_1
X_09654_ _09867_/A _09717_/A vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05817_ _06065_/A _09078_/A _05816_/X vssd1 vssd1 vccd1 vccd1 _05909_/A sky130_fd_sc_hd__o21a_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08439__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _08498_/X _08617_/B _08604_/Y _08630_/A vssd1 vssd1 vccd1 vccd1 _10785_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09585_ _10968_/Q _09642_/A _09492_/A _10967_/Q vssd1 vssd1 vccd1 vccd1 _09587_/A
+ sky130_fd_sc_hd__a22o_1
X_06797_ _06882_/A _06836_/A vssd1 vssd1 vccd1 vccd1 _06823_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05748_ _10703_/Q vssd1 vssd1 vccd1 vccd1 _05749_/A sky130_fd_sc_hd__inv_2
X_08536_ _08624_/B vssd1 vssd1 vccd1 vccd1 _08686_/A sky130_fd_sc_hd__clkbuf_4
X_05679_ _08304_/A _05580_/X _05583_/Y _05803_/A _05678_/X vssd1 vssd1 vccd1 vccd1
+ _05679_/X sky130_fd_sc_hd__o221a_1
X_08467_ _08572_/B _10739_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08398_ _10198_/A vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__clkbuf_1
X_07418_ _07732_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07349_ _07349_/A _07349_/B _07349_/C vssd1 vssd1 vccd1 vccd1 _07350_/B sky130_fd_sc_hd__nor3_1
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10360_ _08491_/X _06818_/A _10355_/X _10927_/Q vssd1 vssd1 vccd1 vccd1 _10927_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07994__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ _08998_/X _09001_/X _09018_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10835_/D
+ sky130_fd_sc_hd__o31a_2
X_10291_ _10289_/X _10300_/B _10291_/S vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05964__C input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08349__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07700__B _07700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08226__A2 _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06237__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10627_ _10806_/CLK _10627_/D vssd1 vssd1 vccd1 vccd1 _10627_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10558_ _10700_/CLK _10558_/D vssd1 vssd1 vccd1 vccd1 _10558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08531__B _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10489_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06720_ _06720_/A _06720_/B vssd1 vssd1 vccd1 vccd1 _06725_/A sky130_fd_sc_hd__xnor2_1
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07163__A _07415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06651_ _06648_/A _06648_/B _06654_/A vssd1 vssd1 vccd1 vccd1 _06652_/B sky130_fd_sc_hd__o21ba_1
XFILLER_37_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05602_ _05602_/A _05602_/B vssd1 vssd1 vccd1 vccd1 _05602_/X sky130_fd_sc_hd__and2_1
XFILLER_92_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09370_ _09606_/B _09607_/A _09369_/X vssd1 vssd1 vccd1 vccd1 _09674_/B sky130_fd_sc_hd__a21oi_2
X_06582_ _06581_/B _06581_/C _06581_/A vssd1 vssd1 vccd1 vccd1 _06593_/B sky130_fd_sc_hd__o21ai_1
X_08321_ _08321_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08321_/X sky130_fd_sc_hd__or2_1
X_05533_ _10545_/Q vssd1 vssd1 vccd1 vccd1 _05547_/A sky130_fd_sc_hd__inv_2
XFILLER_33_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08252_ _08243_/A _08251_/C _05598_/X vssd1 vssd1 vccd1 vccd1 _08252_/Y sky130_fd_sc_hd__a21oi_1
X_05464_ _10647_/Q _10646_/Q _07922_/A _07919_/A vssd1 vssd1 vccd1 vccd1 _05467_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_60_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07610__B _07706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07203_ _07204_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07205_/A sky130_fd_sc_hd__or2_1
XFILLER_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _05883_/A _08043_/A _08179_/Y _08038_/A _08182_/Y vssd1 vssd1 vccd1 vccd1
+ _08185_/A sky130_fd_sc_hd__a221o_1
XFILLER_118_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05395_ _10576_/Q vssd1 vssd1 vccd1 vccd1 _05452_/A sky130_fd_sc_hd__inv_2
XANTENNA__06228__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07134_ _07134_/A _07134_/B vssd1 vssd1 vccd1 vccd1 _07295_/A sky130_fd_sc_hd__xnor2_1
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07065_ _09381_/A _07056_/A _07056_/B vssd1 vssd1 vccd1 vccd1 _07066_/B sky130_fd_sc_hd__a21oi_1
X_06016_ input8/X _08048_/A vssd1 vssd1 vccd1 vccd1 _09098_/A sky130_fd_sc_hd__or2_1
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07967_ _07967_/A _09013_/A vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__nor2_1
XFILLER_75_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09706_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__nand2_1
X_06918_ _10515_/A _07682_/B _06918_/C vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__and3_1
XANTENNA__08153__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08153__A1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _07898_/A _07898_/B vssd1 vssd1 vccd1 vccd1 _10638_/D sky130_fd_sc_hd__nor2_1
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09637_ _09834_/B _09692_/A vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__and2_2
X_06849_ _06900_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _06860_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10849__D _10849_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _09568_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__or2b_1
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08519_ _10797_/Q _08514_/X _08517_/X hold21/A vssd1 vssd1 vccd1 vccd1 _10760_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _09542_/B _09499_/B _09499_/C vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__nand3_1
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06219__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10412_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10343_ _10343_/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__and2_1
XANTENNA__09447__B _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05978__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06152__A _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ _10956_/Q _10940_/Q vssd1 vssd1 vccd1 vccd1 _10287_/C sky130_fd_sc_hd__or2b_1
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05991__A _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10254__A2 _10253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ _08844_/A _08870_/B _08870_/C _08870_/D vssd1 vssd1 vccd1 vccd1 _08871_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_69_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06997__A _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07821_ _06151_/A _06258_/X _07807_/X _07820_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07821_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_57_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07752_ _07586_/A _07586_/B _07751_/X vssd1 vssd1 vccd1 vccd1 _07753_/B sky130_fd_sc_hd__o21ai_1
XFILLER_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06703_ _06893_/A _06893_/B _06702_/X vssd1 vssd1 vccd1 vccd1 _06885_/B sky130_fd_sc_hd__a21o_2
X_07683_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__and2_1
XFILLER_92_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06634_ _06634_/A _06634_/B vssd1 vssd1 vccd1 vccd1 _06635_/B sky130_fd_sc_hd__nand2_1
X_09422_ _09422_/A _09422_/B vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__xnor2_1
XFILLER_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09353_ _09371_/B _09353_/B vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__or2_1
X_08304_ _08304_/A vssd1 vssd1 vccd1 vccd1 _08305_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06565_ _06564_/A _06564_/B _06584_/A vssd1 vssd1 vccd1 vccd1 _06571_/A sky130_fd_sc_hd__o21ai_1
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05516_ _05337_/B _05510_/X _05513_/X _07903_/A vssd1 vssd1 vccd1 vccd1 _10565_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09284_ _09289_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__and2_1
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06496_ _06496_/A vssd1 vssd1 vccd1 vccd1 _06521_/A sky130_fd_sc_hd__clkbuf_2
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08235_/Y sky130_fd_sc_hd__nor2_1
X_05447_ _07922_/A _05324_/X _05318_/X _07925_/A _05446_/X vssd1 vssd1 vccd1 vccd1
+ _05447_/X sky130_fd_sc_hd__o221a_1
XFILLER_119_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08166_ _08166_/A vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__buf_4
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05378_ _10658_/Q _05380_/A vssd1 vssd1 vccd1 vccd1 _05378_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07117_ _10984_/Q _07125_/A _07222_/B _10983_/Q vssd1 vssd1 vccd1 vccd1 _07117_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ _08092_/X _08094_/X _08105_/B _08096_/X vssd1 vssd1 vccd1 vccd1 _08097_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_106_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07048_ _07048_/A _07048_/B vssd1 vssd1 vccd1 vccd1 _07463_/B sky130_fd_sc_hd__xnor2_1
XFILLER_130_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08999_ _09079_/A vssd1 vssd1 vccd1 vccd1 _08999_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08126__A1 _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05316__A _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10961_ _10962_/CLK _10961_/D vssd1 vssd1 vccd1 vccd1 _10961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10892_ _10909_/CLK _10892_/D vssd1 vssd1 vccd1 vccd1 _10892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06147__A _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10814_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__05986__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10326_ _10325_/X _10318_/Y _10316_/B vssd1 vssd1 vccd1 vccd1 _10327_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10257_ _10257_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_66_clock _10981_/CLK vssd1 vssd1 vccd1 vccd1 _10920_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10188_ _07539_/A _10043_/A _10184_/X _10897_/Q vssd1 vssd1 vccd1 vccd1 _10897_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06350_ _06457_/A vssd1 vssd1 vccd1 vccd1 _06895_/A sky130_fd_sc_hd__clkbuf_2
X_05301_ _07991_/A _05369_/A vssd1 vssd1 vccd1 vccd1 _05362_/B sky130_fd_sc_hd__nand2_1
X_06281_ _06338_/A _06281_/B vssd1 vssd1 vccd1 vccd1 _06352_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_clock _10857_/CLK vssd1 vssd1 vccd1 vccd1 _10682_/CLK sky130_fd_sc_hd__clkbuf_16
X_08020_ input32/X _08015_/X _08018_/Y _08019_/X vssd1 vssd1 vccd1 vccd1 _10672_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_71_clock_A _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ _09971_/A vssd1 vssd1 vccd1 vccd1 _09971_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _08927_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07159__A2 _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08853_ input29/X _08785_/X _08786_/X _10820_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08853_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08108__A1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08784_ _08773_/A _08778_/B _08803_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _08784_/X
+ sky130_fd_sc_hd__a31o_1
X_05996_ _08201_/A vssd1 vssd1 vccd1 vccd1 _09403_/A sky130_fd_sc_hd__buf_4
XFILLER_57_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07804_ _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _07804_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08108__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07735_ _07735_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09405_ _09757_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09405_/X sky130_fd_sc_hd__or2_1
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06617_ _06672_/A _06672_/B _06616_/Y vssd1 vssd1 vccd1 vccd1 _06668_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07597_ _07751_/A _07597_/B vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__xor2_4
X_06548_ _06567_/A _06547_/C _06567_/B _06568_/A vssd1 vssd1 vccd1 vccd1 _06549_/B
+ sky130_fd_sc_hd__a22oi_1
X_09336_ _09336_/A _09336_/B vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__xor2_4
XFILLER_138_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08292__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _09267_/A vssd1 vssd1 vccd1 vccd1 _10859_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_138_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08218_ _08218_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08228_/B sky130_fd_sc_hd__nor2_1
X_06479_ _06479_/A _06479_/B vssd1 vssd1 vccd1 vccd1 _06480_/B sky130_fd_sc_hd__and2_1
XFILLER_119_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09198_ _07871_/A _09136_/A _09148_/A _08208_/A _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09198_/X sky130_fd_sc_hd__a221o_1
X_08149_ _08169_/C vssd1 vssd1 vccd1 vccd1 _08149_/Y sky130_fd_sc_hd__inv_2
XFILLER_119_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10862__D _10862_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08910__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10111_ _10039_/Y _10042_/B _10040_/A vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10042_ _10042_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10042_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_130_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input18_A io_wbs_m2s_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08357__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ _10945_/CLK _10944_/D vssd1 vssd1 vccd1 vccd1 _10944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10875_ _10909_/CLK _10875_/D vssd1 vssd1 vccd1 vccd1 _10875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08283__B1 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08820__A _08820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10309_ _10309_/A vssd1 vssd1 vccd1 vccd1 _10309_/Y sky130_fd_sc_hd__inv_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08338__A1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05850_ _10668_/Q _05863_/B vssd1 vssd1 vccd1 vccd1 _05857_/B sky130_fd_sc_hd__or2_1
XFILLER_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05781_ _08315_/B vssd1 vssd1 vccd1 vccd1 _05781_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_18_clock_A _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07520_ _07661_/A _07668_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__or3_1
XFILLER_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07451_ _07598_/A _07451_/B vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07382_ _07382_/A vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__clkinv_2
X_06402_ _06441_/B _06409_/B vssd1 vssd1 vccd1 vccd1 _06690_/A sky130_fd_sc_hd__and2_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09121_ _10518_/B vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__clkbuf_2
X_06333_ _06371_/B _06371_/C _06804_/A vssd1 vssd1 vccd1 vccd1 _06334_/B sky130_fd_sc_hd__o21a_1
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09052_ _10716_/Q _08999_/X _09037_/Y _08701_/A vssd1 vssd1 vccd1 vccd1 _09052_/X
+ sky130_fd_sc_hd__a22o_1
X_06264_ _10917_/Q _10900_/Q vssd1 vssd1 vccd1 vccd1 _06270_/A sky130_fd_sc_hd__nand2_1
XFILLER_116_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08003_ _08235_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__or2_1
X_06195_ input20/X vssd1 vssd1 vccd1 vccd1 _06195_/X sky130_fd_sc_hd__buf_4
XFILLER_104_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10384__A1 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _09953_/Y _09878_/B _09882_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09955_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_131_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08905_ _10826_/Q _10825_/Q _10824_/Q _08876_/A _08902_/B vssd1 vssd1 vccd1 vccd1
+ _08905_/X sky130_fd_sc_hd__o41a_1
XANTENNA__10136__A1 _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _09883_/Y _09809_/B _09884_/X vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__o21ba_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08825_/A _08828_/Y _08841_/C _08688_/A vssd1 vssd1 vccd1 vccd1 _08836_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05979_ _05958_/X _05975_/X _05978_/Y vssd1 vssd1 vccd1 vccd1 _10573_/D sky130_fd_sc_hd__o21a_1
X_08767_ _08758_/A _08761_/Y _08804_/C _08688_/A vssd1 vssd1 vccd1 vccd1 _08767_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08698_ _08698_/A vssd1 vssd1 vccd1 vccd1 _08732_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10500__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07718_ _07718_/A vssd1 vssd1 vccd1 vccd1 _07718_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _07649_/A _07649_/B vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _10694_/CLK _10660_/D vssd1 vssd1 vccd1 vccd1 _10660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09319_ _09536_/B vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10591_ _10878_/CLK _10591_/D vssd1 vssd1 vccd1 vccd1 _10591_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08624__B _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05967__C input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput75 _10861_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[27] sky130_fd_sc_hd__buf_2
Xoutput53 _05956_/X vssd1 vssd1 vccd1 vccd1 io_pwm_high sky130_fd_sc_hd__buf_2
XFILLER_134_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput64 _10851_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput86 _10842_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10025_ _10097_/A _10025_/B vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08087__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10927_ _10930_/CLK _10927_/D vssd1 vssd1 vccd1 vccd1 _10927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06319__B _10907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10858_ _10862_/CLK _10858_/D vssd1 vssd1 vccd1 vccd1 _10858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10791_/CLK _10789_/D vssd1 vssd1 vccd1 vccd1 _10789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08550__A _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10291__S _10291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06951_ _06951_/A _06951_/B vssd1 vssd1 vccd1 vccd1 _06952_/B sky130_fd_sc_hd__and2_1
X_05902_ _08119_/A _05904_/A vssd1 vssd1 vccd1 vccd1 _05902_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09670_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09670_/Y sky130_fd_sc_hd__nor2_1
X_08621_ _10790_/Q _08617_/X _08630_/A vssd1 vssd1 vccd1 vccd1 _08621_/Y sky130_fd_sc_hd__a21oi_1
X_06882_ _06882_/A _06882_/B vssd1 vssd1 vccd1 vccd1 _06883_/B sky130_fd_sc_hd__and2_1
X_05833_ _10675_/Q vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__buf_2
XFILLER_55_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05764_ _05764_/A _05791_/A _05789_/A vssd1 vssd1 vccd1 vccd1 _05765_/D sky130_fd_sc_hd__and3_1
X_08552_ _08586_/A vssd1 vssd1 vccd1 vccd1 _08583_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ _08483_/A _08483_/B vssd1 vssd1 vccd1 vccd1 _08484_/A sky130_fd_sc_hd__and2_1
XANTENNA__08495__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07503_ _07503_/A vssd1 vssd1 vccd1 vccd1 _07606_/A sky130_fd_sc_hd__inv_2
XFILLER_35_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05695_ _08169_/B vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07434_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07729_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07365_ _07366_/A _07366_/B _07366_/C vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__a21oi_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09104_ _09104_/A _09104_/B vssd1 vssd1 vccd1 vccd1 _09104_/Y sky130_fd_sc_hd__nand2_1
X_06316_ _10925_/Q _10908_/Q vssd1 vssd1 vccd1 vccd1 _06317_/B sky130_fd_sc_hd__or2_1
X_07296_ _07296_/A _07296_/B vssd1 vssd1 vccd1 vccd1 _07297_/B sky130_fd_sc_hd__or2_1
X_06247_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06247_/X sky130_fd_sc_hd__clkbuf_4
X_09035_ _09037_/A _09035_/B _09211_/B vssd1 vssd1 vccd1 vccd1 _09209_/B sky130_fd_sc_hd__or3_2
XFILLER_117_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06178_ input47/X vssd1 vssd1 vccd1 vccd1 _06178_/X sky130_fd_sc_hd__buf_4
XFILLER_104_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08970__A1 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _09937_/A vssd1 vssd1 vccd1 vccd1 _10123_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_131_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09868_ _09868_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09870_/C sky130_fd_sc_hd__nor2_1
XFILLER_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08819_ _08819_/A vssd1 vssd1 vccd1 vccd1 _08819_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07804__A _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09799_ _09859_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09937_/A sky130_fd_sc_hd__xnor2_2
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10737_/CLK _10712_/D vssd1 vssd1 vccd1 vccd1 _10712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10643_ _10646_/CLK _10643_/D vssd1 vssd1 vccd1 vccd1 _10643_/Q sky130_fd_sc_hd__dfxtp_1
X_10574_ _10833_/CLK _10574_/D vssd1 vssd1 vccd1 vccd1 _10574_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05994__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08370__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__C1 _07393_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10405__A _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08961__B2 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__a21oi_1
XFILLER_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10140__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05480_ _05480_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _07150_/A _07150_/B vssd1 vssd1 vccd1 vccd1 _07151_/C sky130_fd_sc_hd__xnor2_1
X_06101_ _10694_/Q _10693_/Q _08191_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__or3_1
XFILLER_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _07149_/C vssd1 vssd1 vccd1 vccd1 _07326_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06032_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07983_ _07983_/A vssd1 vssd1 vccd1 vccd1 _08015_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09722_ _09723_/A _09723_/B _09723_/C vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__a21oi_1
XFILLER_86_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06934_ _06934_/A _06934_/B vssd1 vssd1 vccd1 vccd1 _06966_/A sky130_fd_sc_hd__xor2_4
XFILLER_83_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06865_ _06821_/A _06821_/B _06824_/A vssd1 vssd1 vccd1 vccd1 _06866_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09653_ _09653_/A _09600_/A vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__or2b_1
X_05816_ _06065_/A _05454_/A _05911_/A vssd1 vssd1 vccd1 vccd1 _05816_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08604_ _08600_/X _08597_/B _08498_/X vssd1 vssd1 vccd1 vccd1 _08604_/Y sky130_fd_sc_hd__a21oi_1
X_09584_ _09767_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09594_/A sky130_fd_sc_hd__or2_1
XFILLER_43_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08535_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10291_/S sky130_fd_sc_hd__clkbuf_4
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06796_ _06796_/A _06796_/B vssd1 vssd1 vccd1 vccd1 _06836_/A sky130_fd_sc_hd__xor2_2
X_05747_ _08282_/A _10563_/Q _10562_/Q _05746_/Y vssd1 vssd1 vccd1 vccd1 _05747_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05678_ _05771_/A _05588_/X _05580_/X _08304_/A _05677_/X vssd1 vssd1 vccd1 vccd1
+ _05678_/X sky130_fd_sc_hd__a221o_1
X_08466_ _10776_/Q vssd1 vssd1 vccd1 vccd1 _08572_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08397_ _08419_/A vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07417_ _07417_/A vssd1 vssd1 vccd1 vccd1 _07713_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07348_ _07489_/A _07481_/B vssd1 vssd1 vccd1 vccd1 _07482_/A sky130_fd_sc_hd__nor2_1
XFILLER_109_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07279_ _07302_/A _07279_/B _07344_/A vssd1 vssd1 vccd1 vccd1 _07289_/A sky130_fd_sc_hd__nor3_1
XANTENNA__07443__A1 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__B2 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09018_ _07442_/X _09015_/X _10537_/C vssd1 vssd1 vccd1 vccd1 _09018_/X sky130_fd_sc_hd__mux2_1
X_10290_ _10287_/D _10278_/Y _10287_/C vssd1 vssd1 vccd1 vccd1 _10300_/B sky130_fd_sc_hd__a21bo_1
XFILLER_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08171__A2 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05989__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10626_ _10806_/CLK _10626_/D vssd1 vssd1 vccd1 vccd1 _10626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _10666_/CLK _10557_/D vssd1 vssd1 vccd1 vccd1 _10557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10488_ _05958_/X _10475_/X _10487_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10967_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05874__D _05886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06650_ _06650_/A _06650_/B _06650_/C vssd1 vssd1 vccd1 vccd1 _06654_/A sky130_fd_sc_hd__and3_1
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05601_ _10560_/Q _05604_/A vssd1 vssd1 vccd1 vccd1 _05602_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06581_ _06581_/A _06581_/B _06581_/C vssd1 vssd1 vccd1 vccd1 _06593_/A sky130_fd_sc_hd__or3_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08320_ _08263_/A _08327_/B _08316_/Y _08319_/X _08062_/X vssd1 vssd1 vccd1 vccd1
+ _08320_/X sky130_fd_sc_hd__o32a_1
X_05532_ _10547_/Q vssd1 vssd1 vccd1 vccd1 _05549_/A sky130_fd_sc_hd__inv_2
X_08251_ _08251_/A _08251_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08277_/C sky130_fd_sc_hd__and3_1
X_05463_ _07914_/A _07911_/A _07907_/A _07903_/A vssd1 vssd1 vccd1 vccd1 _05467_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07202_ _07201_/Y _07187_/B _07190_/A vssd1 vssd1 vccd1 vccd1 _07204_/B sky130_fd_sc_hd__a21oi_1
X_08182_ _08263_/A _08180_/Y _08189_/B _08258_/A vssd1 vssd1 vccd1 vccd1 _08182_/Y
+ sky130_fd_sc_hd__o31ai_1
X_05394_ _10621_/Q vssd1 vssd1 vccd1 vccd1 _05462_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_134_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07133_ _07133_/A _07133_/B vssd1 vssd1 vccd1 vccd1 _07134_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07064_ _10984_/Q vssd1 vssd1 vccd1 vccd1 _07149_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06015_ input7/X _07967_/A input4/X input9/X vssd1 vssd1 vccd1 vccd1 _08048_/A sky130_fd_sc_hd__or4b_1
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08925__A1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _08414_/A _08939_/C vssd1 vssd1 vccd1 vccd1 _08971_/B sky130_fd_sc_hd__nor2_2
XFILLER_59_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09705_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09707_/B sky130_fd_sc_hd__xnor2_1
X_06917_ _06917_/A _06918_/C vssd1 vssd1 vccd1 vccd1 _06940_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__08153__A2 _08043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07897_ _10606_/Q _07888_/X _07892_/X _07896_/Y vssd1 vssd1 vccd1 vccd1 _07898_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__xor2_2
XFILLER_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06848_ _06848_/A _06848_/B vssd1 vssd1 vccd1 vccd1 _06862_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_66_clock_A _10981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09567_ _09567_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09570_/A sky130_fd_sc_hd__xor2_1
X_06779_ _06779_/A _06779_/B vssd1 vssd1 vccd1 vccd1 _06781_/B sky130_fd_sc_hd__xnor2_1
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08518_ _10796_/Q _08514_/X _08517_/X _10759_/Q vssd1 vssd1 vccd1 vccd1 _10759_/D
+ sky130_fd_sc_hd__a22o_1
X_09498_ _09458_/A _09458_/C _09458_/B vssd1 vssd1 vccd1 vccd1 _09499_/C sky130_fd_sc_hd__a21bo_1
X_08449_ _10771_/Q _10734_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08450_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _06182_/X _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10411_/X sky130_fd_sc_hd__a21bo_1
XFILLER_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10342_ input16/X _10415_/A _10342_/S vssd1 vssd1 vccd1 vccd1 _10343_/B sky130_fd_sc_hd__mux2_1
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08916__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10273_ _06997_/B _10115_/X _10271_/X _10272_/Y vssd1 vssd1 vccd1 vccd1 _10906_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input48_A io_wbs_m2s_sel[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10239__B1 _08514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08301__C1 _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06327__B _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10609_ _10851_/CLK _10609_/D vssd1 vssd1 vccd1 vccd1 _10609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07820_ _10869_/Q _07824_/B vssd1 vssd1 vccd1 vccd1 _07820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06997__B _06997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _07751_/A _07597_/B vssd1 vssd1 vccd1 vccd1 _07751_/X sky130_fd_sc_hd__or2b_1
XFILLER_65_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06702_ _06652_/B _06702_/B vssd1 vssd1 vccd1 vccd1 _06702_/X sky130_fd_sc_hd__and2b_1
XANTENNA__06146__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07682_ _07682_/A _07682_/B _09303_/B vssd1 vssd1 vccd1 vccd1 _09313_/B sky130_fd_sc_hd__and3_1
X_06633_ _06633_/A _06633_/B vssd1 vssd1 vccd1 vccd1 _06634_/B sky130_fd_sc_hd__or2_1
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09422_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ _10906_/Q _10890_/Q vssd1 vssd1 vccd1 vccd1 _09353_/B sky130_fd_sc_hd__and2b_1
X_06564_ _06564_/A _06564_/B _06584_/A vssd1 vssd1 vccd1 vccd1 _06571_/C sky130_fd_sc_hd__or3_1
XANTENNA__07621__B _07702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08303_ _08303_/A vssd1 vssd1 vccd1 vccd1 _10704_/D sky130_fd_sc_hd__clkbuf_1
X_05515_ _05340_/X _05510_/X _05513_/X _07900_/A vssd1 vssd1 vccd1 vccd1 _10564_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09283_ _10827_/Q _09274_/X _09275_/X _09282_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09284_/B sky130_fd_sc_hd__a32o_1
X_06495_ _06502_/B _06502_/C vssd1 vssd1 vccd1 vccd1 _06496_/A sky130_fd_sc_hd__and2_1
X_08234_ _08228_/A _08228_/B _08232_/A vssd1 vssd1 vccd1 vccd1 _08234_/X sky130_fd_sc_hd__a21o_1
X_05446_ _07919_/A _05326_/X _05324_/X _10645_/Q _05445_/X vssd1 vssd1 vccd1 vccd1
+ _05446_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08733__A _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08165_ _08355_/B vssd1 vssd1 vccd1 vccd1 _08165_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05377_ _06039_/A _05383_/A vssd1 vssd1 vccd1 vccd1 _05380_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07116_ _10984_/Q _07229_/B vssd1 vssd1 vccd1 vccd1 _07135_/B sky130_fd_sc_hd__nand2_1
X_08096_ _08096_/A vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07047_ _07472_/A _07472_/B vssd1 vssd1 vccd1 vccd1 _07473_/A sky130_fd_sc_hd__nand2_1
X_08998_ _08062_/X _08972_/X _08974_/X _08997_/X vssd1 vssd1 vccd1 vccd1 _08998_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07949_ _07949_/A vssd1 vssd1 vccd1 vccd1 _10651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10960_ _10960_/CLK _10960_/D vssd1 vssd1 vccd1 vccd1 _10960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10891_ _10909_/CLK _10891_/D vssd1 vssd1 vccd1 vccd1 _10891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _09619_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09620_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09087__A0 _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05332__A _08021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07958__S _07983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05986__B input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06073__B1 _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06163__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10325_ _10944_/Q _10960_/Q vssd1 vssd1 vccd1 vccd1 _10325_/X sky130_fd_sc_hd__or2b_1
XFILLER_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _10954_/Q _10938_/Q vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__and2b_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07706__B _07706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10187_ _09379_/B _10181_/X _10184_/X _10896_/Q vssd1 vssd1 vccd1 vccd1 _10896_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06983__D _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05300_ _10661_/Q _10660_/Q _05886_/A vssd1 vssd1 vccd1 vccd1 _05369_/A sky130_fd_sc_hd__nor3_2
X_06280_ _06558_/B _06360_/A vssd1 vssd1 vccd1 vccd1 _06281_/B sky130_fd_sc_hd__xor2_2
XFILLER_30_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_14_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06064__B1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09983_/A sky130_fd_sc_hd__or2_1
X_08921_ _08921_/A _08921_/B vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09384__A _09417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08852_ _08870_/B _08852_/B vssd1 vssd1 vccd1 vccd1 _08852_/X sky130_fd_sc_hd__xor2_1
XANTENNA__06801__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07803_ _07803_/A _07803_/B vssd1 vssd1 vccd1 vccd1 _10117_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07616__B _09898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08108__A2 _08043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08783_ _08773_/A _08778_/B _08803_/B vssd1 vssd1 vccd1 vccd1 _08783_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_84_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05995_ input51/X vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__inv_4
X_07734_ _07734_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07735_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07665_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__or2_1
XFILLER_26_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09404_ _09402_/A _09402_/B _09402_/C vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__a21oi_1
X_06616_ _06616_/A _06616_/B vssd1 vssd1 vccd1 vccd1 _06616_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07596_ _07596_/A _07718_/A vssd1 vssd1 vccd1 vccd1 _07597_/B sky130_fd_sc_hd__xnor2_4
XFILLER_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06547_ _06568_/A _10973_/Q _06547_/C _06567_/B vssd1 vssd1 vccd1 vccd1 _06549_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ _09316_/A _09337_/B _09334_/X vssd1 vssd1 vccd1 vccd1 _09336_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__08292__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _09289_/A _09266_/B vssd1 vssd1 vccd1 vccd1 _09267_/A sky130_fd_sc_hd__and2_1
X_06478_ _06478_/A _06478_/B vssd1 vssd1 vccd1 vccd1 _06480_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08217_ _08216_/X _08218_/B _08058_/A vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__a21bo_1
X_05429_ _07882_/A _05353_/X _05350_/X _10635_/Q _05428_/X vssd1 vssd1 vccd1 vccd1
+ _05429_/X sky130_fd_sc_hd__a221o_1
X_09197_ _09113_/A _09196_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08148_ _08148_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08169_/C sky130_fd_sc_hd__and2_1
XFILLER_107_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08075_/A _08075_/B _05733_/X vssd1 vssd1 vccd1 vccd1 _08079_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__06055__B1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09294__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ _10110_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10041_ _09964_/X _09967_/B _09965_/A vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__a21o_1
XFILLER_76_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10943_ _10945_/CLK _10943_/D vssd1 vssd1 vccd1 vccd1 _10943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10874_ _10960_/CLK _10874_/D vssd1 vssd1 vccd1 vccd1 _10874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05997__A _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08035__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10308_ _10298_/A _10301_/Y _10297_/A vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10239_ _10246_/C _10238_/X _08514_/A vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__o21ai_1
X_05780_ _10566_/Q vssd1 vssd1 vccd1 vccd1 _05780_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07450_ _07450_/A _07551_/B vssd1 vssd1 vccd1 vccd1 _07451_/B sky130_fd_sc_hd__xor2_1
XFILLER_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07381_ _07381_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07458_/B sky130_fd_sc_hd__xnor2_1
X_06401_ _06845_/A _06627_/B vssd1 vssd1 vccd1 vccd1 _06630_/A sky130_fd_sc_hd__and2_1
X_09120_ _09114_/X _09117_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__o21a_1
X_06332_ _06388_/A vssd1 vssd1 vccd1 vccd1 _06804_/A sky130_fd_sc_hd__clkbuf_2
X_09051_ _09042_/X _09050_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10837_/D sky130_fd_sc_hd__o21a_2
XANTENNA__10963__D _10963_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ _08015_/A vssd1 vssd1 vccd1 vccd1 _08002_/X sky130_fd_sc_hd__clkbuf_2
X_06263_ _10918_/Q _10901_/Q vssd1 vssd1 vccd1 vccd1 _06263_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08026__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06194_ _06191_/X _06183_/X _06193_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10596_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09953_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09953_/Y sky130_fd_sc_hd__inv_2
XFILLER_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09884_ _09812_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__and2b_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08835_ _08825_/A _08828_/Y _08841_/C vssd1 vssd1 vccd1 vccd1 _08835_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08758_/A _08761_/Y _08804_/C vssd1 vssd1 vccd1 vccd1 _08766_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_73_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05978_ _05286_/B _05975_/X _05977_/X vssd1 vssd1 vccd1 vccd1 _05978_/Y sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_50_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10826_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07717_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07720_/A sky130_fd_sc_hd__xnor2_1
X_08697_ _08688_/X _08693_/Y _08696_/X vssd1 vssd1 vccd1 vccd1 _10802_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07648_ _07655_/A _07648_/B vssd1 vssd1 vccd1 vccd1 _07649_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_65_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10889_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07579_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__or2_1
X_09318_ _09443_/B vssd1 vssd1 vccd1 vccd1 _09536_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_41_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10590_ _10813_/CLK _10590_/D vssd1 vssd1 vccd1 vccd1 _10590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09249_ _09249_/A vssd1 vssd1 vccd1 vccd1 _10856_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_126_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08017__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__A0 _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09736__B _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput54 _05954_/X vssd1 vssd1 vccd1 vccd1 io_pwm_low sky130_fd_sc_hd__buf_2
Xoutput65 _10852_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[18] sky130_fd_sc_hd__buf_2
Xoutput76 _10862_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[28] sky130_fd_sc_hd__buf_2
XFILLER_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput87 _10843_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_1_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input30_A io_wbs_m2s_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10024_ _09828_/B _09830_/X _10095_/B vssd1 vssd1 vccd1 vccd1 _10025_/B sky130_fd_sc_hd__a21boi_1
XFILLER_49_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_clock _10857_/CLK vssd1 vssd1 vccd1 vccd1 _10651_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10926_ _10930_/CLK _10926_/D vssd1 vssd1 vccd1 vccd1 _10926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10857_ _10857_/CLK _10857_/D vssd1 vssd1 vccd1 vccd1 _10857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10790_/CLK _10788_/D vssd1 vssd1 vccd1 vccd1 _10788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10138__A _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09205__A0 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06950_ _06950_/A _06952_/A vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__xnor2_1
X_05901_ _10654_/Q vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__buf_2
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06881_ _06881_/A _06881_/B vssd1 vssd1 vccd1 vccd1 _06932_/B sky130_fd_sc_hd__xor2_4
X_05832_ _08342_/A _05836_/A _05827_/Y vssd1 vssd1 vccd1 vccd1 _05947_/B sky130_fd_sc_hd__a21oi_1
XFILLER_121_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08620_ _08620_/A vssd1 vssd1 vccd1 vccd1 _10789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05763_ _08228_/A _10558_/Q _10557_/Q _05744_/Y vssd1 vssd1 vccd1 vccd1 _05789_/A
+ sky130_fd_sc_hd__o22a_1
X_08551_ _10198_/A _08550_/X _08462_/A vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05694_ _10551_/Q vssd1 vssd1 vccd1 vccd1 _05694_/Y sky130_fd_sc_hd__inv_2
X_08482_ _10781_/Q _10744_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08483_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07502_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07910__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07433_ _07433_/A vssd1 vssd1 vccd1 vccd1 _07728_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ _09113_/A _09102_/X _10518_/B vssd1 vssd1 vccd1 vccd1 _09103_/Y sky130_fd_sc_hd__o21ai_1
X_07364_ _07410_/A _07364_/B vssd1 vssd1 vccd1 vccd1 _07366_/C sky130_fd_sc_hd__nand2_1
XFILLER_136_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06315_ _10925_/Q _09344_/B vssd1 vssd1 vccd1 vccd1 _06317_/A sky130_fd_sc_hd__nand2_1
X_07295_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07296_/B sky130_fd_sc_hd__and2_1
XFILLER_108_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06246_ _10612_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06246_/X sky130_fd_sc_hd__or2_1
X_09034_ _09023_/X _09025_/X _09033_/X _06137_/X vssd1 vssd1 vccd1 vccd1 _10836_/D
+ sky130_fd_sc_hd__o31a_2
XANTENNA__05481__A1 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09747__A1 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06177_ _06172_/X _06158_/X _06175_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10592_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09936_ _10009_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09572__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09867_ _09867_/A _09867_/B _09937_/A _09867_/D vssd1 vssd1 vccd1 vccd1 _09868_/B
+ sky130_fd_sc_hd__and4_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08818_ _08817_/A _08817_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08818_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10511__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07804__B _10117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ _09432_/A _09735_/B _09735_/A vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__o21a_1
X_08749_ _06172_/X _08728_/X _08729_/X _08748_/X vssd1 vssd1 vccd1 vccd1 _08749_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10711_ _10845_/CLK _10711_/D vssd1 vssd1 vccd1 vccd1 _10711_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08238__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10642_ _10646_/CLK _10642_/D vssd1 vssd1 vccd1 vccd1 _10642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _10832_/CLK _10573_/D vssd1 vssd1 vccd1 vccd1 _10573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10007_ _10077_/B _10007_/B vssd1 vssd1 vccd1 vccd1 _10009_/C sky130_fd_sc_hd__nand2_1
XFILLER_49_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10909_/CLK _10909_/D vssd1 vssd1 vccd1 vccd1 _10909_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__08229__A1 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08229__B2 _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06100_ _10692_/Q _10691_/Q _10690_/Q _08160_/B vssd1 vssd1 vccd1 vccd1 _08191_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07080_ _07070_/A _07070_/B _07298_/A vssd1 vssd1 vccd1 vccd1 _07089_/A sky130_fd_sc_hd__a21bo_1
X_06031_ _10582_/Q vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07982_ _06187_/X _07965_/X _07981_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10659_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09721_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09723_/C sky130_fd_sc_hd__xnor2_1
X_06933_ _06935_/A _06935_/B _06932_/X vssd1 vssd1 vccd1 vccd1 _06934_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06864_ _06864_/A _06864_/B vssd1 vssd1 vccd1 vccd1 _06867_/B sky130_fd_sc_hd__xnor2_1
X_09652_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09662_/B sky130_fd_sc_hd__and2_1
X_05815_ _05405_/A _05482_/X _05814_/X vssd1 vssd1 vccd1 vccd1 _05911_/A sky130_fd_sc_hd__o21ai_1
XFILLER_94_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08603_ _08603_/A vssd1 vssd1 vccd1 vccd1 _10784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09583_ _10969_/Q _09744_/B _09671_/A vssd1 vssd1 vccd1 vccd1 _09584_/B sky130_fd_sc_hd__a21boi_1
X_06795_ _06763_/A _06763_/B _06766_/A vssd1 vssd1 vccd1 vccd1 _06796_/B sky130_fd_sc_hd__a21oi_2
X_05746_ _08277_/B vssd1 vssd1 vccd1 vccd1 _05746_/Y sky130_fd_sc_hd__inv_2
X_08534_ _10251_/S _10768_/Q _10767_/Q vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__and3_1
XFILLER_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05677_ _08285_/A _05590_/X _05588_/X _05771_/A _05676_/X vssd1 vssd1 vccd1 vccd1
+ _05677_/X sky130_fd_sc_hd__o221a_1
X_08465_ _08465_/A vssd1 vssd1 vccd1 vccd1 _10738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06256__A _08837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08396_ _08383_/X _10739_/Q _08394_/X hold19/X vssd1 vssd1 vccd1 vccd1 _10721_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07416_ _07416_/A vssd1 vssd1 vccd1 vccd1 _07732_/A sky130_fd_sc_hd__buf_4
XFILLER_137_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07347_ _07347_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07481_/B sky130_fd_sc_hd__xor2_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09017_ _10523_/A vssd1 vssd1 vccd1 vccd1 _10537_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_07278_ _07308_/A _07319_/A _07308_/C vssd1 vssd1 vccd1 vccd1 _07344_/A sky130_fd_sc_hd__o21ai_2
XFILLER_136_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06229_ _10605_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06229_/X sky130_fd_sc_hd__or2_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10506__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09919_ _10057_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _10056_/C sky130_fd_sc_hd__nand2_1
XFILLER_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ _10803_/CLK _10625_/D vssd1 vssd1 vccd1 vccd1 _10625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10556_ _10666_/CLK _10556_/D vssd1 vssd1 vccd1 vccd1 _10556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10487_/X sky130_fd_sc_hd__or2_1
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05600_ _10699_/Q vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06580_ _06594_/A _06594_/B _06579_/Y vssd1 vssd1 vccd1 vccd1 _06607_/B sky130_fd_sc_hd__o21bai_1
X_05531_ _10554_/Q vssd1 vssd1 vccd1 vccd1 _05663_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08250_ _08157_/X _08245_/Y _08247_/Y _08249_/X vssd1 vssd1 vccd1 vccd1 _10699_/D
+ sky130_fd_sc_hd__o31a_1
X_05462_ _05462_/A _05462_/B _05462_/C _05462_/D vssd1 vssd1 vccd1 vccd1 _05462_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08181_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08189_/B sky130_fd_sc_hd__nor2_1
X_07201_ _07201_/A vssd1 vssd1 vccd1 vccd1 _07201_/Y sky130_fd_sc_hd__inv_2
X_05393_ _10621_/Q _05393_/B vssd1 vssd1 vccd1 vccd1 _05393_/X sky130_fd_sc_hd__and2_1
X_07132_ _07132_/A _07132_/B vssd1 vssd1 vccd1 vccd1 _07285_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07063_ _07086_/B _07188_/B vssd1 vssd1 vccd1 vccd1 _07070_/A sky130_fd_sc_hd__and2_1
X_06014_ input50/X input48/X vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__nand2_4
XFILLER_133_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07965_ _08034_/B vssd1 vssd1 vccd1 vccd1 _07965_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07635__A _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09704_ _09644_/A _09769_/C _09703_/X vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__o21a_1
X_06916_ _06916_/A _06916_/B vssd1 vssd1 vccd1 vccd1 _06918_/C sky130_fd_sc_hd__nor2_2
X_07896_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07896_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09635_ hold9/A _09572_/X _09631_/X _09634_/Y vssd1 vssd1 vccd1 vccd1 _10873_/D sky130_fd_sc_hd__a22o_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06847_ _06847_/A _06847_/B vssd1 vssd1 vccd1 vccd1 _06848_/B sky130_fd_sc_hd__nor2_1
XFILLER_70_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09566_ _09566_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__xnor2_2
X_06778_ _06792_/A _06778_/B vssd1 vssd1 vccd1 vccd1 _06781_/A sky130_fd_sc_hd__nor2_1
X_05729_ _10546_/Q vssd1 vssd1 vccd1 vccd1 _05729_/Y sky130_fd_sc_hd__inv_2
X_08517_ _10177_/A vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09497_ _09542_/A _09496_/C _09496_/A vssd1 vssd1 vccd1 vccd1 _09499_/B sky130_fd_sc_hd__a21o_1
X_08448_ _08448_/A vssd1 vssd1 vccd1 vccd1 _10733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08379_ _08367_/X _10733_/Q _07865_/X _08378_/X vssd1 vssd1 vccd1 vccd1 _10715_/D
+ sky130_fd_sc_hd__o211a_1
X_10410_ _10941_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10410_/X sky130_fd_sc_hd__and2_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _10341_/A _10341_/B _10341_/C vssd1 vssd1 vccd1 vccd1 _10342_/S sky130_fd_sc_hd__or3_1
XFILLER_105_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10272_ _10287_/A _10271_/B _09480_/X vssd1 vssd1 vccd1 vccd1 _10272_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08377__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ _10830_/CLK _10608_/D vssd1 vssd1 vccd1 vccd1 _10608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10539_ _08974_/X _08969_/Y _09036_/X _06137_/X vssd1 vssd1 vccd1 vccd1 _10987_/D
+ sky130_fd_sc_hd__o31a_4
XANTENNA__10411__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07158__C _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07750_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__xor2_2
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06701_ _06903_/A _06903_/B _06700_/X vssd1 vssd1 vccd1 vccd1 _06893_/B sky130_fd_sc_hd__a21o_2
XANTENNA_clkbuf_leaf_10_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07681_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__xor2_1
XFILLER_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06632_ _06633_/A _06633_/B vssd1 vssd1 vccd1 vccd1 _06634_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09420_ _09420_/A _10885_/Q vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__and2_1
XANTENNA__10966__D _10966_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _10890_/Q _10906_/Q vssd1 vssd1 vccd1 vccd1 _09371_/B sky130_fd_sc_hd__and2b_1
X_06563_ _10974_/Q _10973_/Q _06575_/B _06587_/A vssd1 vssd1 vccd1 vccd1 _06584_/A
+ sky130_fd_sc_hd__and4_1
X_08302_ _08300_/X _08302_/B vssd1 vssd1 vccd1 vccd1 _08303_/A sky130_fd_sc_hd__and2b_1
X_09282_ _08027_/A _09281_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09282_/X sky130_fd_sc_hd__mux2_1
X_05514_ _05343_/Y _05510_/X _05513_/X _07896_/A vssd1 vssd1 vccd1 vccd1 _10563_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _08233_/A _08233_/B vssd1 vssd1 vccd1 vccd1 _08233_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06494_ _10971_/Q vssd1 vssd1 vccd1 vccd1 _06502_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05445_ _07914_/A _05329_/X _05326_/X _10644_/Q _05444_/X vssd1 vssd1 vccd1 vccd1
+ _05445_/X sky130_fd_sc_hd__o221a_1
X_08164_ _08248_/A vssd1 vssd1 vccd1 vccd1 _08164_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05376_ _10626_/Q vssd1 vssd1 vccd1 vccd1 _05461_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08095_ _08095_/A _08095_/B vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07115_ _07222_/B vssd1 vssd1 vccd1 vccd1 _07229_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06253__B _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10056__A _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ _07421_/A _07046_/B vssd1 vssd1 vccd1 vccd1 _07472_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09571__A2 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _05813_/A _08976_/X _08994_/X _08996_/Y _09078_/B vssd1 vssd1 vccd1 vccd1
+ _08997_/X sky130_fd_sc_hd__a221o_1
XFILLER_87_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07948_ _07955_/A _07948_/B vssd1 vssd1 vccd1 vccd1 _07949_/A sky130_fd_sc_hd__or2_1
X_07879_ _10601_/Q _07870_/X _07874_/X _07878_/Y vssd1 vssd1 vccd1 vccd1 _07880_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10890_ _10909_/CLK _10890_/D vssd1 vssd1 vccd1 vccd1 _10890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ _09618_/A _09618_/B _09618_/C vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__or3_1
X_09549_ _09549_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09610_/C sky130_fd_sc_hd__xor2_2
XFILLER_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08643__B _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ _10324_/A _10334_/A vssd1 vssd1 vccd1 vccd1 _10330_/A sky130_fd_sc_hd__or2_1
XFILLER_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10255_ _10938_/Q _10954_/Q vssd1 vssd1 vccd1 vccd1 _10257_/A sky130_fd_sc_hd__and2b_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10186_ _07570_/A _10181_/X _10184_/X _10895_/Q vssd1 vssd1 vccd1 vccd1 _10895_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07869__A_N _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06064__A1 _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06064__B2 _09104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08927_/C sky130_fd_sc_hd__nand2_1
XFILLER_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08210__C1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08851_ _08847_/X _08815_/B _08845_/Y vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__a21o_1
XFILLER_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07802_ _07802_/A _07802_/B vssd1 vssd1 vccd1 vccd1 _07803_/B sky130_fd_sc_hd__xnor2_2
X_05994_ _07880_/A _05994_/B vssd1 vssd1 vccd1 vccd1 _10576_/D sky130_fd_sc_hd__nor2_1
X_08782_ _10812_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08803_/B sky130_fd_sc_hd__xor2_1
XFILLER_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07733_ _07733_/A _07733_/B vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07664_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09403_ _09403_/A _09403_/B vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__nand2_4
XFILLER_53_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06615_ _06681_/A _06674_/C _06674_/A vssd1 vssd1 vccd1 vccd1 _06672_/B sky130_fd_sc_hd__a21bo_1
XFILLER_25_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07595_ _07397_/A _07397_/B _07594_/X vssd1 vssd1 vccd1 vccd1 _07718_/A sky130_fd_sc_hd__a21oi_4
X_06546_ _06546_/A _06602_/A vssd1 vssd1 vccd1 vccd1 _06618_/A sky130_fd_sc_hd__xnor2_2
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09334_ _10883_/Q _07098_/A vssd1 vssd1 vccd1 vccd1 _09334_/X sky130_fd_sc_hd__or2b_1
XANTENNA__08292__A2 _08212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09265_ _10824_/Q _09243_/X _09244_/X _09264_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09266_/B sky130_fd_sc_hd__a32o_1
X_06477_ _06477_/A _06477_/B vssd1 vssd1 vccd1 vccd1 _06478_/B sky130_fd_sc_hd__and2_1
X_08216_ _08218_/A vssd1 vssd1 vccd1 vccd1 _08216_/X sky130_fd_sc_hd__clkbuf_2
X_05428_ _07878_/A _05358_/X _05353_/X _10634_/Q _05427_/X vssd1 vssd1 vccd1 vccd1
+ _05428_/X sky130_fd_sc_hd__o221a_1
X_09196_ _09114_/A _09195_/X _10500_/B vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08150_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08147_/X sky130_fd_sc_hd__or2_1
XFILLER_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05359_ _10632_/Q vssd1 vssd1 vccd1 vccd1 _07875_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08078_ _08073_/X _08076_/X _08077_/X vssd1 vssd1 vccd1 vccd1 _10682_/D sky130_fd_sc_hd__o21a_1
XANTENNA__06055__B2 _09104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07029_ _07044_/A _07030_/C _07417_/A _07021_/A vssd1 vssd1 vccd1 vccd1 _07031_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_121_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _10040_/A _10039_/Y vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__or2b_1
XFILLER_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07823__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10942_ _10962_/CLK _10942_/D vssd1 vssd1 vccd1 vccd1 _10942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10873_ _10958_/CLK _10873_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06174__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08035__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10307_ _10307_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__nor2_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _10236_/X _10237_/Y _10279_/S vssd1 vssd1 vccd1 vccd1 _10238_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10169_ _07098_/A _10167_/X _08517_/X _10883_/Q vssd1 vssd1 vccd1 vccd1 _10883_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06400_ _06441_/B vssd1 vssd1 vccd1 vccd1 _06845_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08259__C1 _08258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07380_ _07459_/B _07490_/A _07327_/X vssd1 vssd1 vccd1 vccd1 _07381_/B sky130_fd_sc_hd__a21bo_1
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06331_ _06342_/A _06342_/B vssd1 vssd1 vccd1 vccd1 _06388_/A sky130_fd_sc_hd__xnor2_1
X_09050_ _10484_/A _10474_/B _10495_/B _10506_/A _09049_/X vssd1 vssd1 vccd1 vccd1
+ _09050_/X sky130_fd_sc_hd__a221o_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06262_ _06262_/A _06262_/B vssd1 vssd1 vccd1 vccd1 _06305_/A sky130_fd_sc_hd__nand2_4
X_08001_ input24/X _07987_/X _08000_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10665_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06193_ _06193_/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06193_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09952_ _09952_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__xnor2_1
X_08903_ _10827_/Q _08919_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__nor2_1
XFILLER_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09883_ _09883_/A vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__inv_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ _10818_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08841_/C sky130_fd_sc_hd__xor2_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08765_ _10810_/Q _08801_/B vssd1 vssd1 vccd1 vccd1 _08804_/C sky130_fd_sc_hd__xor2_2
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05977_ _08445_/A vssd1 vssd1 vccd1 vccd1 _05977_/X sky130_fd_sc_hd__buf_2
XFILLER_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07716_ _07442_/X _07574_/B _07715_/X vssd1 vssd1 vccd1 vccd1 _07717_/B sky130_fd_sc_hd__a21o_1
X_08696_ _06147_/X _08694_/X _08695_/X _10802_/Q _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08696_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06259__A _10978_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07647_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__xnor2_1
XFILLER_41_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07578_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07580_/A sky130_fd_sc_hd__nand2_1
X_09317_ _09736_/B _09388_/A vssd1 vssd1 vccd1 vccd1 _09396_/B sky130_fd_sc_hd__nand2_2
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06529_ _06527_/A _06489_/B _06540_/A _06600_/A vssd1 vssd1 vccd1 vccd1 _06529_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09248_ _09259_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__and2_1
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09226_/S sky130_fd_sc_hd__buf_2
XFILLER_5_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08640__C _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput55 _10987_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_122_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput66 _10853_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[19] sky130_fd_sc_hd__buf_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput77 _10863_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[29] sky130_fd_sc_hd__buf_2
XFILLER_122_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10023_ _10023_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _10095_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input23_A io_wbs_m2s_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09150__B1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_57_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10925_ _10930_/CLK _10925_/D vssd1 vssd1 vccd1 vccd1 _10925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08384__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10856_ _10862_/CLK _10856_/D vssd1 vssd1 vccd1 vccd1 _10856_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10787_ _10790_/CLK _10787_/D vssd1 vssd1 vccd1 vccd1 _10787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05900_ _05900_/A _05900_/B vssd1 vssd1 vccd1 vccd1 _05900_/X sky130_fd_sc_hd__and2_1
XFILLER_95_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06880_ _07799_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _06934_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08192__B2 _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__A1 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05831_ _08027_/A _05831_/B _05831_/C vssd1 vssd1 vccd1 vccd1 _05836_/A sky130_fd_sc_hd__or3_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05762_ _05746_/Y _10562_/Q _10561_/Q _05751_/Y _05761_/X vssd1 vssd1 vccd1 vccd1
+ _05791_/A sky130_fd_sc_hd__o221a_1
X_08550_ _08661_/A vssd1 vssd1 vccd1 vccd1 _08550_/X sky130_fd_sc_hd__clkbuf_2
X_05693_ _05693_/A vssd1 vssd1 vccd1 vccd1 _08173_/A sky130_fd_sc_hd__buf_2
X_08481_ _08481_/A vssd1 vssd1 vccd1 vccd1 _10743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07501_ _07501_/A _07505_/A vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__and2_1
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07432_ _07563_/A vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ _09114_/A _09101_/X _09118_/A vssd1 vssd1 vccd1 vccd1 _09102_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07363_ _07361_/Y _07363_/B _07363_/C vssd1 vssd1 vccd1 vccd1 _07364_/B sky130_fd_sc_hd__nand3b_1
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06314_ _10908_/Q vssd1 vssd1 vccd1 vccd1 _09344_/B sky130_fd_sc_hd__clkbuf_4
X_07294_ _07309_/A _07309_/C _07309_/B vssd1 vssd1 vccd1 vccd1 _07310_/A sky130_fd_sc_hd__a21oi_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06245_ input35/X _06238_/X _06244_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10611_/D
+ sky130_fd_sc_hd__o211a_1
X_09033_ _07726_/A _09032_/X _10537_/C vssd1 vssd1 vccd1 vccd1 _09033_/X sky130_fd_sc_hd__mux2_1
X_06176_ _10343_/A vssd1 vssd1 vccd1 vccd1 _06176_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08707__B1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09866_ _09931_/A _09937_/A _10139_/S _09736_/B vssd1 vssd1 vccd1 vccd1 _09868_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08183__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08183__A1 _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08817_ _08817_/A _08817_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08817_/X sky130_fd_sc_hd__and3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09797_ _09797_/A _09797_/B vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__xnor2_2
XFILLER_46_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08748_ _10807_/Q vssd1 vssd1 vccd1 vccd1 _08748_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _10801_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08679_/X sky130_fd_sc_hd__and2_1
XFILLER_54_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10710_ _10710_/CLK _10710_/D vssd1 vssd1 vccd1 vccd1 _10710_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10641_ _10646_/CLK _10641_/D vssd1 vssd1 vccd1 vccd1 _10641_/Q sky130_fd_sc_hd__dfxtp_1
X_10572_ _10865_/CLK _10572_/D vssd1 vssd1 vccd1 vccd1 _10572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07997__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08174__B2 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08174__A1 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__or2_1
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10908_ _10924_/CLK _10908_/D vssd1 vssd1 vccd1 vccd1 _10908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10839_ _10839_/CLK _10839_/D vssd1 vssd1 vccd1 vccd1 _10839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09938__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07437__B1 _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06030_ _10581_/Q _06020_/X _06029_/X vssd1 vssd1 vccd1 vccd1 _10581_/D sky130_fd_sc_hd__o21a_1
XFILLER_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07981_ _07981_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07981_/X sky130_fd_sc_hd__or2_1
XFILLER_87_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10960_/CLK sky130_fd_sc_hd__clkbuf_16
X_09720_ _09716_/Y _09718_/Y _09719_/X vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__o21a_1
X_06932_ _06890_/B _06932_/B vssd1 vssd1 vccd1 vccd1 _06932_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08289__A _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10969__D _10969_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ _06863_/A _06863_/B vssd1 vssd1 vccd1 vccd1 _06864_/B sky130_fd_sc_hd__nor2_1
X_09651_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09662_/A sky130_fd_sc_hd__nor2_1
X_05814_ _05408_/Y _05643_/A _05813_/X vssd1 vssd1 vccd1 vccd1 _05814_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08602_ _08617_/B _08649_/A _08602_/C vssd1 vssd1 vccd1 vccd1 _08603_/A sky130_fd_sc_hd__and3b_1
XFILLER_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09582_ _10970_/Q _09744_/A vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06794_ _06832_/A _06794_/B vssd1 vssd1 vccd1 vccd1 _06796_/A sky130_fd_sc_hd__xor2_2
XFILLER_27_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05745_ _10702_/Q vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__07921__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ _08881_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _10767_/D sky130_fd_sc_hd__nor2_1
XFILLER_82_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05676_ _08277_/A _05593_/X _05590_/X _08285_/A _05675_/X vssd1 vssd1 vccd1 vccd1
+ _05676_/X sky130_fd_sc_hd__a221o_1
X_08464_ _08477_/A _08464_/B vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__or2_1
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _08395_/A _10755_/Q vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__or2_1
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07415_ _07415_/A _07472_/A _07415_/C _07434_/A vssd1 vssd1 vccd1 vccd1 _07428_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07346_ _07488_/B _07529_/A _07488_/A vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__o21ai_2
XFILLER_136_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_clock _10857_/CLK vssd1 vssd1 vccd1 vccd1 _10987_/CLK sky130_fd_sc_hd__clkbuf_16
X_09016_ _09016_/A _09016_/B vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__or2_1
X_07277_ _07277_/A _07277_/B vssd1 vssd1 vccd1 vccd1 _07308_/C sky130_fd_sc_hd__xnor2_1
XFILLER_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06228_ input28/X _06225_/X _06227_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10604_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06159_ _10589_/Q vssd1 vssd1 vccd1 vccd1 _06160_/A sky130_fd_sc_hd__inv_2
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _10031_/A sky130_fd_sc_hd__xnor2_2
XFILLER_59_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09849_ _09901_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09851_/C sky130_fd_sc_hd__xor2_1
XFILLER_58_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10624_ _10803_/CLK _10624_/D vssd1 vssd1 vccd1 vccd1 _10624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ _10695_/CLK _10555_/D vssd1 vssd1 vccd1 vccd1 _10555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06182__A input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ _06147_/X _10475_/X _10484_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10966_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08837__A _08837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05530_ _10567_/Q vssd1 vssd1 vccd1 vccd1 _05769_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05461_ _05461_/A _05461_/B _05461_/C _05461_/D vssd1 vssd1 vccd1 vccd1 _05462_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08180_ _08180_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _08180_/Y sky130_fd_sc_hd__nor2_1
X_05392_ _05392_/A _05392_/B vssd1 vssd1 vccd1 vccd1 _05393_/B sky130_fd_sc_hd__nor2_1
X_07200_ _07200_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _07204_/A sky130_fd_sc_hd__xnor2_1
X_07131_ _07377_/A _07229_/B _07147_/A vssd1 vssd1 vccd1 vccd1 _07132_/B sky130_fd_sc_hd__and3_1
XFILLER_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07062_ _07164_/B vssd1 vssd1 vccd1 vccd1 _07188_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06013_ _06008_/X _05975_/X _06012_/Y vssd1 vssd1 vccd1 vccd1 _10579_/D sky130_fd_sc_hd__o21a_1
XFILLER_114_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10193__B2 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07964_ _07964_/A vssd1 vssd1 vccd1 vccd1 _08034_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_114_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07895_ _07898_/A _07895_/B vssd1 vssd1 vccd1 vccd1 _10637_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _09703_/A _09703_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__or3b_1
X_06915_ _06915_/A _06915_/B _06942_/A vssd1 vssd1 vccd1 vccd1 _06916_/B sky130_fd_sc_hd__nor3_1
XFILLER_28_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09634_ _09634_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__nor2_1
X_06846_ _10508_/A _07784_/B _06845_/C vssd1 vssd1 vccd1 vccd1 _06847_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09565_ _09625_/A _09625_/B _09626_/A vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__o21a_1
X_06777_ _06900_/A _07783_/B _06775_/C vssd1 vssd1 vccd1 vccd1 _06778_/B sky130_fd_sc_hd__a21oi_1
X_05728_ _06037_/A vssd1 vssd1 vccd1 vccd1 _05728_/X sky130_fd_sc_hd__clkbuf_2
X_08516_ _10795_/Q _08514_/X _08509_/X _10758_/Q vssd1 vssd1 vccd1 vccd1 _10758_/D
+ sky130_fd_sc_hd__a22o_1
X_09496_ _09496_/A _09542_/A _09496_/C vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__nand3_1
X_05659_ _05896_/A _05628_/X _05626_/X _08148_/A _05658_/X vssd1 vssd1 vccd1 vccd1
+ _05659_/X sky130_fd_sc_hd__o221a_1
X_08447_ _08460_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08448_/A sky130_fd_sc_hd__or2_1
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08378_ _08381_/A hold27/X vssd1 vssd1 vccd1 vccd1 _08378_/X sky130_fd_sc_hd__or2_1
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10517__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ _07562_/A _07327_/X _07511_/A _07328_/Y vssd1 vssd1 vccd1 vccd1 _07333_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10420__A2 _10724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ _10914_/Q vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10271_ _10287_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10271_/X sky130_fd_sc_hd__or2_1
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08657__A _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07561__A _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_6_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _10830_/CLK _10607_/D vssd1 vssd1 vccd1 vccd1 _10607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10538_ _07592_/A _10522_/A _10537_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10986_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10469_ _10961_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10469_/X sky130_fd_sc_hd__or2_1
XFILLER_69_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10357__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07591__A2 _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06700_ _06665_/B _06700_/B vssd1 vssd1 vccd1 vccd1 _06700_/X sky130_fd_sc_hd__and2b_1
X_07680_ _07680_/A _07680_/B vssd1 vssd1 vccd1 vccd1 _07681_/B sky130_fd_sc_hd__xnor2_1
XFILLER_92_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06631_ _06631_/A _06631_/B vssd1 vssd1 vccd1 vccd1 _06633_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09350_ _09371_/A _09372_/B vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__or2_1
X_06562_ _06585_/A _06585_/B _06573_/C vssd1 vssd1 vccd1 vccd1 _06564_/B sky130_fd_sc_hd__and3_1
X_08301_ input32/X _08248_/A _08052_/A _08297_/A _08175_/A vssd1 vssd1 vccd1 vccd1
+ _08302_/B sky130_fd_sc_hd__o221a_1
X_09281_ _08332_/A _07919_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09281_/X sky130_fd_sc_hd__mux2_1
X_05513_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05513_/X sky130_fd_sc_hd__clkbuf_2
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08251_/C sky130_fd_sc_hd__nor2_2
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06493_ _06527_/A _06513_/D _06493_/C vssd1 vssd1 vccd1 vccd1 _06510_/A sky130_fd_sc_hd__and3_1
XFILLER_33_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05444_ _10643_/Q _05329_/X _05438_/X _07911_/A _05443_/X vssd1 vssd1 vccd1 vccd1
+ _05444_/X sky130_fd_sc_hd__a221o_1
XANTENNA__06815__A _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08163_ _08158_/X _08169_/C _08162_/Y vssd1 vssd1 vccd1 vccd1 _08163_/Y sky130_fd_sc_hd__a21oi_1
X_05375_ _10627_/Q vssd1 vssd1 vccd1 vccd1 _05461_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ _08098_/A _08095_/B vssd1 vssd1 vccd1 vccd1 _08094_/X sky130_fd_sc_hd__or2_1
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07114_ _07216_/B vssd1 vssd1 vccd1 vccd1 _07222_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_134_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07045_ _07573_/A _07434_/A _07509_/A vssd1 vssd1 vccd1 vccd1 _07046_/B sky130_fd_sc_hd__and3_1
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10166__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08996_ _05721_/Y _06212_/B _08995_/X vssd1 vssd1 vccd1 vccd1 _08996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07947_ input41/X _05279_/A _07964_/A vssd1 vssd1 vccd1 vccd1 _07948_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07878_ _07878_/A vssd1 vssd1 vccd1 vccd1 _07878_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06829_ _06882_/A _06883_/A _06882_/B vssd1 vssd1 vccd1 vccd1 _06884_/A sky130_fd_sc_hd__and3_1
XFILLER_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09617_ _09545_/B _09617_/B vssd1 vssd1 vccd1 vccd1 _09618_/C sky130_fd_sc_hd__and2b_1
X_09548_ _09432_/A _09508_/B _09508_/A vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__o21ai_2
XFILLER_34_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09479_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06073__A2 _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10323_ _10945_/Q _10961_/Q vssd1 vssd1 vccd1 vccd1 _10334_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10254_ _07061_/A _10253_/A _10253_/Y _08563_/X vssd1 vssd1 vccd1 vccd1 _10904_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06460__A _10978_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10185_ _09920_/B _10181_/X _10184_/X _10894_/Q vssd1 vssd1 vccd1 vccd1 _10894_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06064__A2 _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08850_ _10820_/Q _08865_/B vssd1 vssd1 vccd1 vccd1 _08870_/B sky130_fd_sc_hd__xor2_2
XFILLER_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07801_ _07801_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__xnor2_1
X_05993_ _05992_/X _09107_/A _05993_/S vssd1 vssd1 vccd1 vccd1 _05994_/B sky130_fd_sc_hd__mux2_1
X_08781_ _08778_/X _08779_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10811_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07732_ _07732_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07733_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07663_ _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09402_ _09402_/A _09402_/B _09402_/C vssd1 vssd1 vccd1 vccd1 _09402_/X sky130_fd_sc_hd__and3_1
X_06614_ _06614_/A _06614_/B _06614_/C vssd1 vssd1 vccd1 vccd1 _06674_/A sky130_fd_sc_hd__nand3_1
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07594_ _07396_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07594_/X sky130_fd_sc_hd__and2b_1
X_09333_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__nor2_2
XFILLER_61_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ _06545_/A _06520_/X vssd1 vssd1 vccd1 vccd1 _06546_/A sky130_fd_sc_hd__or2b_1
X_09264_ _05844_/A _09262_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09264_/X sky130_fd_sc_hd__mux2_1
X_06476_ _06688_/A _06688_/B vssd1 vssd1 vccd1 vccd1 _06658_/A sky130_fd_sc_hd__or2b_1
X_08215_ _08215_/A vssd1 vssd1 vccd1 vccd1 _10695_/D sky130_fd_sc_hd__clkbuf_1
X_05427_ _07875_/A _05360_/X _05358_/X _10633_/Q _05426_/X vssd1 vssd1 vccd1 vccd1
+ _05427_/X sky130_fd_sc_hd__a221o_1
X_09195_ _10946_/Q _09143_/Y _09194_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09195_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _08146_/A vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__buf_2
XANTENNA__09856__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05358_ _05358_/A _05358_/B vssd1 vssd1 vccd1 vccd1 _05358_/X sky130_fd_sc_hd__and2_1
X_08077_ _10526_/A _08047_/X _08052_/X _08075_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08077_/X sky130_fd_sc_hd__o221a_1
XANTENNA__06055__A2 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05289_ _05279_/A _05454_/A _05400_/A vssd1 vssd1 vccd1 vccd1 _05289_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_136_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07028_ _07028_/A _07028_/B vssd1 vssd1 vccd1 vccd1 _07417_/A sky130_fd_sc_hd__xnor2_2
XFILLER_115_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08979_ _10616_/Q _09020_/B vssd1 vssd1 vccd1 vccd1 _08979_/X sky130_fd_sc_hd__or2_1
XFILLER_76_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08000__A _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10941_ _10962_/CLK _10941_/D vssd1 vssd1 vccd1 vccd1 _10941_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08935__A _08935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10872_ _10958_/CLK _10872_/D vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08670__A _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_53_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10306_ _10959_/Q _10943_/Q vssd1 vssd1 vccd1 vccd1 _10307_/B sky130_fd_sc_hd__and2b_1
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _10225_/A _10228_/Y _10225_/B vssd1 vssd1 vccd1 vccd1 _10237_/Y sky130_fd_sc_hd__o21bai_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10168_ _07394_/X _10167_/X _08517_/X _10882_/Q vssd1 vssd1 vccd1 vccd1 _10882_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10099_ _10100_/A _10100_/B _10100_/C vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__a21o_1
XANTENNA__05534__A _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09006__A _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06330_ _10930_/Q _07112_/A vssd1 vssd1 vccd1 vccd1 _06342_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06365__A _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06261_ _10919_/Q _10902_/Q vssd1 vssd1 vccd1 vccd1 _06262_/B sky130_fd_sc_hd__or2_1
X_08000_ _08000_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08000_/X sky130_fd_sc_hd__or2_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06192_ _10596_/Q vssd1 vssd1 vccd1 vccd1 _06193_/A sky130_fd_sc_hd__inv_2
XFILLER_116_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08982__A1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _09671_/A _10023_/B _09949_/Y _10027_/A vssd1 vssd1 vccd1 vccd1 _09952_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_98_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08902_ _10827_/Q _08902_/B vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__and2_1
XFILLER_112_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09882_ _09882_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__xor2_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07924__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08833_ _08829_/X _08832_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10817_/D sky130_fd_sc_hd__o21a_1
XFILLER_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05976_ input51/X vssd1 vssd1 vccd1 vccd1 _08445_/A sky130_fd_sc_hd__clkbuf_2
X_08764_ _08762_/X _08763_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10809_/D sky130_fd_sc_hd__o21a_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07715_ _09379_/B _07571_/B _07715_/C _07715_/D vssd1 vssd1 vccd1 vccd1 _07715_/X
+ sky130_fd_sc_hd__and4bb_1
X_08695_ _08820_/A vssd1 vssd1 vccd1 vccd1 _08695_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07646_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07577_ _07577_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07579_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06528_ _06785_/A _06540_/A vssd1 vssd1 vccd1 vccd1 _06528_/Y sky130_fd_sc_hd__nand2_1
X_09316_ _09316_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09388_/A sky130_fd_sc_hd__xor2_2
X_09247_ _10821_/Q _09243_/X _09244_/X _09246_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09248_/B sky130_fd_sc_hd__a32o_1
X_06459_ _10977_/Q _06459_/B vssd1 vssd1 vccd1 vccd1 _06670_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09178_ _09113_/A _09177_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09178_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08490__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _08132_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08129_/X sky130_fd_sc_hd__or2_1
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput67 _10835_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[1] sky130_fd_sc_hd__buf_2
Xoutput56 _10834_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[0] sky130_fd_sc_hd__buf_2
XFILLER_122_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput78 _10836_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_103_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10022_ _10022_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10532__A1 _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input16_A io_wbs_m2s_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09150__A1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10924_ _10924_/CLK _10924_/D vssd1 vssd1 vccd1 vccd1 _10924_/Q sky130_fd_sc_hd__dfxtp_1
X_10855_ _10855_/CLK _10855_/D vssd1 vssd1 vccd1 vccd1 _10855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08110__C1 _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10790_/CLK _10786_/D vssd1 vssd1 vccd1 vccd1 _10786_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05830_ _05830_/A vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10170__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05950__A1 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05761_ _05749_/A _10564_/Q _10563_/Q _08282_/A vssd1 vssd1 vccd1 vccd1 _05761_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_48_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07500_ _07504_/B _07535_/A _07504_/A vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__o21ai_2
X_05692_ _05692_/A vssd1 vssd1 vccd1 vccd1 _05693_/A sky130_fd_sc_hd__inv_2
X_08480_ _08483_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08481_/A sky130_fd_sc_hd__and2_1
XFILLER_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07431_ _07562_/A vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07362_ _07363_/B _07363_/C _07361_/Y vssd1 vssd1 vccd1 vccd1 _07410_/A sky130_fd_sc_hd__a21bo_1
XFILLER_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09101_ _10938_/Q _10369_/B _09100_/Y _08968_/A vssd1 vssd1 vccd1 vccd1 _09101_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06313_ _06313_/A _06313_/B vssd1 vssd1 vccd1 vccd1 _06755_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07293_ _07317_/A vssd1 vssd1 vccd1 vccd1 _07309_/C sky130_fd_sc_hd__inv_2
XFILLER_31_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06244_ _10611_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06244_/X sky130_fd_sc_hd__or2_1
X_09032_ _10504_/A _09031_/X _09087_/S vssd1 vssd1 vccd1 vccd1 _09032_/X sky130_fd_sc_hd__mux2_1
XFILLER_116_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06175_ hold5/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10211__B1 _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09934_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__or2_1
XFILLER_131_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10514__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09867_/D vssd1 vssd1 vccd1 vccd1 _10139_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA_input8_A io_wbs_m2s_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08183__A2 _08043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08816_ _10816_/Q _08856_/B vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__xor2_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06194__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09796_ _09372_/C _09733_/B _09372_/B vssd1 vssd1 vccd1 vccd1 _09797_/B sky130_fd_sc_hd__a21o_1
X_05959_ input50/X input48/X vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__and2_4
XFILLER_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08747_ _08759_/A _08747_/B _08778_/A vssd1 vssd1 vccd1 vccd1 _08747_/X sky130_fd_sc_hd__and3b_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08678_/A vssd1 vssd1 vccd1 vccd1 _08698_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07629_ _07662_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07630_/B sky130_fd_sc_hd__nor2_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _10851_/CLK _10640_/D vssd1 vssd1 vccd1 vccd1 _10640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06436__C _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _10865_/CLK _10571_/D vssd1 vssd1 vccd1 vccd1 _10571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09199__A1 _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10005_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10505__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10907_ _10920_/CLK _10907_/D vssd1 vssd1 vccd1 vccd1 _10907_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10838_ _10842_/CLK _10838_/D vssd1 vssd1 vccd1 vccd1 _10838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10769_ _10855_/CLK _10769_/D vssd1 vssd1 vccd1 vccd1 _10769_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07437__A1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07980_ _06182_/X _07965_/X _07979_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10658_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_99_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06931_ _06936_/A _06936_/B _06930_/Y vssd1 vssd1 vccd1 vccd1 _06935_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09650_ _09620_/A _09648_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__a21o_1
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
X_08601_ _10783_/Q _08600_/X _10784_/Q vssd1 vssd1 vccd1 vccd1 _08602_/C sky130_fd_sc_hd__a21o_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06862_ _06862_/A _06862_/B vssd1 vssd1 vccd1 vccd1 _06863_/B sky130_fd_sc_hd__nor2_1
X_05813_ _05813_/A _10574_/Q vssd1 vssd1 vccd1 vccd1 _05813_/X sky130_fd_sc_hd__xor2_1
XANTENNA__05923__A1 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09581_ _09638_/C _09703_/A vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__nor2_1
X_06793_ _06833_/A _06793_/B vssd1 vssd1 vccd1 vccd1 _06794_/B sky130_fd_sc_hd__and2_1
X_05744_ _08218_/A vssd1 vssd1 vccd1 vccd1 _05744_/Y sky130_fd_sc_hd__inv_2
X_08532_ _08531_/X _08547_/A _10767_/Q vssd1 vssd1 vccd1 vccd1 _08533_/B sky130_fd_sc_hd__mux2_1
XFILLER_70_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08463_ _10775_/Q hold1/A _08473_/S vssd1 vssd1 vccd1 vccd1 _08464_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10985__D _10985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05675_ _08277_/B _05596_/X _05593_/X _08277_/A _05674_/X vssd1 vssd1 vccd1 vccd1
+ _05675_/X sky130_fd_sc_hd__o221a_1
XFILLER_63_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ _07414_/A _07051_/A vssd1 vssd1 vccd1 vccd1 _07430_/A sky130_fd_sc_hd__or2b_1
XFILLER_35_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08394_ _08394_/A vssd1 vssd1 vccd1 vccd1 _08394_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07345_ _07345_/A _07345_/B vssd1 vssd1 vccd1 vccd1 _07488_/A sky130_fd_sc_hd__xor2_1
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_07276_ _07318_/B _07324_/A _07318_/A vssd1 vssd1 vccd1 vccd1 _07319_/A sky130_fd_sc_hd__a21oi_2
X_06227_ _10604_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06227_/X sky130_fd_sc_hd__or2_1
X_09015_ _10502_/A _09012_/X _09087_/S vssd1 vssd1 vccd1 vccd1 _09015_/X sky130_fd_sc_hd__mux2_1
XFILLER_132_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06158_ _06204_/B vssd1 vssd1 vccd1 vccd1 _06158_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06089_ _06089_/A _06089_/B _06089_/C _06089_/D vssd1 vssd1 vccd1 vccd1 _06089_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_105_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09917_ _09855_/A _09855_/B _09852_/A vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__a21o_1
XFILLER_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09848_ _09848_/A _09848_/B _09848_/C vssd1 vssd1 vccd1 vccd1 _09901_/B sky130_fd_sc_hd__and3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08561__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09787_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09104__A _09104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10623_ _10803_/CLK _10623_/D vssd1 vssd1 vccd1 vccd1 _10623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ _10695_/CLK _10554_/D vssd1 vssd1 vccd1 vccd1 _10554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10485_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 _10985_/CLK sky130_fd_sc_hd__clkbuf_2
XANTENNA__10432__B _10432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05460_ _07871_/A _05460_/B _05460_/C _05460_/D vssd1 vssd1 vccd1 vccd1 _05460_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05391_ _06038_/A _05391_/B vssd1 vssd1 vccd1 vccd1 _05392_/B sky130_fd_sc_hd__and2_1
XFILLER_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07130_ _07134_/A _07133_/A _07133_/B _07123_/B _07144_/A vssd1 vssd1 vccd1 vccd1
+ _07132_/A sky130_fd_sc_hd__o32ai_4
X_07061_ _07061_/A _07061_/B vssd1 vssd1 vccd1 vccd1 _07164_/B sky130_fd_sc_hd__xnor2_4
XFILLER_126_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06012_ _06011_/X _05993_/S _05977_/X vssd1 vssd1 vccd1 vccd1 _06012_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09032__A0 _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07963_ _07963_/A vssd1 vssd1 vccd1 vccd1 _10655_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09335__A1 _09316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07894_ _10605_/Q _07888_/X _07892_/X _07893_/Y vssd1 vssd1 vccd1 vccd1 _07895_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09702_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__xor2_1
X_06914_ _06914_/A _06914_/B vssd1 vssd1 vccd1 vccd1 _06939_/A sky130_fd_sc_hd__xnor2_4
XFILLER_110_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06845_ _06845_/A _07784_/B _06845_/C vssd1 vssd1 vccd1 vccd1 _06847_/A sky130_fd_sc_hd__and3_1
X_09633_ _09631_/A _09631_/B _09631_/C vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__o21a_1
XFILLER_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__xor2_4
XFILLER_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08515_ _08638_/B _08514_/X _08509_/X _10757_/Q vssd1 vssd1 vccd1 vccd1 _10757_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06776_ _06776_/A vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__clkbuf_2
X_05727_ _08130_/A _05739_/B _05549_/A _08117_/A vssd1 vssd1 vccd1 vccd1 _05732_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ _09610_/A _09492_/A _09494_/D _09494_/B vssd1 vssd1 vccd1 vccd1 _09496_/C
+ sky130_fd_sc_hd__a31o_1
X_05658_ _05631_/X _05657_/X _05628_/X _05896_/A vssd1 vssd1 vccd1 vccd1 _05658_/X
+ sky130_fd_sc_hd__a22o_1
X_08446_ _10770_/Q _10733_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08447_/B sky130_fd_sc_hd__mux2_1
X_08377_ _08367_/X _10732_/Q _07865_/X _08376_/X vssd1 vssd1 vccd1 vccd1 _10714_/D
+ sky130_fd_sc_hd__o211a_1
X_05589_ _10703_/Q vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07328_ _07326_/A _07394_/A _07327_/X _07086_/B vssd1 vssd1 vccd1 vccd1 _07328_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_23_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07259_ _07197_/A _07076_/B _07197_/C vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ _10287_/B _10268_/A _10279_/S vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10533__A _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08003__A _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08301__A2 _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__A _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_63_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10909_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10606_ _10830_/CLK _10606_/D vssd1 vssd1 vccd1 vccd1 _10606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10537_ _10537_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10537_/X sky130_fd_sc_hd__or3_1
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10468_ _06195_/X _10459_/X _10467_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10960_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10399_ _10399_/A vssd1 vssd1 vccd1 vccd1 _10399_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06630_ _06630_/A _06630_/B vssd1 vssd1 vccd1 vccd1 _06631_/B sky130_fd_sc_hd__or2_1
XFILLER_92_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_48_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06561_ _06587_/B _06561_/B _06561_/C vssd1 vssd1 vccd1 vccd1 _06573_/C sky130_fd_sc_hd__and3b_1
XFILLER_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09280_ _09280_/A vssd1 vssd1 vccd1 vccd1 _10861_/D sky130_fd_sc_hd__clkbuf_1
X_08300_ _08263_/X _08315_/C _08296_/Y _08299_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08300_/X sky130_fd_sc_hd__o311a_1
X_05512_ _05348_/X _05510_/X _05506_/X _07893_/A vssd1 vssd1 vccd1 vccd1 _10562_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_06492_ _06567_/A _06515_/B vssd1 vssd1 vccd1 vccd1 _06493_/C sky130_fd_sc_hd__nand2_1
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08231_ _08227_/X _08229_/X _08230_/X vssd1 vssd1 vccd1 vccd1 _10697_/D sky130_fd_sc_hd__o21a_1
X_05443_ _10642_/Q _05438_/X _05442_/Y vssd1 vssd1 vccd1 vccd1 _05443_/X sky130_fd_sc_hd__o21ba_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08162_ _08158_/X _08169_/C _08067_/X vssd1 vssd1 vccd1 vccd1 _08162_/Y sky130_fd_sc_hd__o21ai_1
X_05374_ _05374_/A _05374_/B vssd1 vssd1 vccd1 vccd1 _05374_/X sky130_fd_sc_hd__and2_1
X_08093_ _08093_/A vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__06067__B1 _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07113_ _07113_/A _07113_/B vssd1 vssd1 vccd1 vccd1 _07216_/B sky130_fd_sc_hd__xnor2_2
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07927__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ _07044_/A vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05290__A1 _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10166__A2 _10115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _08995_/A vssd1 vssd1 vccd1 vccd1 _08995_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07946_ _07946_/A vssd1 vssd1 vccd1 vccd1 _10650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07877_ _07880_/A _07877_/B vssd1 vssd1 vccd1 vccd1 _10632_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06828_ _06828_/A _06828_/B vssd1 vssd1 vccd1 vccd1 _06882_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09616_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__xnor2_1
XFILLER_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06759_ _06759_/A _06759_/B vssd1 vssd1 vccd1 vccd1 _06779_/B sky130_fd_sc_hd__nor2_1
X_09547_ _09676_/A _09547_/B vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09438_/A _09438_/B _09477_/X vssd1 vssd1 vccd1 vccd1 _09479_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08429_ _10772_/Q _10771_/Q _08547_/B vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__and3_1
XANTENNA__10528__A _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ _10961_/Q _10945_/Q vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__and2b_1
XFILLER_106_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10253_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input46_A io_wbs_m2s_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10184_ _10355_/A vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05820__A _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07747__A _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08780_ _08992_/A vssd1 vssd1 vccd1 vccd1 _08780_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07800_ _06934_/A _06934_/B _07799_/Y vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__a21oi_1
XFILLER_111_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05992_ input45/X _05992_/B vssd1 vssd1 vccd1 vccd1 _05992_/X sky130_fd_sc_hd__xor2_1
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07731_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07662_ _07662_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07663_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09401_ _09437_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09402_/C sky130_fd_sc_hd__or2_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06613_ _06614_/A _06614_/B _06614_/C vssd1 vssd1 vccd1 vccd1 _06674_/C sky130_fd_sc_hd__a21o_1
X_07593_ _07593_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _07596_/A sky130_fd_sc_hd__xnor2_4
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06544_ _06544_/A _06544_/B vssd1 vssd1 vccd1 vccd1 _06622_/B sky130_fd_sc_hd__xnor2_1
X_09332_ _10900_/Q _10884_/Q vssd1 vssd1 vccd1 vccd1 _09333_/B sky130_fd_sc_hd__and2b_1
XFILLER_80_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06826__A _07682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09287_/S sky130_fd_sc_hd__clkbuf_2
X_06475_ _06666_/B _06671_/A _06666_/A vssd1 vssd1 vccd1 vccd1 _06688_/B sky130_fd_sc_hd__a21bo_1
XFILLER_138_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08214_ _08211_/X _08214_/B vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__and2b_1
X_05426_ _07871_/A _05363_/X _05360_/X _10632_/Q _05425_/X vssd1 vssd1 vccd1 vccd1
+ _05426_/X sky130_fd_sc_hd__o221a_1
X_09194_ _10962_/Q _09194_/B vssd1 vssd1 vccd1 vccd1 _09194_/Y sky130_fd_sc_hd__nor2_1
X_08145_ _08145_/A vssd1 vssd1 vccd1 vccd1 _10688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05357_ _06052_/A _05848_/B _10665_/Q vssd1 vssd1 vccd1 vccd1 _05358_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _08038_/X _08074_/X _08075_/Y _08044_/X _06065_/X vssd1 vssd1 vccd1 vccd1
+ _08076_/X sky130_fd_sc_hd__a32o_1
X_05288_ _06065_/A _05283_/Y _05287_/Y vssd1 vssd1 vccd1 vccd1 _05400_/A sky130_fd_sc_hd__a21o_1
XFILLER_107_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07027_ _09344_/B _07007_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _07028_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_130_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08978_ _08978_/A vssd1 vssd1 vccd1 vccd1 _09020_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05905__A _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07929_ _08284_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _10647_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _10955_/CLK _10940_/D vssd1 vssd1 vccd1 vccd1 _10940_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10871_ _10958_/CLK _10871_/D vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09112__A _09112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _10943_/Q _10959_/Q vssd1 vssd1 vccd1 vccd1 _10307_/A sky130_fd_sc_hd__and2b_1
XFILLER_79_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10236_ _10225_/A _10246_/B _10225_/B vssd1 vssd1 vccd1 vccd1 _10236_/X sky130_fd_sc_hd__o21ba_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07951__A0 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08398__A _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10098_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10100_/C sky130_fd_sc_hd__or2_1
XFILLER_47_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06047__A1_N _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08259__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06260_ _10919_/Q _10902_/Q vssd1 vssd1 vccd1 vccd1 _06262_/A sky130_fd_sc_hd__nand2_2
XFILLER_129_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06191_ input19/X vssd1 vssd1 vccd1 vccd1 _06191_/X sky130_fd_sc_hd__buf_4
X_09950_ _09744_/A _09949_/A _09830_/X vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__o21a_1
X_08901_ _09154_/A vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__buf_4
XFILLER_124_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09881_ _09811_/B _09452_/A _09452_/B _10097_/A vssd1 vssd1 vccd1 vccd1 _09882_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08832_ input25/X _08830_/X _08831_/X _10817_/Q vssd1 vssd1 vccd1 vccd1 _08832_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05975_ _05993_/S vssd1 vssd1 vccd1 vccd1 _05975_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08763_ _06182_/X _08728_/X _08729_/X _10809_/Q vssd1 vssd1 vccd1 vccd1 _08763_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07714_ _07713_/B _07713_/Y _07714_/S vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08694_ _08819_/A vssd1 vssd1 vccd1 vccd1 _08694_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07645_ _07645_/A _07645_/B vssd1 vssd1 vccd1 vccd1 _07647_/B sky130_fd_sc_hd__xnor2_2
XFILLER_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07576_ _07576_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06527_ _06527_/A vssd1 vssd1 vccd1 vccd1 _06785_/A sky130_fd_sc_hd__clkbuf_2
X_09315_ _10899_/Q _10883_/Q vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__xor2_4
X_09246_ _05851_/A _09245_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09246_/X sky130_fd_sc_hd__mux2_1
X_06458_ _06458_/A _06458_/B vssd1 vssd1 vccd1 vccd1 _06646_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__05484__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05409_ _10617_/Q vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09177_ _09114_/A _09176_/X _10500_/B vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__o21a_1
X_06389_ _06412_/A _06389_/B vssd1 vssd1 vccd1 vccd1 _06502_/C sky130_fd_sc_hd__xnor2_1
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08128_ _08128_/A vssd1 vssd1 vccd1 vccd1 _10686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ _08059_/A _08082_/D vssd1 vssd1 vccd1 vccd1 _08072_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput57 _10844_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput79 _10864_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[30] sky130_fd_sc_hd__buf_2
Xoutput68 _10854_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_115_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10021_ _10021_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__or2_1
XFILLER_103_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09107__A _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10923_ _10930_/CLK _10923_/D vssd1 vssd1 vccd1 vccd1 _10923_/Q sky130_fd_sc_hd__dfxtp_1
X_10854_ _10854_/CLK _10854_/D vssd1 vssd1 vccd1 vccd1 _10854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _10790_/CLK _10785_/D vssd1 vssd1 vccd1 vccd1 _10785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10219_ _10216_/X _10217_/X _10329_/S vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05760_ _08232_/A _10559_/Q _10558_/Q _08228_/A vssd1 vssd1 vccd1 vccd1 _05764_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05691_ _08169_/A vssd1 vssd1 vccd1 vccd1 _05692_/A sky130_fd_sc_hd__buf_2
XFILLER_90_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ _07430_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07361_ _07406_/A _07361_/B vssd1 vssd1 vccd1 vccd1 _07361_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09100_ _10954_/Q _09124_/A vssd1 vssd1 vccd1 vccd1 _09100_/Y sky130_fd_sc_hd__nor2_1
X_06312_ _10926_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _06313_/B sky130_fd_sc_hd__or2_1
XFILLER_31_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08591__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09031_ _10482_/A _09030_/X _09086_/S vssd1 vssd1 vccd1 vccd1 _09031_/X sky130_fd_sc_hd__mux2_1
X_07292_ _07326_/A _07076_/B _07390_/B _07563_/A vssd1 vssd1 vccd1 vccd1 _07298_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06243_ input34/X _06238_/X _06242_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10610_/D
+ sky130_fd_sc_hd__o211a_1
X_06174_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06193_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10211__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07935__A _10432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__xor2_1
XFILLER_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09864_ _09864_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09867_/D sky130_fd_sc_hd__xnor2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08815_ _08815_/A _08815_/B vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__nand2_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09795_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09883_/A sky130_fd_sc_hd__xor2_4
X_08746_ _08743_/Y _08744_/X _08740_/X _08741_/X vssd1 vssd1 vccd1 vccd1 _08747_/B
+ sky130_fd_sc_hd__a211o_1
X_05958_ _10531_/A vssd1 vssd1 vccd1 vccd1 _05958_/X sky130_fd_sc_hd__buf_4
XFILLER_54_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07670__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05889_ _10659_/Q _05891_/A _05886_/B _05886_/A vssd1 vssd1 vccd1 vccd1 _05889_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08670_/X _08675_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10800_/D sky130_fd_sc_hd__o21a_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07628_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _07698_/A sky130_fd_sc_hd__xor2_2
XFILLER_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07559_ _07724_/A _07559_/B vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__or2_1
X_10570_ _10865_/CLK _10570_/D vssd1 vssd1 vccd1 vccd1 _10570_/Q sky130_fd_sc_hd__dfxtp_2
X_09229_ _09229_/A vssd1 vssd1 vccd1 vccd1 _10853_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09199__A2 _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08006__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10004_ _09940_/B _10078_/A _10003_/X vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__o21a_1
XFILLER_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10906_ _10920_/CLK _10906_/D vssd1 vssd1 vccd1 vccd1 _10906_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10837_ _10839_/CLK _10837_/D vssd1 vssd1 vccd1 vccd1 _10837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10768_ _10768_/CLK _10768_/D vssd1 vssd1 vccd1 vccd1 _10768_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09300__A _09300_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10699_ _10707_/CLK _10699_/D vssd1 vssd1 vccd1 vccd1 _10699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10181__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ _06930_/A _06930_/B vssd1 vssd1 vccd1 vccd1 _06930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08600_ _08600_/A vssd1 vssd1 vccd1 vccd1 _08600_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06861_ _06862_/A _06862_/B vssd1 vssd1 vccd1 vccd1 _06863_/A sky130_fd_sc_hd__and2_1
X_05812_ _10649_/Q vssd1 vssd1 vccd1 vccd1 _05813_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09580_ _10970_/Q _09744_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__nand2_1
X_06792_ _06792_/A _06792_/B vssd1 vssd1 vccd1 vccd1 _06793_/B sky130_fd_sc_hd__or2_1
XFILLER_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05743_ _08224_/B vssd1 vssd1 vccd1 vccd1 _08218_/A sky130_fd_sc_hd__clkbuf_2
X_08531_ _08531_/A _08661_/A vssd1 vssd1 vccd1 vccd1 _08531_/X sky130_fd_sc_hd__or2_1
XANTENNA__08322__B1 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05674_ _05598_/X _05599_/X _05596_/X _10701_/Q _05673_/X vssd1 vssd1 vccd1 vccd1
+ _05674_/X sky130_fd_sc_hd__a221o_1
X_08462_ _08462_/A vssd1 vssd1 vccd1 vccd1 _08477_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ _07549_/A _07413_/B vssd1 vssd1 vccd1 vccd1 _07598_/A sky130_fd_sc_hd__and2_1
X_08393_ _08383_/X hold1/X _08380_/X _08392_/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o211a_1
XFILLER_50_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07344_ _07344_/A _07344_/B vssd1 vssd1 vccd1 vccd1 _07345_/A sky130_fd_sc_hd__and2_1
XANTENNA__09210__A _09274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07275_ _07275_/A _07275_/B vssd1 vssd1 vccd1 vccd1 _07318_/A sky130_fd_sc_hd__xnor2_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06226_ _06253_/B vssd1 vssd1 vccd1 vccd1 _06236_/B sky130_fd_sc_hd__clkbuf_1
X_09014_ _09016_/A _10341_/C vssd1 vssd1 vccd1 vccd1 _09087_/S sky130_fd_sc_hd__or2_1
XFILLER_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06157_ _05958_/X _06131_/X _06156_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10588_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09050__B2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__A1 _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06088_ _05778_/Y _10679_/Q _07985_/A _08180_/A _06087_/X vssd1 vssd1 vccd1 vccd1
+ _06089_/D sky130_fd_sc_hd__a221o_1
XFILLER_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09916_ _09916_/A _09916_/B vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__nor2_1
XFILLER_98_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10499__A1 _06124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09847_ _09716_/Y _09780_/X _09781_/Y _09718_/Y vssd1 vssd1 vccd1 vccd1 _09848_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08496__A _08514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ _09851_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__nor2_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _08831_/A vssd1 vssd1 vccd1 vccd1 _08729_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10622_ _10803_/CLK _10622_/D vssd1 vssd1 vccd1 vccd1 _10622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _10694_/CLK _10553_/D vssd1 vssd1 vccd1 vccd1 _10553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10484_ _10484_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10484_/X sky130_fd_sc_hd__or2_1
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09041__A1 _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05390_ _10653_/Q vssd1 vssd1 vccd1 vccd1 _06038_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07060_ _07112_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07061_/B sky130_fd_sc_hd__nand2_1
X_06011_ _06011_/A vssd1 vssd1 vccd1 vccd1 _06011_/X sky130_fd_sc_hd__buf_4
XANTENNA__05841__A1 _08018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_44_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07962_ _08443_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _07963_/A sky130_fd_sc_hd__or2_1
XFILLER_102_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09701_ _09844_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__nand2_1
X_07893_ _07893_/A vssd1 vssd1 vccd1 vccd1 _07893_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06913_ _06913_/A _06923_/B vssd1 vssd1 vccd1 vccd1 _06914_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09335__A2 _09337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09632_ _09757_/A vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__buf_2
X_06844_ _10510_/A _07783_/B _06844_/C vssd1 vssd1 vccd1 vccd1 _06845_/C sky130_fd_sc_hd__and3_1
X_09563_ _09563_/A _09563_/B vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08514_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08514_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06775_ _06775_/A _06776_/A _06775_/C vssd1 vssd1 vccd1 vccd1 _06792_/A sky130_fd_sc_hd__and3_1
XFILLER_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05726_ _05726_/A vssd1 vssd1 vccd1 vccd1 _08117_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09494_ _09610_/A _09494_/B _09696_/A _09494_/D vssd1 vssd1 vccd1 vccd1 _09542_/A
+ sky130_fd_sc_hd__nand4_2
X_05657_ _10687_/Q _05631_/B _05632_/Y _05726_/A _05656_/X vssd1 vssd1 vccd1 vccd1
+ _05657_/X sky130_fd_sc_hd__a221o_1
X_08445_ _08445_/A vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05588_ _05588_/A _05588_/B vssd1 vssd1 vccd1 vccd1 _05588_/X sky130_fd_sc_hd__and2_1
X_08376_ _08381_/A _10748_/Q vssd1 vssd1 vccd1 vccd1 _08376_/X sky130_fd_sc_hd__or2_1
XFILLER_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07327_ _07327_/A vssd1 vssd1 vccd1 vccd1 _07327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07258_ _07258_/A _07258_/B vssd1 vssd1 vccd1 vccd1 _07273_/A sky130_fd_sc_hd__xor2_1
XANTENNA__05832__A1 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06209_ input9/X _10432_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09104_/B sky130_fd_sc_hd__nand3_1
X_07189_ _07197_/A _07587_/B _07188_/C vssd1 vssd1 vccd1 vccd1 _07190_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10169__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05899__A1 _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _10826_/CLK _10605_/D vssd1 vssd1 vccd1 vccd1 _10605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _07729_/A _10522_/A _10535_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10985_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10960_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__or2_1
XANTENNA__08222__C1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05818__A _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _10938_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10398_/X sky130_fd_sc_hd__and2_1
XFILLER_123_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05339__B1 _10671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08864__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06560_ _06587_/A _06587_/B _06587_/C _07676_/A vssd1 vssd1 vccd1 vccd1 _06585_/B
+ sky130_fd_sc_hd__a31o_1
X_05511_ _05346_/X _05510_/X _05506_/X _07889_/A vssd1 vssd1 vccd1 vccd1 _10561_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06491_ _06568_/A vssd1 vssd1 vccd1 vccd1 _06527_/A sky130_fd_sc_hd__clkbuf_2
X_08230_ input24/X _08164_/X _08165_/X _06061_/A _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08230_/X sky130_fd_sc_hd__o221a_1
X_05442_ _05834_/A _05442_/B vssd1 vssd1 vccd1 vccd1 _05442_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08161_ _07979_/A _08306_/B _08159_/X _08173_/B _06011_/X vssd1 vssd1 vccd1 vccd1
+ _08161_/X sky130_fd_sc_hd__o221a_1
X_05373_ _10659_/Q _05373_/B vssd1 vssd1 vccd1 vccd1 _05374_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08092_ _08092_/A vssd1 vssd1 vccd1 vccd1 _08092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07112_ _07112_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07113_/B sky130_fd_sc_hd__nand2_1
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05814__A1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07043_ _07043_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07048_/B sky130_fd_sc_hd__nor2_1
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08104__A _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08764__B1 _08676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ _08994_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _08994_/X sky130_fd_sc_hd__or2_1
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07945_ _07955_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07946_/A sky130_fd_sc_hd__or2_1
XFILLER_75_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07876_ _10600_/Q _07870_/X _07874_/X _07875_/Y vssd1 vssd1 vccd1 vccd1 _07877_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__xor2_1
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06827_ _06844_/C _06856_/C vssd1 vssd1 vccd1 vccd1 _06883_/A sky130_fd_sc_hd__xor2_1
XFILLER_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06758_ _06758_/A _06758_/B _06758_/C _06786_/A vssd1 vssd1 vccd1 vccd1 _06759_/B
+ sky130_fd_sc_hd__and4_1
X_09546_ _09546_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__nand2_2
X_05709_ _08169_/B vssd1 vssd1 vccd1 vccd1 _05709_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ _09436_/A _09477_/B vssd1 vssd1 vccd1 vccd1 _09477_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08428_ _10770_/Q _10769_/Q _10768_/Q _10767_/Q vssd1 vssd1 vccd1 vccd1 _08547_/B
+ sky130_fd_sc_hd__and4_1
X_06689_ _06690_/A _06690_/B vssd1 vssd1 vccd1 vccd1 _06691_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05502__B1 _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08359_ _05528_/A _08349_/X _08358_/Y vssd1 vssd1 vccd1 vccd1 _08359_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _07570_/A _10283_/X _10320_/X _10293_/X vssd1 vssd1 vccd1 vccd1 _10911_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10252_ _10252_/A _10252_/B vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08949__A input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _07028_/A _10181_/X _10177_/X _10893_/Q vssd1 vssd1 vccd1 vccd1 _10893_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_input39_A io_wbs_m2s_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06230__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07853__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10519_ _10537_/B vssd1 vssd1 vccd1 vccd1 _10531_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08210__A2 _08061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05991_ _07899_/A vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__buf_2
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07730_ _07730_/A _07730_/B vssd1 vssd1 vccd1 vccd1 _07731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07661_ _07661_/A _07661_/B vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09400_ _09399_/B _09400_/B vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__and2b_1
X_07592_ _07592_/A _07592_/B vssd1 vssd1 vccd1 vccd1 _07593_/B sky130_fd_sc_hd__nand2_2
X_06612_ _06612_/A _06612_/B vssd1 vssd1 vccd1 vccd1 _06614_/C sky130_fd_sc_hd__nor2_2
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06543_ _06544_/B _06544_/A vssd1 vssd1 vccd1 vccd1 _06624_/A sky130_fd_sc_hd__or2b_1
X_09331_ _10884_/Q _10900_/Q vssd1 vssd1 vccd1 vccd1 _09333_/A sky130_fd_sc_hd__and2b_1
XFILLER_61_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09262_ _08304_/A _07907_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09262_/X sky130_fd_sc_hd__mux2_1
X_06474_ _06474_/A _06474_/B vssd1 vssd1 vccd1 vccd1 _06666_/A sky130_fd_sc_hd__nand2_1
X_08213_ input22/X _08212_/X _08124_/X _08208_/A _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08214_/B sky130_fd_sc_hd__o221a_1
XFILLER_119_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05425_ _05460_/B _05366_/Y _05363_/X _10631_/Q _05424_/X vssd1 vssd1 vccd1 vccd1
+ _05425_/X sky130_fd_sc_hd__a221o_1
X_09193_ _09202_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _10848_/D sky130_fd_sc_hd__nor2_4
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__and2_1
XANTENNA__07938__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05356_ _05363_/A vssd1 vssd1 vccd1 vccd1 _05848_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08075_/Y sky130_fd_sc_hd__xnor2_1
X_05287_ _05401_/A _05406_/A vssd1 vssd1 vccd1 vccd1 _05287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07026_ _07509_/A _07421_/A _07025_/Y vssd1 vssd1 vccd1 vccd1 _07042_/A sky130_fd_sc_hd__a21oi_1
XFILLER_88_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08977_ _09124_/A _09124_/B _09124_/C vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__or3_2
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07928_ hold17/X _07906_/A _05525_/A _07874_/A vssd1 vssd1 vccd1 vccd1 _07929_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07859_ _10878_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _10889_/CLK _10870_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_1
X_09529_ _09568_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _09529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_15_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10832_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10304_ _07028_/A _10283_/X _10303_/Y _10293_/X vssd1 vssd1 vccd1 vccd1 _10909_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10235_ _10233_/X _10235_/B vssd1 vssd1 vccd1 vccd1 _10246_/C sky130_fd_sc_hd__and2b_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07951__A1 _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10166_ _10881_/Q _10115_/X _10165_/Y _10043_/X vssd1 vssd1 vccd1 vccd1 _10881_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06199__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10097_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__and2_1
XFILLER_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06190_ _06187_/X _06183_/X _06189_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10595_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10184__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ _08897_/Y _08898_/X _08899_/X vssd1 vssd1 vccd1 vccd1 _10826_/D sky130_fd_sc_hd__o21a_1
X_09880_ _09880_/A vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__buf_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08831_ _08831_/A vssd1 vssd1 vccd1 vccd1 _08831_/X sky130_fd_sc_hd__clkbuf_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05974_ _06120_/S vssd1 vssd1 vccd1 vccd1 _05993_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08762_ _08804_/A _08804_/B _08760_/X _08761_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08762_/X sky130_fd_sc_hd__o311a_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08693_ _08693_/A _08693_/B vssd1 vssd1 vccd1 vccd1 _08693_/Y sky130_fd_sc_hd__xnor2_1
X_07713_ _07713_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07713_/Y sky130_fd_sc_hd__nand2_1
XFILLER_93_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07644_ _07662_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07645_/B sky130_fd_sc_hd__or2_1
XANTENNA__09213__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07170__A2 _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07575_ _07574_/A _07574_/B _07574_/C vssd1 vssd1 vccd1 vccd1 _07576_/B sky130_fd_sc_hd__a21oi_1
X_06526_ _06541_/C _06512_/B _06511_/A vssd1 vssd1 vccd1 vccd1 _06535_/B sky130_fd_sc_hd__o21a_1
X_09314_ _09314_/A _09314_/B vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09245_ _08278_/A _07896_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09245_/X sky130_fd_sc_hd__mux2_1
X_06457_ _06457_/A _06465_/A vssd1 vssd1 vccd1 vccd1 _06458_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05408_ _10648_/Q vssd1 vssd1 vccd1 vccd1 _05408_/Y sky130_fd_sc_hd__inv_2
X_09176_ _10944_/Q _09143_/Y _09175_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09176_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06388_ _06388_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06389_/B sky130_fd_sc_hd__nand2_1
X_08127_ _08122_/X _08127_/B vssd1 vssd1 vccd1 vccd1 _08128_/A sky130_fd_sc_hd__and2b_1
XFILLER_107_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05339_ _10670_/Q _05854_/A _10671_/Q vssd1 vssd1 vccd1 vccd1 _05340_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10094__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08058_ _08058_/A vssd1 vssd1 vccd1 vccd1 _08058_/X sky130_fd_sc_hd__buf_2
XFILLER_107_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput58 _10845_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[11] sky130_fd_sc_hd__buf_2
XFILLER_89_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07009_ _07030_/C vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput69 _10855_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10020_ _10021_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__nand2_1
XFILLER_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08011__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10922_ _10924_/CLK _10922_/D vssd1 vssd1 vccd1 vccd1 _10922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09123__A _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10853_ _10855_/CLK _10853_/D vssd1 vssd1 vccd1 vccd1 _10853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10791_/CLK _10784_/D vssd1 vssd1 vccd1 vccd1 _10784_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08110__A1 _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10218_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10329_/S sky130_fd_sc_hd__buf_2
XFILLER_121_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10149_ _10023_/A _10023_/B _10095_/A _10098_/A vssd1 vssd1 vccd1 vccd1 _10151_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05690_ _05528_/X _05564_/Y _05689_/X vssd1 vssd1 vccd1 vccd1 _10728_/D sky130_fd_sc_hd__o21ai_4
XANTENNA__08885__C1 _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07360_ _07360_/A _07407_/A vssd1 vssd1 vccd1 vccd1 _07361_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06311_ _10926_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _06313_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08591__B _10253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09030_ _10949_/Q _10432_/C _09008_/A _10933_/Q vssd1 vssd1 vccd1 vccd1 _09030_/X
+ sky130_fd_sc_hd__a22o_1
X_07291_ _07366_/B _07291_/B _07291_/C vssd1 vssd1 vccd1 vccd1 _07369_/B sky130_fd_sc_hd__and3_1
XFILLER_136_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06242_ _10610_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06242_/X sky130_fd_sc_hd__or2_1
XANTENNA__06392__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06173_ _10592_/Q vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__inv_2
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08168__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05736__A _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09208__A _09208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09863_ _09863_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__xnor2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08814_ _08814_/A vssd1 vssd1 vccd1 vccd1 _08814_/X sky130_fd_sc_hd__buf_2
XFILLER_58_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09794_ _09731_/A _09731_/B _09793_/X vssd1 vssd1 vccd1 vccd1 _09795_/B sky130_fd_sc_hd__a21o_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _08740_/X _08741_/X _08743_/Y _08744_/X vssd1 vssd1 vccd1 vccd1 _08759_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05957_ input42/X vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__buf_4
X_05888_ _08180_/A _05888_/B vssd1 vssd1 vccd1 vccd1 _05888_/X sky130_fd_sc_hd__or2_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _08992_/A vssd1 vssd1 vccd1 vccd1 _08676_/X sky130_fd_sc_hd__buf_2
XFILLER_81_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_39_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05471__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07627_ _07715_/D _07627_/B vssd1 vssd1 vccd1 vccd1 _07628_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07558_ _07557_/B _07558_/B vssd1 vssd1 vccd1 vccd1 _07559_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10435__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06509_ _06510_/A _06510_/B vssd1 vssd1 vccd1 vccd1 _06511_/A sky130_fd_sc_hd__nand2_1
X_07489_ _07489_/A _07489_/B vssd1 vssd1 vccd1 vccd1 _07490_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09228_ _09228_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09229_/A sky130_fd_sc_hd__and2_2
X_09159_ _05461_/A _09136_/X _09148_/X _05692_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09159_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _09930_/B _10123_/B _10139_/S _09716_/A vssd1 vssd1 vccd1 vccd1 _10003_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_92_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input21_A io_wbs_m2s_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08331__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905_ _10920_/CLK _10905_/D vssd1 vssd1 vccd1 vccd1 _10905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10836_ _10836_/CLK _10836_/D vssd1 vssd1 vccd1 vccd1 _10836_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10767_ _10833_/CLK _10767_/D vssd1 vssd1 vccd1 vccd1 _10767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10698_ _10700_/CLK _10698_/D vssd1 vssd1 vccd1 vccd1 _10698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06860_ _06860_/A _06860_/B vssd1 vssd1 vccd1 vccd1 _06862_/B sky130_fd_sc_hd__xnor2_1
X_05811_ _05818_/A _05818_/B vssd1 vssd1 vccd1 vccd1 _05907_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06791_ _06792_/A _06792_/B vssd1 vssd1 vccd1 vccd1 _06833_/A sky130_fd_sc_hd__nand2_1
X_05742_ _05742_/A _05742_/B _05742_/C _05741_/Y vssd1 vssd1 vccd1 vccd1 _05788_/C
+ sky130_fd_sc_hd__or4b_1
X_08530_ _10766_/Q _08419_/B _08529_/X vssd1 vssd1 vccd1 vccd1 _10766_/D sky130_fd_sc_hd__a21o_1
XFILLER_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05673_ _08251_/B _05602_/X _05599_/X _08251_/A _05672_/X vssd1 vssd1 vccd1 vccd1
+ _05673_/X sky130_fd_sc_hd__o221a_1
XANTENNA__05291__A _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08461_ _08461_/A vssd1 vssd1 vccd1 vccd1 _10737_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07412_ _07412_/A _07412_/B _07412_/C vssd1 vssd1 vccd1 vccd1 _07413_/B sky130_fd_sc_hd__or3_1
XFILLER_23_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08395_/A _10754_/Q vssd1 vssd1 vccd1 vccd1 _08392_/X sky130_fd_sc_hd__or2_1
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07343_ _07528_/B _07528_/C _07528_/A vssd1 vssd1 vccd1 vccd1 _07529_/A sky130_fd_sc_hd__a21oi_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ _07323_/B _07331_/A _07323_/A vssd1 vssd1 vccd1 vccd1 _07324_/A sky130_fd_sc_hd__a21o_1
XFILLER_129_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06225_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06225_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09013_ _09013_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _10341_/C sky130_fd_sc_hd__or2_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06156_ _06156_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06156_/Y sky130_fd_sc_hd__nand2_1
X_06087_ _08315_/A _08023_/A _05813_/A _05721_/Y vssd1 vssd1 vccd1 vccd1 _06087_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09915_ _09915_/A _09915_/B _09915_/C vssd1 vssd1 vccd1 vccd1 _09916_/B sky130_fd_sc_hd__nor3_1
XFILLER_86_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09846_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__or2_1
XFILLER_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09778_/B sky130_fd_sc_hd__and2_1
X_06989_ _10979_/Q vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _08830_/A vssd1 vssd1 vccd1 vccd1 _08728_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08659_/A vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__buf_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10621_ _10803_/CLK _10621_/D vssd1 vssd1 vccd1 vccd1 _10621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10552_ _10694_/CLK _10552_/D vssd1 vssd1 vccd1 vccd1 _10552_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10423__A2 _10725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10483_ _06143_/X _10475_/X _10482_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10965_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06000__A _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08068__B1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ _10819_/CLK _10819_/D vssd1 vssd1 vccd1 vccd1 _10819_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10457__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06010_ _08236_/A vssd1 vssd1 vccd1 vccd1 _06011_/A sky130_fd_sc_hd__inv_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07766__A _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__A _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07961_ _10537_/A _06050_/X _07983_/A vssd1 vssd1 vccd1 vccd1 _07962_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09700_ _09769_/A _09810_/B _09769_/B _09764_/A vssd1 vssd1 vccd1 vccd1 _09701_/B
+ sky130_fd_sc_hd__a22o_1
X_06912_ _06916_/A _06912_/B vssd1 vssd1 vccd1 vccd1 _06923_/B sky130_fd_sc_hd__xor2_4
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07892_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07892_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08597__A _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06843_ _10513_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _06848_/A sky130_fd_sc_hd__nand2_1
X_09631_ _09631_/A _09631_/B _09631_/C vssd1 vssd1 vccd1 vccd1 _09631_/X sky130_fd_sc_hd__or3_1
XANTENNA__10350__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09562_ _09562_/A _09562_/B _09562_/C vssd1 vssd1 vccd1 vccd1 _09563_/A sky130_fd_sc_hd__nand3_1
X_06774_ _06785_/A _06774_/B vssd1 vssd1 vccd1 vccd1 _06775_/C sky130_fd_sc_hd__and2_1
X_05725_ _10548_/Q vssd1 vssd1 vccd1 vccd1 _05739_/B sky130_fd_sc_hd__inv_2
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08513_ _10794_/Q vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09493_ _09454_/A _09454_/B _09390_/A vssd1 vssd1 vccd1 vccd1 _09494_/D sky130_fd_sc_hd__a21o_1
X_05656_ _06037_/A _05636_/Y _05632_/Y _10686_/Q _05655_/X vssd1 vssd1 vccd1 vccd1
+ _05656_/X sky130_fd_sc_hd__o221a_1
X_08444_ _08444_/A vssd1 vssd1 vccd1 vccd1 _10732_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__06845__A _06845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05587_ _10564_/Q _05593_/A _10565_/Q vssd1 vssd1 vccd1 vccd1 _05588_/B sky130_fd_sc_hd__o21ai_1
X_08375_ _08367_/X _10731_/Q _07865_/X _08374_/X vssd1 vssd1 vccd1 vccd1 _10713_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07326_ _07326_/A vssd1 vssd1 vccd1 vccd1 _07562_/A sky130_fd_sc_hd__buf_2
XFILLER_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07257_ _07275_/A _07275_/B vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__nor2_1
XFILLER_133_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06208_ _10341_/A vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__buf_4
X_07188_ _07188_/A _07188_/B _07188_/C vssd1 vssd1 vccd1 vccd1 _07190_/A sky130_fd_sc_hd__and3_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06139_ _10585_/Q vssd1 vssd1 vccd1 vccd1 _06140_/A sky130_fd_sc_hd__inv_2
XFILLER_78_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _09829_/A _10023_/A vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__or2_1
XFILLER_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09131__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _10669_/CLK _10604_/D vssd1 vssd1 vccd1 vccd1 _10604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10535_ _10535_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10535_/X sky130_fd_sc_hd__or3_1
XFILLER_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10466_ _06191_/X _10459_/X _10465_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10959_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10397_ _10389_/X _10718_/Q _10394_/X _10396_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10937_/D sky130_fd_sc_hd__o221a_1
XFILLER_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output52_A _10581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09306__A _09306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05510_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05510_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06490_ _10974_/Q vssd1 vssd1 vccd1 vccd1 _06568_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05441_ _10673_/Q _05844_/B _08318_/A vssd1 vssd1 vccd1 vccd1 _05442_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08160_ _08160_/A _08160_/B vssd1 vssd1 vccd1 vccd1 _08173_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05372_ _10628_/Q vssd1 vssd1 vccd1 vccd1 _05460_/D sky130_fd_sc_hd__dlymetal6s2s_1
X_07111_ _07150_/A vssd1 vssd1 vccd1 vccd1 _07135_/A sky130_fd_sc_hd__inv_2
X_08091_ _08091_/A vssd1 vssd1 vccd1 vccd1 _10683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_134_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07042_ _07042_/A _07042_/B vssd1 vssd1 vccd1 vccd1 _07043_/B sky130_fd_sc_hd__nor2_1
XFILLER_115_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08993_ _08970_/X _08983_/X _08991_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10834_/D
+ sky130_fd_sc_hd__o31a_2
XFILLER_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07944_ input38/X _06065_/X _07964_/A vssd1 vssd1 vccd1 vccd1 _07945_/B sky130_fd_sc_hd__mux2_1
X_07875_ _07875_/A vssd1 vssd1 vccd1 vccd1 _07875_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_18_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06826_ _07682_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _06856_/C sky130_fd_sc_hd__nand2_2
X_09614_ _09656_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06757_ _06758_/A _06758_/C _06786_/A _06769_/A vssd1 vssd1 vccd1 vccd1 _06759_/A
+ sky130_fd_sc_hd__a22oi_1
X_09545_ _09617_/B _09545_/B vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__xor2_2
XFILLER_36_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05708_ _05708_/A _05708_/B vssd1 vssd1 vccd1 vccd1 _05708_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ _09476_/A _09476_/B vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__nand2_1
X_06688_ _06688_/A _06688_/B vssd1 vssd1 vccd1 vccd1 _06690_/B sky130_fd_sc_hd__xnor2_1
X_05639_ _10682_/Q vssd1 vssd1 vccd1 vccd1 _05719_/A sky130_fd_sc_hd__clkbuf_2
X_08427_ _10782_/Q _10781_/Q _10780_/Q _10779_/Q vssd1 vssd1 vccd1 vccd1 _08432_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10097__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08358_ _05528_/A _08349_/X _08092_/A vssd1 vssd1 vccd1 vccd1 _08358_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08289_ _08289_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07309_ _07309_/A _07309_/B _07309_/C vssd1 vssd1 vccd1 vccd1 _07310_/B sky130_fd_sc_hd__and3_1
XFILLER_20_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10320_ _10320_/A _10320_/B vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__xor2_1
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10251_ _10249_/Y _10250_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _10252_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10182_ _07008_/A _10181_/X _10177_/X _10892_/Q vssd1 vssd1 vccd1 vccd1 _10892_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08030__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10518_ _10537_/B _10518_/B vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10449_ _05982_/A _10446_/X _10448_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10952_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05990_ _08462_/A vssd1 vssd1 vccd1 vccd1 _07899_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_85_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10470__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09171__A1 _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ _07668_/A _07667_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07661_/B sky130_fd_sc_hd__o21ai_1
XFILLER_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07591_ _09420_/A _07475_/B _07475_/C vssd1 vssd1 vccd1 vccd1 _07592_/B sky130_fd_sc_hd__o21ai_1
XFILLER_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06611_ _06856_/A _06522_/B _06513_/D _06769_/A vssd1 vssd1 vccd1 vccd1 _06612_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09330_ _10965_/Q _09536_/B vssd1 vssd1 vccd1 vccd1 _09451_/B sky130_fd_sc_hd__nand2_1
X_06542_ _06542_/A _06542_/B vssd1 vssd1 vccd1 vccd1 _06544_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09261_ _10441_/A vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08212_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08212_/X sky130_fd_sc_hd__buf_2
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06473_ _06670_/A _06670_/B vssd1 vssd1 vccd1 vccd1 _06671_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05424_ _05460_/C _05369_/Y _05366_/Y _10630_/Q _05423_/X vssd1 vssd1 vccd1 vccd1
+ _05424_/X sky130_fd_sc_hd__o221a_1
X_09192_ _09112_/A _09188_/Y _09191_/X vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08143_ input46/X _08086_/X _08109_/X _06035_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08144_/B sky130_fd_sc_hd__o221a_1
X_05355_ _10664_/Q vssd1 vssd1 vccd1 vccd1 _06052_/A sky130_fd_sc_hd__clkbuf_2
X_08074_ _08074_/A vssd1 vssd1 vccd1 vccd1 _08074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05286_ _10649_/Q _05286_/B vssd1 vssd1 vccd1 vccd1 _05406_/A sky130_fd_sc_hd__nor2_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ _07044_/A _07039_/C vssd1 vssd1 vccd1 vccd1 _07025_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_130_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05474__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08976_ _08976_/A vssd1 vssd1 vccd1 vccd1 _08976_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07927_ _08284_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _10646_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06289__B _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _07848_/X _05461_/A _07844_/X _07857_/Y vssd1 vssd1 vccd1 vccd1 _10627_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08785__A _08819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05723__A1 _05721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06809_ _10911_/Q vssd1 vssd1 vccd1 vccd1 _07570_/A sky130_fd_sc_hd__clkbuf_4
X_07789_ _07789_/A _07789_/B vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__nand2_1
XFILLER_44_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05723__B2 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ _09479_/A _09479_/B _09476_/A vssd1 vssd1 vccd1 vccd1 _09529_/B sky130_fd_sc_hd__o21ai_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08122__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08009__B _08021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09459_ _09458_/B _09458_/C _09458_/A vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__a21o_1
XFILLER_138_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10303_ _10303_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10303_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10234_ _10936_/Q _10952_/Q vssd1 vssd1 vccd1 vccd1 _10235_/B sky130_fd_sc_hd__or2b_1
XANTENNA_input51_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10165_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10165_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_120_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10096_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__nor2_1
XFILLER_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08695__A _08820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08830_/A vssd1 vssd1 vccd1 vccd1 _08830_/X sky130_fd_sc_hd__clkbuf_2
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05294__A _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05973_ _10432_/B _08981_/A vssd1 vssd1 vccd1 vccd1 _06120_/S sky130_fd_sc_hd__nand2_2
X_08761_ _08804_/B _08760_/X _08804_/A vssd1 vssd1 vccd1 vccd1 _08761_/Y sky130_fd_sc_hd__o21ai_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08692_ _08679_/X _08692_/B vssd1 vssd1 vccd1 vccd1 _08693_/B sky130_fd_sc_hd__and2b_1
X_07712_ _07601_/A _07601_/B _07711_/X vssd1 vssd1 vccd1 vccd1 _07757_/A sky130_fd_sc_hd__o21ba_1
XFILLER_38_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07643_ _07643_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07647_/A sky130_fd_sc_hd__xnor2_1
XFILLER_80_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09314_/B sky130_fd_sc_hd__nor2_1
X_07574_ _07574_/A _07574_/B _07574_/C vssd1 vssd1 vccd1 vccd1 _07576_/A sky130_fd_sc_hd__and3_1
X_06525_ _06620_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _06621_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09244_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06456_ _06456_/A _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06465_/A sky130_fd_sc_hd__and3_1
XFILLER_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05407_ _10617_/Q _05480_/A vssd1 vssd1 vccd1 vccd1 _05407_/X sky130_fd_sc_hd__or2_1
X_09175_ _10960_/Q _09194_/B vssd1 vssd1 vccd1 vccd1 _09175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08126_ _10535_/A _08123_/X _08124_/X _08117_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08127_/B sky130_fd_sc_hd__o221a_1
XFILLER_119_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10375__A _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06387_ _06387_/A _06387_/B vssd1 vssd1 vccd1 vccd1 _06412_/B sky130_fd_sc_hd__or2_1
X_05338_ _10639_/Q vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_35_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05269_ _10679_/Q vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__clkinv_4
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08057_ _08352_/B vssd1 vssd1 vccd1 vccd1 _08058_/A sky130_fd_sc_hd__buf_2
XFILLER_89_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07008_ _07008_/A _07008_/B vssd1 vssd1 vccd1 vccd1 _07030_/C sky130_fd_sc_hd__xnor2_2
XFILLER_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput59 _10846_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[12] sky130_fd_sc_hd__buf_2
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08959_ _09736_/B vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10921_ _10924_/CLK _10921_/D vssd1 vssd1 vccd1 vccd1 _10921_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10852_ _10852_/CLK _10852_/D vssd1 vssd1 vccd1 vccd1 _10852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10797_/CLK _10783_/D vssd1 vssd1 vccd1 vccd1 _10783_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08110__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10217_ _10202_/X _10206_/Y _10203_/X vssd1 vssd1 vccd1 vccd1 _10217_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__07385__B1 _09304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10148_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10152_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10079_ _10079_/A _10079_/B vssd1 vssd1 vccd1 vccd1 _10081_/C sky130_fd_sc_hd__xnor2_1
XFILLER_48_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08334__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10444__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06310_ _06730_/A _06730_/B _06730_/C _06731_/B vssd1 vssd1 vccd1 vccd1 _06734_/B
+ sky130_fd_sc_hd__a31o_2
X_07290_ _07287_/A _07287_/B _07289_/X vssd1 vssd1 vccd1 vccd1 _07291_/C sky130_fd_sc_hd__a21bo_1
X_06241_ input33/X _06238_/X _06240_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10609_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_clock _10985_/CLK vssd1 vssd1 vccd1 vccd1 _10848_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06172_ input46/X vssd1 vssd1 vccd1 vccd1 _06172_/X sky130_fd_sc_hd__buf_4
XANTENNA__09062__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07612__A1 _07539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10978_/CLK sky130_fd_sc_hd__clkbuf_16
X_09931_ _09931_/A _10139_/S vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__nand2_1
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09862_ _09346_/B _09797_/B _09861_/X vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__o21a_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08813_ _08810_/X _08812_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10815_/D sky130_fd_sc_hd__a21oi_1
X_09793_ _09730_/B _09793_/B vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__and2b_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05956_ _05956_/A vssd1 vssd1 vccd1 vccd1 _05956_/X sky130_fd_sc_hd__clkbuf_1
X_08744_ _10807_/Q _08744_/B vssd1 vssd1 vccd1 vccd1 _08744_/X sky130_fd_sc_hd__or2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05887_ _07985_/A _05886_/Y _05883_/X vssd1 vssd1 vccd1 vccd1 _05888_/B sky130_fd_sc_hd__o21a_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08675_ _06008_/A _08672_/X _08674_/X _10800_/Q vssd1 vssd1 vccd1 vccd1 _08675_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10768_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07626_ _07700_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__xor2_2
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07557_ _07558_/B _07557_/B vssd1 vssd1 vccd1 vccd1 _07724_/A sky130_fd_sc_hd__and2b_1
XFILLER_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06508_ _06519_/A _06508_/B vssd1 vssd1 vccd1 vccd1 _06510_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_29_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10811_/CLK sky130_fd_sc_hd__clkbuf_16
X_07488_ _07488_/A _07488_/B _07529_/A vssd1 vssd1 vccd1 vccd1 _07489_/B sky130_fd_sc_hd__or3_1
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09227_ _10818_/Q _09210_/X _09212_/X _09226_/X _09203_/X vssd1 vssd1 vccd1 vccd1
+ _09228_/B sky130_fd_sc_hd__a32o_1
X_06439_ _10975_/Q _06561_/C _06440_/A _06461_/B vssd1 vssd1 vccd1 vccd1 _06442_/A
+ sky130_fd_sc_hd__a22o_1
X_09158_ _09113_/X _09157_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09158_/Y sky130_fd_sc_hd__o21ai_1
X_08109_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08109_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09089_ _09081_/X _09088_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10840_/D sky130_fd_sc_hd__o21a_4
XFILLER_135_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08564__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _10484_/A _10139_/S vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__nand2_1
XFILLER_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09108__B2 _10719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input14_A io_wbs_m2s_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10904_ _10924_/CLK _10904_/D vssd1 vssd1 vccd1 vccd1 _10904_/Q sky130_fd_sc_hd__dfxtp_1
X_10835_ _10839_/CLK _10835_/D vssd1 vssd1 vccd1 vccd1 _10835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09292__A0 _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10766_ _10935_/CLK _10766_/D vssd1 vssd1 vccd1 vccd1 _10766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10697_ _10710_/CLK _10697_/D vssd1 vssd1 vccd1 vccd1 _10697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05810_ _10652_/Q vssd1 vssd1 vccd1 vccd1 _05905_/A sky130_fd_sc_hd__buf_2
XANTENNA__08307__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06790_ _06772_/A _06762_/A _07773_/B _06856_/A vssd1 vssd1 vccd1 vccd1 _06792_/B
+ sky130_fd_sc_hd__o211a_1
X_05741_ _08059_/A _05741_/B vssd1 vssd1 vccd1 vccd1 _05741_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08322__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05672_ _10699_/Q _05602_/X _05605_/X _05671_/X vssd1 vssd1 vccd1 vccd1 _05672_/X
+ sky130_fd_sc_hd__a22o_1
X_08460_ _08460_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_2_0_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08391_ _08383_/X _10737_/Q _08380_/X _08390_/X vssd1 vssd1 vccd1 vccd1 _10719_/D
+ sky130_fd_sc_hd__o211a_1
X_07411_ _07412_/B _07412_/C _07412_/A vssd1 vssd1 vccd1 vccd1 _07549_/A sky130_fd_sc_hd__o21ai_1
X_07342_ _07488_/B _07342_/B vssd1 vssd1 vccd1 vccd1 _07528_/A sky130_fd_sc_hd__or2_1
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07273_ _07273_/A _07273_/B vssd1 vssd1 vccd1 vccd1 _07323_/A sky130_fd_sc_hd__xnor2_1
X_06224_ input26/X _06207_/X _06223_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10603_/D
+ sky130_fd_sc_hd__o211a_1
X_09012_ _10480_/A _09009_/X _09086_/S vssd1 vssd1 vccd1 vccd1 _09012_/X sky130_fd_sc_hd__mux2_1
XFILLER_117_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06155_ _10588_/Q vssd1 vssd1 vccd1 vccd1 _06156_/A sky130_fd_sc_hd__inv_2
XFILLER_132_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06086_ _08093_/A _05291_/A _06065_/X _06066_/Y _06085_/X vssd1 vssd1 vccd1 vccd1
+ _06089_/C sky130_fd_sc_hd__a221o_1
XFILLER_117_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09219__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _09915_/A _09915_/B _09915_/C vssd1 vssd1 vccd1 vccd1 _09916_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07962__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09845_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09901_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input6_A io_wbs_m2s_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09776_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06988_ _07563_/A _07433_/A vssd1 vssd1 vccd1 vccd1 _07562_/C sky130_fd_sc_hd__nand2_1
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05939_ _05771_/A _05841_/X _05940_/B _08315_/B _05938_/X vssd1 vssd1 vccd1 vccd1
+ _05939_/X sky130_fd_sc_hd__a221o_1
X_08727_ _08740_/A _08724_/X _08740_/B _08726_/Y _08658_/X vssd1 vssd1 vccd1 vccd1
+ _08727_/X sky130_fd_sc_hd__o311a_1
XFILLER_85_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08849__B1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08778_/A vssd1 vssd1 vccd1 vccd1 _08658_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _07609_/A _07609_/B vssd1 vssd1 vccd1 vccd1 _07706_/B sky130_fd_sc_hd__xnor2_4
X_08589_ _10782_/Q _08586_/B _08588_/Y vssd1 vssd1 vccd1 vccd1 _10782_/D sky130_fd_sc_hd__o21a_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08077__A1 _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _10652_/CLK _10620_/D vssd1 vssd1 vccd1 vccd1 _10620_/Q sky130_fd_sc_hd__dfxtp_1
X_10551_ _10694_/CLK _10551_/D vssd1 vssd1 vccd1 vccd1 _10551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10482_ _10482_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10482_/X sky130_fd_sc_hd__or2_1
XFILLER_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08001__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06012__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_4_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08208__A _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10818_ _10826_/CLK _10818_/D vssd1 vssd1 vccd1 vccd1 _10818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06079__B1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10749_ _10791_/CLK _10749_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10354__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ _07960_/A vssd1 vssd1 vccd1 vccd1 _10654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06911_ _06748_/X _06771_/B _06910_/X vssd1 vssd1 vccd1 vccd1 _06913_/A sky130_fd_sc_hd__a21bo_2
XFILLER_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07891_ _07898_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _10636_/D sky130_fd_sc_hd__nor2_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09630_ _09686_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09631_/C sky130_fd_sc_hd__nor2_1
X_06842_ _06842_/A vssd1 vssd1 vccd1 vccd1 _07776_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09561_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__xnor2_4
X_06773_ _06900_/A _06842_/A _06773_/C vssd1 vssd1 vccd1 vccd1 _06902_/A sky130_fd_sc_hd__and3_2
XFILLER_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05724_ _10687_/Q vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__clkbuf_2
X_08512_ _10793_/Q _08506_/X _08509_/X _10756_/Q vssd1 vssd1 vccd1 vccd1 _10756_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09492_ _09492_/A vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05655_ _10685_/Q _05636_/Y _05637_/Y _08095_/A _05654_/X vssd1 vssd1 vccd1 vccd1
+ _05655_/X sky130_fd_sc_hd__a221o_1
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__or2_1
XFILLER_90_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05586_ _10704_/Q vssd1 vssd1 vccd1 vccd1 _05771_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _08381_/A hold28/X vssd1 vssd1 vccd1 vccd1 _08374_/X sky130_fd_sc_hd__or2_1
XFILLER_23_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07325_ _07338_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07528_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07256_ _07230_/X _07256_/B vssd1 vssd1 vccd1 vccd1 _07275_/B sky130_fd_sc_hd__and2b_1
XFILLER_118_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06207_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06207_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10383__A _10934_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ _07201_/A _07187_/B vssd1 vssd1 vccd1 vccd1 _07188_/C sky130_fd_sc_hd__xnor2_1
XFILLER_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06138_ _06124_/X _06131_/X _06134_/Y _06137_/X vssd1 vssd1 vccd1 vccd1 _10584_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06069_ _06062_/X _06063_/X _06069_/C _06069_/D vssd1 vssd1 vccd1 vccd1 _06070_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09828_ _09977_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__xor2_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ _10826_/CLK _10603_/D vssd1 vssd1 vccd1 vccd1 _10603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10534_ _07727_/A _10522_/X _10533_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10984_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_13_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10465_ _10959_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10465_/X sky130_fd_sc_hd__or2_1
XANTENNA__10293__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08222__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10396_ _10937_/Q _10379_/B _10395_/X vssd1 vssd1 vccd1 vccd1 _10396_/X sky130_fd_sc_hd__a21bo_1
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09306__B _09316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05440_ _10674_/Q vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__buf_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05371_ _07985_/A _05374_/A vssd1 vssd1 vccd1 vccd1 _05371_/Y sky130_fd_sc_hd__xnor2_2
X_07110_ _10983_/Q _07125_/A vssd1 vssd1 vccd1 vccd1 _07150_/A sky130_fd_sc_hd__nand2_1
X_08090_ _08090_/A _08090_/B vssd1 vssd1 vccd1 vccd1 _08091_/A sky130_fd_sc_hd__and2_1
XFILLER_134_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07041_ _07424_/A _07041_/B vssd1 vssd1 vccd1 vccd1 _07048_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08213__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08213__B2 _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09992__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08992_ _08992_/A vssd1 vssd1 vccd1 vccd1 _08992_/X sky130_fd_sc_hd__buf_2
XFILLER_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07943_ _07943_/A vssd1 vssd1 vccd1 vccd1 _10649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07874_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07874_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06825_ _06845_/A _06842_/A vssd1 vssd1 vccd1 vccd1 _06844_/C sky130_fd_sc_hd__nand2_1
X_09613_ _09613_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09614_/B sky130_fd_sc_hd__or3_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06756_ _06756_/A _06806_/B vssd1 vssd1 vccd1 vccd1 _06786_/A sky130_fd_sc_hd__xnor2_2
X_09544_ _09501_/A _09501_/C _09501_/B vssd1 vssd1 vccd1 vccd1 _09545_/B sky130_fd_sc_hd__a21boi_2
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05707_ _05702_/A _10556_/Q _10555_/Q _08196_/A vssd1 vssd1 vccd1 vccd1 _05708_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09232__A _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09475_ _09475_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09476_/B sky130_fd_sc_hd__nand2_1
X_06687_ _06941_/B _06944_/A _06941_/A vssd1 vssd1 vccd1 vccd1 _06942_/A sky130_fd_sc_hd__a21oi_2
XFILLER_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05638_ _10684_/Q vssd1 vssd1 vccd1 vccd1 _08095_/A sky130_fd_sc_hd__clkbuf_2
X_08426_ _10778_/Q _10777_/Q _10776_/Q _10775_/Q vssd1 vssd1 vccd1 vccd1 _08432_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08357_ _08881_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _10710_/D sky130_fd_sc_hd__nor2_1
X_05569_ _10709_/Q vssd1 vssd1 vccd1 vccd1 _08339_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08288_ _08278_/A _08278_/B _08287_/A vssd1 vssd1 vccd1 vccd1 _08288_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07308_ _07308_/A _07319_/A _07308_/C vssd1 vssd1 vccd1 vccd1 _07344_/B sky130_fd_sc_hd__or3_1
X_07239_ _07235_/C _07382_/A _07224_/X vssd1 vssd1 vccd1 vccd1 _07239_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10250_ _10235_/B _10237_/Y _10233_/X vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__a21o_1
XFILLER_133_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10181_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07191__A1 _07229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10517_ _10517_/A vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10448_ _10952_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10448_/X sky130_fd_sc_hd__or2_1
XFILLER_124_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07954__A0 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379_ _10933_/Q _10379_/B vssd1 vssd1 vccd1 vccd1 _10379_/X sky130_fd_sc_hd__and2_1
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09317__A _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06610_ _06758_/B vssd1 vssd1 vccd1 vccd1 _06769_/A sky130_fd_sc_hd__clkbuf_2
X_07590_ _10901_/Q vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__clkinv_2
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10198__A _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06541_ _06785_/A _06719_/C _06541_/C vssd1 vssd1 vccd1 vccd1 _06542_/B sky130_fd_sc_hd__and3_1
X_09260_ _09260_/A vssd1 vssd1 vccd1 vccd1 _10858_/D sky130_fd_sc_hd__clkbuf_4
X_06472_ _06472_/A _06472_/B vssd1 vssd1 vccd1 vccd1 _06670_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08211_ _08114_/X _08224_/C _08207_/Y _08210_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08211_/X sky130_fd_sc_hd__o311a_1
X_05423_ _10629_/Q _05369_/Y _05371_/Y _05460_/D _05422_/X vssd1 vssd1 vccd1 vccd1
+ _05423_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09191_ _10813_/Q _09168_/X _09079_/X _10726_/Q _09190_/X vssd1 vssd1 vccd1 vccd1
+ _09191_/X sky130_fd_sc_hd__a221o_1
X_08142_ _07974_/A _08044_/A _08141_/X vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__a21o_1
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05354_ _10633_/Q vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08073_ _08038_/X _08065_/B _08072_/Y _06033_/X vssd1 vssd1 vccd1 vccd1 _08073_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05285_ _10573_/Q vssd1 vssd1 vccd1 vccd1 _05286_/B sky130_fd_sc_hd__inv_2
XFILLER_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07024_ _07169_/A vssd1 vssd1 vccd1 vccd1 _07044_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08975_ _08995_/A vssd1 vssd1 vccd1 vccd1 _08976_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07926_ hold25/X _07906_/A _07910_/X _07925_/Y vssd1 vssd1 vccd1 vccd1 _07927_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07857_ _06189_/A _07849_/X _07850_/X _07856_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ _07857_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06808_ _07670_/A _06853_/A vssd1 vssd1 vccd1 vccd1 _06814_/A sky130_fd_sc_hd__nand2_1
X_07788_ _06741_/A _06833_/A _06833_/B _06834_/B vssd1 vssd1 vccd1 vccd1 _07789_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_31_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05490__A _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09527_ _09527_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__xnor2_1
X_06739_ _06758_/C vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09458_ _09458_/A _09458_/B _09458_/C vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__nand3_1
X_08409_ _08397_/X _10744_/Q _08992_/A _08408_/X vssd1 vssd1 vccd1 vccd1 _10726_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09389_ _10964_/Q _09396_/A _09411_/A vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__and3_1
XFILLER_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10232__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08025__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _10299_/X _10301_/Y _10329_/S vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10233_ _10952_/Q _10936_/Q vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__and2b_1
XFILLER_133_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10164_ _10164_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input44_A io_wbs_m2s_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07880__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10095_ _10095_/A _10095_/B vssd1 vssd1 vccd1 vccd1 _10097_/B sky130_fd_sc_hd__xor2_1
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05972_ _09107_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__clkbuf_2
X_08760_ _10808_/Q _08748_/X _08928_/B vssd1 vssd1 vccd1 vccd1 _08760_/X sky130_fd_sc_hd__o21a_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08691_ _08689_/Y _08691_/B vssd1 vssd1 vccd1 vccd1 _08693_/A sky130_fd_sc_hd__and2b_1
X_07711_ _07603_/A _07711_/B vssd1 vssd1 vccd1 vccd1 _07711_/X sky130_fd_sc_hd__and2b_1
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07642_ _07527_/B _07648_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07643_/B sky130_fd_sc_hd__o21ai_1
XFILLER_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09312_ _10351_/A vssd1 vssd1 vccd1 vccd1 _09312_/X sky130_fd_sc_hd__buf_2
X_07573_ _07573_/A _07726_/B _07573_/C vssd1 vssd1 vccd1 vccd1 _07574_/C sky130_fd_sc_hd__and3_1
XFILLER_61_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06524_ _06520_/X _06602_/A _06545_/A vssd1 vssd1 vccd1 vccd1 _06620_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ _09274_/A vssd1 vssd1 vccd1 vccd1 _09243_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10462__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06455_ _06468_/A _06450_/B _06478_/A vssd1 vssd1 vccd1 vccd1 _06458_/A sky130_fd_sc_hd__a21o_1
X_05406_ _05406_/A _05406_/B vssd1 vssd1 vccd1 vccd1 _05480_/A sky130_fd_sc_hd__nor2_1
X_09174_ _09202_/A _09174_/B vssd1 vssd1 vccd1 vccd1 _10846_/D sky130_fd_sc_hd__nor2_4
X_06386_ _06386_/A _06386_/B vssd1 vssd1 vccd1 vccd1 _06412_/A sky130_fd_sc_hd__xor2_2
X_08125_ _08201_/A vssd1 vssd1 vccd1 vccd1 _08125_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05337_ _07903_/A _05337_/B vssd1 vssd1 vccd1 vccd1 _05337_/X sky130_fd_sc_hd__or2_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08056_ _08039_/X _08045_/X _08055_/X vssd1 vssd1 vccd1 vccd1 _10680_/D sky130_fd_sc_hd__o21a_1
XANTENNA__07965__A _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07007_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07008_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08958_ _09867_/B vssd1 vssd1 vccd1 vccd1 _09736_/B sky130_fd_sc_hd__buf_2
X_07909_ _07916_/A _07909_/B vssd1 vssd1 vccd1 vccd1 _10641_/D sky130_fd_sc_hd__nor2_1
X_08889_ _08889_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _08889_/X sky130_fd_sc_hd__and2_1
XFILLER_69_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10920_ _10920_/CLK _10920_/D vssd1 vssd1 vccd1 vccd1 _10920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08894__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10851_ _10851_/CLK _10851_/D vssd1 vssd1 vccd1 vccd1 _10851_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10855_/CLK _10782_/D vssd1 vssd1 vccd1 vccd1 _10782_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10453__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08031__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10216_ _10203_/X _10226_/A _10202_/X vssd1 vssd1 vccd1 vccd1 _10216_/X sky130_fd_sc_hd__a21bo_1
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10147_ _10049_/C _10050_/A _09976_/Y vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__a21o_1
XFILLER_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10078_ _10078_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _10079_/B sky130_fd_sc_hd__or2b_1
XFILLER_48_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_1_0_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08885__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10444__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06240_ _10609_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06240_/X sky130_fd_sc_hd__or2_1
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10476__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06171_ _06168_/X _06158_/X _06170_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10591_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08270__C1 _08258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09930_ _09856_/C _09930_/B _09930_/C vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__nand3b_1
XFILLER_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09861_ _10892_/Q _07008_/A vssd1 vssd1 vccd1 vccd1 _09861_/X sky130_fd_sc_hd__or2b_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08812_ input23/X _08672_/X _08674_/X _08815_/A vssd1 vssd1 vccd1 vccd1 _08812_/Y
+ sky130_fd_sc_hd__a22oi_1
X_09792_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__xor2_4
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05955_ _06019_/A _10728_/Q vssd1 vssd1 vccd1 vccd1 _05956_/A sky130_fd_sc_hd__and2_1
X_08743_ _10807_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08743_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08325__B1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05886_ _05886_/A _05886_/B vssd1 vssd1 vccd1 vccd1 _05886_/Y sky130_fd_sc_hd__nor2_1
X_08674_ _08831_/A vssd1 vssd1 vccd1 vccd1 _08674_/X sky130_fd_sc_hd__buf_2
XFILLER_66_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _07625_/A _07625_/B vssd1 vssd1 vccd1 vccd1 _07700_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08089__C1 _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07556_ _07556_/A _07556_/B vssd1 vssd1 vccd1 vccd1 _07557_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10435__A1 _06124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06507_ _06507_/A _06521_/A vssd1 vssd1 vccd1 vccd1 _06508_/B sky130_fd_sc_hd__or2_1
XFILLER_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _08244_/A _09225_/X _09226_/S vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10386__A _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07487_ _07495_/A _07495_/B vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06438_ _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06440_/A sky130_fd_sc_hd__and2_1
X_09157_ _09114_/X _09156_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10199__B1 _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06369_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _06896_/A sky130_fd_sc_hd__and2_1
XFILLER_135_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ _06038_/X _08043_/A _08103_/Y _08038_/A _08107_/X vssd1 vssd1 vccd1 vccd1
+ _08111_/A sky130_fd_sc_hd__a221o_1
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09088_ _07729_/A _09087_/X _10537_/C vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__mux2_1
X_08039_ _08074_/A _08065_/B _05736_/A _08038_/X vssd1 vssd1 vccd1 vccd1 _08039_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10001_ _10076_/A _10001_/B vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__xnor2_1
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10920_/CLK _10903_/D vssd1 vssd1 vccd1 vccd1 _10903_/Q sky130_fd_sc_hd__dfxtp_1
X_10834_ _10987_/CLK _10834_/D vssd1 vssd1 vccd1 vccd1 _10834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10765_ _10935_/CLK _10765_/D vssd1 vssd1 vccd1 vccd1 _10765_/Q sky130_fd_sc_hd__dfxtp_1
X_10696_ _10710_/CLK _10696_/D vssd1 vssd1 vccd1 vccd1 _10696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clock_A _10981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10362__B1 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06030__A1 _10581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05740_ _08082_/C vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05671_ _10698_/Q _05605_/B _05606_/X _08224_/A _05670_/X vssd1 vssd1 vccd1 vccd1
+ _05671_/X sky130_fd_sc_hd__a221o_1
X_08390_ _08395_/A _10753_/Q vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__or2_1
XFILLER_63_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07410_ _07410_/A _07410_/B vssd1 vssd1 vccd1 vccd1 _07412_/A sky130_fd_sc_hd__xor2_1
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07341_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07342_/B sky130_fd_sc_hd__and2_1
XFILLER_137_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07272_ _07330_/A _07335_/A vssd1 vssd1 vccd1 vccd1 _07331_/A sky130_fd_sc_hd__or2_1
XFILLER_129_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06223_ _10603_/Q _06223_/B vssd1 vssd1 vccd1 vccd1 _06223_/X sky130_fd_sc_hd__or2_1
X_09011_ _09194_/B _10432_/C vssd1 vssd1 vccd1 vccd1 _09086_/S sky130_fd_sc_hd__nand2_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06154_ _06147_/X _06131_/X _06151_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10587_/D
+ sky130_fd_sc_hd__o211a_1
X_06085_ _08188_/A _07988_/A vssd1 vssd1 vccd1 vccd1 _06085_/X sky130_fd_sc_hd__xor2_1
XFILLER_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09913_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09915_/C sky130_fd_sc_hd__xor2_1
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09844_ _09844_/A _09844_/B _09844_/C vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__and3_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09775_ _09775_/A _09843_/A vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__xor2_1
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06987_ _07020_/B vssd1 vssd1 vccd1 vccd1 _07433_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05938_ _08285_/A _05853_/X _05841_/X _05771_/A _05937_/X vssd1 vssd1 vccd1 vccd1
+ _05938_/X sky130_fd_sc_hd__o221a_1
X_08726_ _08724_/X _08740_/B _08740_/A vssd1 vssd1 vccd1 vccd1 _08726_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_73_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05869_ _08000_/A _05872_/A vssd1 vssd1 vccd1 vccd1 _05869_/Y sky130_fd_sc_hd__nand2_1
X_08657_ _08686_/A _08659_/A vssd1 vssd1 vccd1 vccd1 _08778_/A sky130_fd_sc_hd__and2_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07608_ _07615_/A _06962_/X _07624_/A vssd1 vssd1 vccd1 vccd1 _07609_/B sky130_fd_sc_hd__a21oi_2
X_08588_ _10782_/Q _08586_/B _08583_/A vssd1 vssd1 vccd1 vccd1 _08588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06088__A1 _05778_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07539_ _07539_/A _07607_/A vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__and2_1
XANTENNA__06088__B2 _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _10657_/CLK _10550_/D vssd1 vssd1 vccd1 vccd1 _10550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09209_ _09037_/A _09209_/B vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__and2b_2
X_10481_ _06008_/X _10475_/X _10480_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10964_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08314__A input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06012__A1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clock _10985_/CLK vssd1 vssd1 vccd1 vccd1 _10852_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05523__B1 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_75_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10797_/CLK sky130_fd_sc_hd__clkbuf_16
X_10817_ _10826_/CLK _10817_/D vssd1 vssd1 vccd1 vccd1 _10817_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06079__B2 _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06009__A _10579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10748_ _10791_/CLK _10748_/D vssd1 vssd1 vccd1 vccd1 _10748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07112__B _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05826__A1 _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10679_ _10710_/CLK _10679_/D vssd1 vssd1 vccd1 vccd1 _10679_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_126_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10855_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06910_ _10502_/A _07776_/B _07783_/B _07780_/C vssd1 vssd1 vccd1 vccd1 _06910_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07890_ _10604_/Q _07888_/X _07874_/X _07889_/Y vssd1 vssd1 vccd1 vccd1 _07891_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10806_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06841_ _06841_/A vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06772_ _06772_/A _06772_/B vssd1 vssd1 vccd1 vccd1 _06773_/C sky130_fd_sc_hd__xnor2_1
X_09560_ _09560_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__xnor2_4
X_05723_ _05721_/Y _10542_/Q _10541_/Q _05736_/A vssd1 vssd1 vccd1 vccd1 _05732_/B
+ sky130_fd_sc_hd__a22o_1
X_08511_ _10792_/Q _08506_/X _08509_/X _10755_/Q vssd1 vssd1 vccd1 vccd1 _10755_/D
+ sky130_fd_sc_hd__a22o_1
X_09491_ _09618_/A _09491_/B vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__nor2_1
X_08442_ _10769_/Q _10732_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08443_/B sky130_fd_sc_hd__mux2_1
XFILLER_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05654_ _10684_/Q _05637_/Y _05649_/X _05718_/A _05653_/X vssd1 vssd1 vccd1 vccd1
+ _05654_/X sky130_fd_sc_hd__o221a_1
X_05585_ _08315_/A vssd1 vssd1 vccd1 vccd1 _05803_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08373_ _08367_/X _10730_/Q _07865_/X _08372_/X vssd1 vssd1 vccd1 vccd1 _10712_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07324_ _07324_/A _07324_/B vssd1 vssd1 vccd1 vccd1 _07338_/B sky130_fd_sc_hd__and2_1
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07255_ _07258_/A _07258_/B _07214_/A vssd1 vssd1 vccd1 vccd1 _07256_/B sky130_fd_sc_hd__o21a_1
X_06206_ input22/X vssd1 vssd1 vccd1 vccd1 _06206_/X sky130_fd_sc_hd__clkbuf_4
X_07186_ _07186_/A _07186_/B _07186_/C vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__and3_1
XFILLER_132_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06137_ _10529_/A vssd1 vssd1 vccd1 vccd1 _06137_/X sky130_fd_sc_hd__clkbuf_2
X_06068_ _05693_/A _07981_/A _06065_/X _06066_/Y _06067_/X vssd1 vssd1 vccd1 vccd1
+ _06069_/D sky130_fd_sc_hd__o221a_1
XANTENNA__07973__A _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08519__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09827_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__and2_1
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09758_ _09755_/X _09757_/X _10875_/Q _09406_/X vssd1 vssd1 vccd1 vccd1 _10875_/D
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08709_ _08709_/A _08725_/A vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__nor2_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09689_ _09689_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__or2b_1
XFILLER_27_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10602_ _10826_/CLK _10602_/D vssd1 vssd1 vccd1 vccd1 _10602_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10533_ _10533_/A _10537_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__or3_1
XFILLER_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10464_ _06187_/X _10459_/X _10463_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10958_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_26_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08979__A _10616_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09322__B _09323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05370_ _10660_/Q vssd1 vssd1 vccd1 vccd1 _07985_/A sky130_fd_sc_hd__clkinv_2
XFILLER_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10484__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07040_ _07416_/A _07433_/A _07434_/A _07567_/A vssd1 vssd1 vccd1 vccd1 _07041_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__08213__A2 _08212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06224__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08991_ _10799_/Q _08985_/X _08988_/X _10712_/Q _08990_/X vssd1 vssd1 vccd1 vccd1
+ _08991_/X sky130_fd_sc_hd__a221o_1
X_07942_ _07955_/A _07942_/B vssd1 vssd1 vccd1 vccd1 _07943_/A sky130_fd_sc_hd__or2_1
XFILLER_110_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07873_ _07880_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _10631_/D sky130_fd_sc_hd__nor2_1
XANTENNA__06202__A input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06824_ _06824_/A _06824_/B vssd1 vssd1 vccd1 vccd1 _06875_/A sky130_fd_sc_hd__or2_1
X_09612_ _09613_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__o21ai_2
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09543_ _09618_/B _09543_/B vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06755_ _06755_/A _06755_/B vssd1 vssd1 vccd1 vccd1 _06806_/B sky130_fd_sc_hd__xnor2_2
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05706_ _05877_/A vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__inv_2
X_09474_ _09475_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__or2_1
X_06686_ _06686_/A _06686_/B vssd1 vssd1 vccd1 vccd1 _06941_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05637_ _10545_/Q _05637_/B vssd1 vssd1 vccd1 vccd1 _05637_/Y sky130_fd_sc_hd__xnor2_1
X_08425_ _08624_/B vssd1 vssd1 vccd1 vccd1 _08661_/A sky130_fd_sc_hd__buf_4
X_08356_ _08348_/Y _08086_/X _08157_/A _08354_/X _08355_/X vssd1 vssd1 vccd1 vccd1
+ _08357_/B sky130_fd_sc_hd__o221a_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05568_ _08351_/A vssd1 vssd1 vccd1 vccd1 _08350_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07307_ _07307_/A _07307_/B vssd1 vssd1 vccd1 vccd1 _07347_/A sky130_fd_sc_hd__xnor2_1
X_08287_ _08287_/A _08295_/C vssd1 vssd1 vccd1 vccd1 _08287_/Y sky130_fd_sc_hd__nor2_1
X_05499_ _05374_/X _05497_/X _05490_/A _05461_/A vssd1 vssd1 vccd1 vccd1 _10552_/D
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10394__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07238_ _07211_/A _07125_/A _07244_/B _07237_/X vssd1 vssd1 vccd1 vccd1 _07264_/B
+ sky130_fd_sc_hd__a31oi_2
X_07169_ _07169_/A _07169_/B vssd1 vssd1 vccd1 vccd1 _07184_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06215__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10180_ _07013_/A _10174_/X _10177_/X _10891_/Q vssd1 vssd1 vccd1 vccd1 _10891_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09142__B _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10516_ _06168_/X _10497_/B _10515_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10978_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10447_ _10472_/B vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07954__A1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10378_ _10365_/X _10713_/Q _10375_/X _10377_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10932_/D sky130_fd_sc_hd__o221a_1
XANTENNA__08502__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06022__A _08837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06540_ _06540_/A vssd1 vssd1 vccd1 vccd1 _06719_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06471_ _06474_/A _06474_/B vssd1 vssd1 vccd1 vccd1 _06666_/B sky130_fd_sc_hd__or2_1
X_08210_ _08218_/B _08061_/A _08208_/Y _08209_/Y _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08210_/X sky130_fd_sc_hd__a311o_1
X_05422_ _10628_/Q _05371_/Y _05374_/X _05461_/A _05421_/X vssd1 vssd1 vccd1 vccd1
+ _05422_/X sky130_fd_sc_hd__o221a_1
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09190_ _08198_/A _09226_/S _09203_/A _09189_/X vssd1 vssd1 vccd1 vccd1 _09190_/X
+ sky130_fd_sc_hd__o211a_1
X_08141_ _08058_/A _08137_/Y _08140_/Y _08113_/A _08096_/A vssd1 vssd1 vccd1 vccd1
+ _08141_/X sky130_fd_sc_hd__a221o_1
X_05353_ _05353_/A _05353_/B vssd1 vssd1 vccd1 vccd1 _05353_/X sky130_fd_sc_hd__and2_1
X_08072_ _08075_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08072_/Y sky130_fd_sc_hd__xnor2_1
X_05284_ _10650_/Q _10574_/Q vssd1 vssd1 vccd1 vccd1 _05401_/A sky130_fd_sc_hd__xor2_1
XFILLER_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07023_ _07222_/A vssd1 vssd1 vccd1 vccd1 _07169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08412__A _10432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08974_ _08974_/A vssd1 vssd1 vccd1 vccd1 _08974_/X sky130_fd_sc_hd__clkbuf_2
X_07925_ _07925_/A vssd1 vssd1 vccd1 vccd1 _07925_/Y sky130_fd_sc_hd__clkinv_2
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07856_ _10877_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09243__A _09274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07787_ _07787_/A _07787_/B vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__xnor2_1
X_06807_ _06818_/A _06817_/B vssd1 vssd1 vccd1 vccd1 _06853_/A sky130_fd_sc_hd__or2_1
XFILLER_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _09625_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__xnor2_2
X_06738_ _06752_/A _06738_/B vssd1 vssd1 vccd1 vccd1 _06758_/C sky130_fd_sc_hd__xnor2_2
XFILLER_43_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08122__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09457_ _09456_/B _09456_/C _09456_/A vssd1 vssd1 vccd1 vccd1 _09458_/C sky130_fd_sc_hd__a21o_1
X_08408_ _08408_/A hold21/X vssd1 vssd1 vccd1 vccd1 _08408_/X sky130_fd_sc_hd__or2_1
XFILLER_52_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06669_ _06686_/A _06686_/B vssd1 vssd1 vccd1 vccd1 _06915_/B sky130_fd_sc_hd__and2_1
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09388_ _09388_/A _09388_/B vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__xnor2_2
X_08339_ _08339_/A _08339_/B _08339_/C vssd1 vssd1 vccd1 vccd1 _08350_/B sky130_fd_sc_hd__and3_1
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08306__B _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10232__A2 _10115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10301_ _10301_/A _10301_/B vssd1 vssd1 vccd1 vccd1 _10301_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10232_ _07056_/A _10115_/X _10231_/X _10043_/X vssd1 vssd1 vccd1 vccd1 _10902_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10163_ _10112_/A _10112_/B _10162_/X vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__a21oi_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input37_A io_wbs_m2s_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09138__B1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10094_ _10097_/A _10025_/B vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__or2b_1
XFILLER_47_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08361__A1 _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09153__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__A_N _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08821__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06017__A _10341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05971_ _08965_/A _09124_/B vssd1 vssd1 vccd1 vccd1 _09107_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _07607_/A _07604_/B _07539_/A vssd1 vssd1 vccd1 vccd1 _07758_/A sky130_fd_sc_hd__o21ai_2
XFILLER_93_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08690_ _10802_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08691_/B sky130_fd_sc_hd__nand2_1
XFILLER_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07641_ _07641_/A _07641_/B vssd1 vssd1 vccd1 vccd1 _07693_/B sky130_fd_sc_hd__xnor2_2
XFILLER_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07572_ _09379_/B _07572_/B vssd1 vssd1 vccd1 vccd1 _07574_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10002__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ _10043_/A _09309_/Y _09326_/A _10192_/A hold16/A vssd1 vssd1 vccd1 vccd1
+ _10866_/D sky130_fd_sc_hd__a32o_1
X_06523_ _06532_/A _06523_/B _06523_/C vssd1 vssd1 vccd1 vccd1 _06545_/A sky130_fd_sc_hd__and3_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09242_ _09242_/A vssd1 vssd1 vccd1 vccd1 _10855_/D sky130_fd_sc_hd__clkbuf_1
X_06454_ _06477_/A _06477_/B vssd1 vssd1 vccd1 vccd1 _06478_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05405_ _05405_/A _05643_/A vssd1 vssd1 vccd1 vccd1 _05406_/B sky130_fd_sc_hd__nor2_1
X_09173_ _09112_/X _09167_/Y _09172_/X vssd1 vssd1 vccd1 vccd1 _09174_/B sky130_fd_sc_hd__a21oi_1
X_06385_ _06305_/A _06274_/B _06374_/B _06303_/A vssd1 vssd1 vccd1 vccd1 _06386_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_135_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08124_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08124_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05336_ _05336_/A _05336_/B vssd1 vssd1 vccd1 vccd1 _05337_/B sky130_fd_sc_hd__and2_1
XFILLER_135_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ _06124_/A _08047_/X _08052_/X _08082_/D _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08055_/X sky130_fd_sc_hd__o221a_1
XFILLER_134_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07006_ _07197_/A vssd1 vssd1 vccd1 vccd1 _07567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07981__A _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08957_ _09610_/B vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__clkbuf_2
X_07908_ _10609_/Q _07906_/X _07892_/X _07907_/Y vssd1 vssd1 vccd1 vccd1 _07909_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08888_ _10825_/Q _08888_/B vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__or2_1
XFILLER_57_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07839_ _06170_/A _07828_/X _07829_/X _07838_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07839_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__10150__A1 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10850_ _10851_/CLK _10850_/D vssd1 vssd1 vccd1 vccd1 _10850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10781_ _10781_/CLK _10781_/D vssd1 vssd1 vccd1 vccd1 _10781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09867_/A _09610_/B _09555_/B _09599_/B vssd1 vssd1 vccd1 vccd1 _09613_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08052__A _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10215_ _10226_/B _10226_/C vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10146_ _10146_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ _10982_/CLK _10979_/D vssd1 vssd1 vccd1 vccd1 _10979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06170_ _06170_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06170_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06970__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_74_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _09735_/A _09735_/B _09859_/Y _09432_/A vssd1 vssd1 vccd1 vccd1 _09864_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_86_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10380__A1 _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08811_ _10815_/Q vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__clkbuf_2
X_09791_ _09711_/B _09727_/B _09711_/A vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__o21bai_4
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05954_ _05954_/A vssd1 vssd1 vccd1 vccd1 _05954_/X sky130_fd_sc_hd__clkbuf_1
X_08742_ _08744_/B vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08673_ _08686_/A _08830_/A vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__nor2_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05885_ _05885_/A vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__buf_2
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10132__A1 _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ _07624_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _07625_/B sky130_fd_sc_hd__nor2_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08089__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07555_ _07732_/A _07555_/B _07713_/B vssd1 vssd1 vccd1 vccd1 _07556_/B sky130_fd_sc_hd__and3_1
X_07486_ _07485_/A _07485_/B _07493_/B _07493_/A vssd1 vssd1 vccd1 vccd1 _07495_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_06506_ _06517_/A _06506_/B vssd1 vssd1 vccd1 vccd1 _06507_/A sky130_fd_sc_hd__nand2_1
X_09225_ _08242_/A _07885_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09225_/X sky130_fd_sc_hd__mux2_1
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06437_ _10975_/Q _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06472_/A sky130_fd_sc_hd__and3_1
XFILLER_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07976__A _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ _10942_/Q _09143_/Y _09155_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09156_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06368_ _06451_/C _06368_/B vssd1 vssd1 vccd1 vccd1 _06895_/B sky130_fd_sc_hd__nor2_2
X_08107_ _08113_/A _08104_/Y _08115_/B _06024_/A vssd1 vssd1 vccd1 vccd1 _08107_/X
+ sky130_fd_sc_hd__a31o_1
X_05319_ _10646_/Q vssd1 vssd1 vccd1 vccd1 _07925_/A sky130_fd_sc_hd__clkbuf_2
X_09087_ _10513_/A _09086_/X _09087_/S vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__mux2_1
X_06299_ _10920_/Q _10903_/Q vssd1 vssd1 vccd1 vccd1 _06304_/B sky130_fd_sc_hd__or2_1
X_08038_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10000_ _09801_/A _09933_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _10001_/B sky130_fd_sc_hd__a21oi_2
XFILLER_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__xnor2_1
XFILLER_57_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10902_ _10920_/CLK _10902_/D vssd1 vssd1 vccd1 vccd1 _10902_/Q sky130_fd_sc_hd__dfxtp_1
X_10833_ _10833_/CLK _10833_/D vssd1 vssd1 vccd1 vccd1 _10833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10764_ _10935_/CLK _10764_/D vssd1 vssd1 vccd1 vccd1 _10764_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10426__A2 _10726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10695_ _10695_/CLK _10695_/D vssd1 vssd1 vccd1 vccd1 _10695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06030__A2 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10129_ _10129_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10251__S _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10114__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05670_ _08224_/B _05610_/X _05606_/X _10697_/Q _05669_/X vssd1 vssd1 vccd1 vccd1
+ _05670_/X sky130_fd_sc_hd__o221a_1
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10487__A _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10417__A2 _10723_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07340_ _07525_/A _07525_/B _07526_/A vssd1 vssd1 vccd1 vccd1 _07528_/C sky130_fd_sc_hd__a21o_1
X_09010_ _09124_/A vssd1 vssd1 vccd1 vccd1 _09194_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07271_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07335_/A sky130_fd_sc_hd__or2_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06222_ input25/X _06207_/X _06220_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10602_/D
+ sky130_fd_sc_hd__o211a_1
X_06153_ _10343_/A vssd1 vssd1 vccd1 vccd1 _06153_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06254__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08794__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06084_ _05291_/A _08093_/A _05766_/Y _05830_/A vssd1 vssd1 vccd1 vccd1 _06089_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09912_ _09842_/A _09842_/B _09841_/A vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__a21oi_2
XFILLER_112_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09843_ _09843_/A _09775_/A vssd1 vssd1 vccd1 vccd1 _09844_/C sky130_fd_sc_hd__or2b_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09771_/B _09773_/X _09705_/B _09708_/A vssd1 vssd1 vccd1 vccd1 _09843_/A
+ sky130_fd_sc_hd__o31a_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _06997_/B _06986_/B vssd1 vssd1 vccd1 vccd1 _07020_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05937_ _08277_/A _05935_/B _05853_/X _08285_/A _05936_/X vssd1 vssd1 vccd1 vccd1
+ _05937_/X sky130_fd_sc_hd__a221o_1
X_08725_ _08725_/A _08725_/B vssd1 vssd1 vccd1 vccd1 _08740_/B sky130_fd_sc_hd__and2_1
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05868_ _10665_/Q vssd1 vssd1 vccd1 vccd1 _08000_/A sky130_fd_sc_hd__buf_2
X_08656_ _10369_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _08659_/A sky130_fd_sc_hd__nand2_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _10781_/Q _08583_/B _08586_/Y vssd1 vssd1 vccd1 vccd1 _10781_/D sky130_fd_sc_hd__o21a_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07607_ _07607_/A _07607_/B vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__nand2_2
X_05799_ _05717_/B _05798_/Y _05708_/A vssd1 vssd1 vccd1 vccd1 _05799_/X sky130_fd_sc_hd__o21a_1
X_07538_ _07606_/A _07606_/B vssd1 vssd1 vccd1 vccd1 _07607_/A sky130_fd_sc_hd__or2_1
XFILLER_50_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06088__A2 _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ _07746_/A _07469_/B vssd1 vssd1 vccd1 vccd1 _07497_/A sky130_fd_sc_hd__xor2_1
XFILLER_108_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ _09208_/A vssd1 vssd1 vccd1 vccd1 _10850_/D sky130_fd_sc_hd__clkbuf_1
X_10480_ _10480_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10480_/X sky130_fd_sc_hd__or2_1
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09139_ _10808_/Q _08985_/X _08988_/X _10721_/Q _09138_/X vssd1 vssd1 vccd1 vccd1
+ _09139_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06115__A _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05954__A _05954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08537__A1 _10291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10798_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_91_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_22_clock_A _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08068__A3 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10816_ _10878_/CLK _10816_/D vssd1 vssd1 vccd1 vccd1 _10816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06079__A2 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10747_ _10791_/CLK _10747_/D vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _10710_/CLK _10678_/D vssd1 vssd1 vccd1 vccd1 _10678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06840_ _07789_/A _06840_/B vssd1 vssd1 vccd1 vccd1 _06864_/A sky130_fd_sc_hd__and2_1
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06771_ _06940_/A _06771_/B vssd1 vssd1 vccd1 vccd1 _06772_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05722_ _05913_/A vssd1 vssd1 vccd1 vccd1 _05736_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08510_ _10791_/Q _08506_/X _08509_/X _10754_/Q vssd1 vssd1 vccd1 vccd1 _10754_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09490_ _09489_/A _09642_/A _09492_/A _09555_/A vssd1 vssd1 vccd1 vccd1 _09491_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__08161__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05653_ _05651_/Y _05652_/X _05649_/X _05718_/A vssd1 vssd1 vccd1 vccd1 _05653_/X
+ sky130_fd_sc_hd__a22o_1
X_08441_ _08476_/S vssd1 vssd1 vccd1 vccd1 _08455_/S sky130_fd_sc_hd__buf_2
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05584_ _10706_/Q vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__buf_2
X_08372_ _08381_/A _10746_/Q vssd1 vssd1 vccd1 vccd1 _08372_/X sky130_fd_sc_hd__or2_1
XFILLER_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07323_ _07323_/A _07323_/B _07331_/A vssd1 vssd1 vccd1 vccd1 _07324_/B sky130_fd_sc_hd__nand3_1
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07254_ _07254_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07258_/B sky130_fd_sc_hd__and2_1
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06205_ _06202_/X _06183_/X _06204_/Y _06200_/X vssd1 vssd1 vccd1 vccd1 _10598_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08415__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__CLK _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ _07185_/A _07185_/B vssd1 vssd1 vccd1 vccd1 _07201_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06136_ _08166_/A vssd1 vssd1 vccd1 vccd1 _10529_/A sky130_fd_sc_hd__buf_2
X_06067_ _05756_/A _08235_/A _05818_/A _08082_/A vssd1 vssd1 vccd1 vccd1 _06067_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07975__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08150__A _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09192__A1 _09112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09826_ _09815_/A _09815_/B _09825_/X vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__a21o_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09757_ _09757_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09757_/X sky130_fd_sc_hd__or2_1
X_06969_ _07007_/A vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__buf_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08708_ _10804_/Q _08732_/B vssd1 vssd1 vccd1 vccd1 _08725_/B sky130_fd_sc_hd__xor2_1
XFILLER_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09688_ _10043_/A _09686_/X _09755_/B _10192_/A _10874_/Q vssd1 vssd1 vccd1 vccd1
+ _10874_/D sky130_fd_sc_hd__a32o_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08638_/B _10793_/Q _08600_/A _08642_/D _10795_/Q vssd1 vssd1 vccd1 vccd1
+ _08640_/B sky130_fd_sc_hd__a41o_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10601_ _10814_/CLK _10601_/D vssd1 vssd1 vccd1 vccd1 _10601_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10532_ _07713_/A _10522_/X _10531_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10983_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10463_ _10958_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10463_/X sky130_fd_sc_hd__or2_1
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10394_ _10535_/A _10394_/B _10394_/C vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__and3_1
XFILLER_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05441__B1 _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09183__A1 _09112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08997__A1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08235__A _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08749__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08990_ _10765_/Q _09037_/A _08990_/C vssd1 vssd1 vccd1 vccd1 _08990_/X sky130_fd_sc_hd__and3_1
XFILLER_114_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07941_ input27/X _05813_/A _07964_/A vssd1 vssd1 vccd1 vccd1 _07942_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07872_ _10599_/Q _07870_/X _07848_/A _07871_/Y vssd1 vssd1 vccd1 vccd1 _07873_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06823_ _06823_/A _06823_/B vssd1 vssd1 vccd1 vccd1 _06824_/B sky130_fd_sc_hd__nor2_1
X_09611_ _09611_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09613_/C sky130_fd_sc_hd__nor2_1
XFILLER_28_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06754_ _06317_/B _06729_/B _06317_/A vssd1 vssd1 vccd1 vccd1 _06755_/B sky130_fd_sc_hd__a21bo_1
X_09542_ _09542_/A _09542_/B _09542_/C vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__and3_1
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05705_ _05704_/Y _05663_/A _10553_/Q _08181_/A vssd1 vssd1 vccd1 vccd1 _05708_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08685__B1 _08676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09473_ _09524_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09475_/B sky130_fd_sc_hd__xnor2_2
X_06685_ _06943_/B _06943_/C _06943_/A vssd1 vssd1 vccd1 vccd1 _06944_/A sky130_fd_sc_hd__a21o_1
X_05636_ _05636_/A _05636_/B vssd1 vssd1 vccd1 vccd1 _05636_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__05499__B1 _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__xnor2_4
X_05567_ _10710_/Q vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__buf_2
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08355_/X sky130_fd_sc_hd__or2_1
X_07306_ _07349_/B _07349_/C _07349_/A vssd1 vssd1 vccd1 vccd1 _07461_/B sky130_fd_sc_hd__o21a_1
X_08286_ _08287_/A _08295_/C vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__and2_1
X_05498_ _05378_/Y _05497_/X _05490_/X _05461_/B vssd1 vssd1 vccd1 vccd1 _10551_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_07237_ _07236_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07237_/X sky130_fd_sc_hd__and2b_1
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07984__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07168_ _07196_/A _07334_/A _07195_/A vssd1 vssd1 vccd1 vccd1 _07192_/B sky130_fd_sc_hd__a21o_1
XFILLER_133_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06119_ _07880_/A _06119_/B vssd1 vssd1 vccd1 vccd1 _10582_/D sky130_fd_sc_hd__nor2_1
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_74_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10790_/CLK sky130_fd_sc_hd__clkbuf_16
X_07099_ _07219_/B vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09809_ _09883_/A _09809_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__xor2_2
XFILLER_86_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_12_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10781_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_27_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10808_/CLK sky130_fd_sc_hd__clkbuf_16
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__or2_1
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10446_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10538__A1 _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10377_ _06008_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10377_/X sky130_fd_sc_hd__a21bo_1
XFILLER_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06470_ _06470_/A _06470_/B vssd1 vssd1 vccd1 vccd1 _06474_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05421_ _05461_/B _05378_/Y _05374_/X _10627_/Q _05420_/X vssd1 vssd1 vccd1 vccd1
+ _05421_/X sky130_fd_sc_hd__a221o_1
X_08140_ _08148_/B _08140_/B vssd1 vssd1 vccd1 vccd1 _08140_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05352_ _10666_/Q _05358_/A vssd1 vssd1 vccd1 vccd1 _05353_/B sky130_fd_sc_hd__nand2_1
X_08071_ _08082_/B vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__clkbuf_2
X_05283_ _10574_/Q vssd1 vssd1 vccd1 vccd1 _05283_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07022_ _10980_/Q vssd1 vssd1 vccd1 vccd1 _07222_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06213__A _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _09211_/A vssd1 vssd1 vccd1 vccd1 _08974_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07924_ _08284_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _10645_/D sky130_fd_sc_hd__nor2_1
XFILLER_102_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_69_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07855_ _07848_/X _05461_/B _07844_/X _07854_/Y vssd1 vssd1 vccd1 vccd1 _10626_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07786_ _07786_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _07787_/B sky130_fd_sc_hd__xnor2_1
X_06806_ _06806_/A _06806_/B vssd1 vssd1 vccd1 vccd1 _06817_/B sky130_fd_sc_hd__or2_1
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09525_ _09626_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__nand2_1
X_06737_ _06745_/B _06746_/A _07675_/A vssd1 vssd1 vccd1 vccd1 _06738_/B sky130_fd_sc_hd__a21o_1
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07979__A _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06668_ _06668_/A _06668_/B vssd1 vssd1 vccd1 vccd1 _06686_/B sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_69_clock_A _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ _09456_/A _09456_/B _09456_/C vssd1 vssd1 vccd1 vccd1 _09458_/B sky130_fd_sc_hd__nand3_1
X_05619_ _05663_/B _05619_/B vssd1 vssd1 vccd1 vccd1 _05619_/X sky130_fd_sc_hd__and2_1
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _09090_/A vssd1 vssd1 vccd1 vccd1 _08992_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06599_ _06599_/A _06599_/B vssd1 vssd1 vccd1 vccd1 _06616_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07698__B _07698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ _09387_/A _09424_/A vssd1 vssd1 vccd1 vccd1 _09388_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08338_ _06033_/X _08334_/X _08336_/Y _08337_/X vssd1 vssd1 vccd1 vccd1 _10708_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _08278_/B _08253_/X _08267_/Y _08268_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08269_/X sky130_fd_sc_hd__a311o_1
XFILLER_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10300_ _10300_/A _10300_/B vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ _10246_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__xor2_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06123__A input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10162_ _10110_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__and2b_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09138__A1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ _10121_/S _10093_/B vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__nor2_2
XFILLER_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05962__A input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09074__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10429_ _10408_/A _10727_/Q _10427_/X _10428_/X _06257_/X vssd1 vssd1 vccd1 vccd1
+ _10946_/D sky130_fd_sc_hd__o221a_1
XFILLER_112_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09129__B2 _10720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05970_ _06126_/D vssd1 vssd1 vccd1 vccd1 _09124_/B sky130_fd_sc_hd__clkbuf_2
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07640_ _07645_/A _07644_/B _07662_/A vssd1 vssd1 vccd1 vccd1 _07641_/B sky130_fd_sc_hd__a21oi_1
XFILLER_53_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ _07678_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07572_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09310_ _09313_/B _09396_/A _09310_/C vssd1 vssd1 vccd1 vccd1 _09326_/A sky130_fd_sc_hd__or3_1
XFILLER_15_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_70_clock_A _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06522_ _06600_/A _06522_/B _06522_/C vssd1 vssd1 vccd1 vccd1 _06602_/A sky130_fd_sc_hd__and3_1
XFILLER_34_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ _09259_/A _09241_/B vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__and2_4
X_06453_ _06453_/A _06453_/B vssd1 vssd1 vccd1 vccd1 _06477_/B sky130_fd_sc_hd__or2_1
XFILLER_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05404_ _10573_/Q vssd1 vssd1 vccd1 vccd1 _05643_/A sky130_fd_sc_hd__clkbuf_2
X_09172_ _08771_/A _09168_/X _09079_/X _10724_/Q _09171_/X vssd1 vssd1 vccd1 vccd1
+ _09172_/X sky130_fd_sc_hd__a221o_1
XANTENNA__06208__A _10341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06384_ _06719_/A vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__buf_4
X_08123_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08123_/X sky130_fd_sc_hd__buf_2
X_05335_ _08298_/A _05340_/A vssd1 vssd1 vccd1 vccd1 _05336_/B sky130_fd_sc_hd__nand2_1
X_08054_ _08175_/A vssd1 vssd1 vccd1 vccd1 _08054_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08812__B1 _08674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ _07188_/A vssd1 vssd1 vccd1 vccd1 _07197_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08040__A1 _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08956_ _09449_/A vssd1 vssd1 vccd1 vccd1 _09610_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_111_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07907_ _07907_/A vssd1 vssd1 vccd1 vccd1 _07907_/Y sky130_fd_sc_hd__clkinv_2
X_08887_ _10825_/Q _08902_/B vssd1 vssd1 vccd1 vccd1 _08889_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07838_ hold9/X _07845_/B vssd1 vssd1 vccd1 vccd1 _07838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10438__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07769_ _07769_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07771_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09508_ _09508_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09599_/B sky130_fd_sc_hd__xor2_2
X_10780_ _10781_/CLK _10780_/D vssd1 vssd1 vccd1 vccd1 _10780_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09438_/A _09438_/B _10351_/A vssd1 vssd1 vccd1 vccd1 _09439_/X sky130_fd_sc_hd__o21a_1
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05957__A input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08031__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10214_ _10214_/A vssd1 vssd1 vccd1 vccd1 _10226_/C sky130_fd_sc_hd__inv_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06042__B1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10076_ _10076_/A _10001_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__or2b_1
XANTENNA__08334__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10978_ _10978_/CLK _10978_/D vssd1 vssd1 vccd1 vccd1 _10978_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09339__A _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_17_clock_A _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08022__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08810_ _08810_/A _08814_/A _08817_/B vssd1 vssd1 vccd1 vccd1 _08810_/X sky130_fd_sc_hd__or3b_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09790_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__xor2_4
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05953_ _06019_/A _10540_/Q vssd1 vssd1 vccd1 vccd1 _05954_/A sky130_fd_sc_hd__and2_1
X_08741_ _10806_/Q _10805_/Q _10804_/Q _08701_/A _08744_/B vssd1 vssd1 vccd1 vccd1
+ _08741_/X sky130_fd_sc_hd__o41a_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08325__A2 _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05884_ _07988_/A _05883_/X _05878_/B vssd1 vssd1 vccd1 vccd1 _05884_/Y sky130_fd_sc_hd__a21boi_1
X_08672_ _08830_/A vssd1 vssd1 vccd1 vccd1 _08672_/X sky130_fd_sc_hd__buf_2
XFILLER_66_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07623_ _07623_/A _07623_/B vssd1 vssd1 vccd1 vccd1 _07700_/A sky130_fd_sc_hd__xor2_2
XFILLER_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08089__A1 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ _07426_/A _07425_/B _07425_/A vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__o21ba_1
X_07485_ _07485_/A _07485_/B vssd1 vssd1 vccd1 vccd1 _07493_/B sky130_fd_sc_hd__xnor2_2
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06505_ _06521_/A _06517_/C _06503_/Y _06517_/B _06758_/A vssd1 vssd1 vccd1 vccd1
+ _06519_/A sky130_fd_sc_hd__o2111a_1
X_09224_ _09224_/A vssd1 vssd1 vccd1 vccd1 _10852_/D sky130_fd_sc_hd__buf_2
X_06436_ _06436_/A _06456_/A _07682_/B _06460_/B vssd1 vssd1 vccd1 vccd1 _06468_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09155_ _10958_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09155_/Y sky130_fd_sc_hd__nor2_1
X_06367_ _06367_/A _06917_/A vssd1 vssd1 vccd1 vccd1 _06368_/B sky130_fd_sc_hd__nand2_2
X_05318_ _05318_/A _05318_/B vssd1 vssd1 vccd1 vccd1 _05318_/X sky130_fd_sc_hd__and2_1
X_08106_ _08116_/B vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__inv_2
XFILLER_107_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _10491_/A _09085_/X _09086_/S vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__mux2_1
X_06298_ _10920_/Q _10903_/Q vssd1 vssd1 vccd1 vccd1 _06304_/A sky130_fd_sc_hd__nand2_1
X_08037_ _08037_/A vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__buf_2
XFILLER_116_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07992__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09988_ _10065_/C _10065_/B vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08939_ input6/X input5/X _08939_/C input15/X vssd1 vssd1 vccd1 vccd1 _09142_/D sky130_fd_sc_hd__or4b_4
XANTENNA__06401__A _06845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10901_ _10920_/CLK _10901_/D vssd1 vssd1 vccd1 vccd1 _10901_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10832_ _10832_/CLK _10832_/D vssd1 vssd1 vccd1 vccd1 _10832_/Q sky130_fd_sc_hd__dfxtp_2
X_10763_ _10935_/CLK _10763_/D vssd1 vssd1 vccd1 vccd1 _10763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10694_ _10694_/CLK _10694_/D vssd1 vssd1 vccd1 vccd1 _10694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07055__A2 _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08004__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10128_ _10075_/A _10074_/A _10074_/B _10085_/A vssd1 vssd1 vccd1 vccd1 _10146_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08307__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10059_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__nor2_1
XFILLER_48_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09341__B _10909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07270_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07334_/B sky130_fd_sc_hd__or2_1
X_06221_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06221_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06152_ _08166_/A vssd1 vssd1 vccd1 vccd1 _10343_/A sky130_fd_sc_hd__buf_4
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06083_ _05766_/Y _05830_/A _07976_/A _05711_/Y vssd1 vssd1 vccd1 vccd1 _06089_/A
+ sky130_fd_sc_hd__a2bb2o_1
X_09911_ _09911_/A _09911_/B vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__nand2_1
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08701__A _08701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ _09842_/A _09842_/B vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__xnor2_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06221__A _07977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09773_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09773_/X sky130_fd_sc_hd__and2_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _10804_/Q _08701_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08724_/X sky130_fd_sc_hd__o21a_1
XFILLER_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _07007_/A _06997_/C vssd1 vssd1 vccd1 vccd1 _06986_/B sky130_fd_sc_hd__nand2_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05936_ _08277_/B _05858_/Y _05860_/X _05934_/X _05935_/X vssd1 vssd1 vccd1 vccd1
+ _05936_/X sky130_fd_sc_hd__o221a_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05867_ _08233_/A _05866_/X _05863_/X _10699_/Q vssd1 vssd1 vccd1 vccd1 _05867_/X
+ sky130_fd_sc_hd__a22o_1
X_08655_ _08971_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__and2_1
XFILLER_54_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _08586_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _08586_/Y sky130_fd_sc_hd__nor2_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _07606_/A _07606_/B vssd1 vssd1 vccd1 vccd1 _07607_/B sky130_fd_sc_hd__nand2_1
X_05798_ _05798_/A _05798_/B vssd1 vssd1 vccd1 vccd1 _05798_/Y sky130_fd_sc_hd__nor2_1
X_07537_ _07505_/X _07536_/X _07622_/A vssd1 vssd1 vccd1 vccd1 _07606_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07987__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__or2b_1
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _09228_/A _09207_/B vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__and2_1
X_06419_ _06386_/A _06386_/B _06418_/Y vssd1 vssd1 vccd1 vccd1 _06420_/B sky130_fd_sc_hd__o21a_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07399_ _07377_/A _07587_/B _07398_/B _07560_/A vssd1 vssd1 vccd1 vccd1 _07399_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09138_ _07976_/A _09123_/X _09127_/X _09137_/X vssd1 vssd1 vccd1 vccd1 _09138_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09069_ _09639_/B vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08537__A2 _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input12_A io_wbs_m2s_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08058__A _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10815_ _10819_/CLK _10815_/D vssd1 vssd1 vccd1 vccd1 _10815_/Q sky130_fd_sc_hd__dfxtp_1
X_10746_ _10797_/CLK _10746_/D vssd1 vssd1 vccd1 vccd1 _10746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10677_ _10707_/CLK _10677_/D vssd1 vssd1 vccd1 vccd1 _10677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05848__C _05886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08521__A _08935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06976__A _10906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _07682_/A _06842_/A vssd1 vssd1 vccd1 vccd1 _06940_/A sky130_fd_sc_hd__nand2_2
X_05721_ _08082_/C vssd1 vssd1 vccd1 vccd1 _05721_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_82_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10498__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05652_ _05652_/A _05652_/B _05652_/C vssd1 vssd1 vccd1 vccd1 _05652_/X sky130_fd_sc_hd__or3_1
X_08440_ _08440_/A vssd1 vssd1 vccd1 vccd1 _10731_/D sky130_fd_sc_hd__clkbuf_1
X_05583_ _05681_/B _05583_/B vssd1 vssd1 vccd1 vccd1 _05583_/Y sky130_fd_sc_hd__nor2_1
X_08371_ _08547_/A vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__clkbuf_1
X_07322_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07338_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07253_ _07264_/B _07514_/A _07264_/A vssd1 vssd1 vccd1 vccd1 _07254_/B sky130_fd_sc_hd__a21o_1
XFILLER_118_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06204_ _06204_/A _06204_/B vssd1 vssd1 vccd1 vccd1 _06204_/Y sky130_fd_sc_hd__nand2_1
X_07184_ _07184_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07185_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08415__B input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06135_ _09403_/A vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__buf_2
XFILLER_132_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06066_ _08082_/B vssd1 vssd1 vccd1 vccd1 _06066_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09825_ _09814_/B _09825_/B vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__and2b_1
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A io_wbs_m2s_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09756_ _09755_/A _09755_/B _09755_/C vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__a21oi_1
X_06968_ _09381_/A vssd1 vssd1 vccd1 vccd1 _07007_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05919_ _08095_/A _05906_/X _05904_/Y _06037_/A _05918_/X vssd1 vssd1 vccd1 vccd1
+ _05919_/X sky130_fd_sc_hd__a221o_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08707_ _08705_/X _08706_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10803_/D sky130_fd_sc_hd__a21oi_1
XFILLER_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09687_ _09686_/A _09686_/B _09686_/C vssd1 vssd1 vccd1 vccd1 _09755_/B sky130_fd_sc_hd__o21ai_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _10795_/Q _08638_/B _08638_/C vssd1 vssd1 vccd1 vccd1 _08638_/X sky130_fd_sc_hd__and3_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06899_ _06899_/A _06899_/B vssd1 vssd1 vccd1 vccd1 _06928_/A sky130_fd_sc_hd__xnor2_4
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08569_ _08572_/B _08565_/X _08583_/A vssd1 vssd1 vccd1 vccd1 _08569_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ _10811_/CLK _10600_/D vssd1 vssd1 vccd1 vccd1 _10600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10531_ _10531_/A _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10531_/X sky130_fd_sc_hd__or3_1
XANTENNA__10262__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06126__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10462_ _06182_/X _10459_/X _10461_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10957_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10393_ _10389_/X _10717_/Q _10390_/X _10391_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10936_/D sky130_fd_sc_hd__o221a_1
XANTENNA__05965__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10729_ _10935_/CLK _10729_/D vssd1 vssd1 vccd1 vccd1 _10729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08235__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07940_ _08445_/A vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__clkbuf_2
X_07871_ _07871_/A vssd1 vssd1 vccd1 vccd1 _07871_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_95_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06822_ _06823_/A _06823_/B vssd1 vssd1 vccd1 vccd1 _06824_/A sky130_fd_sc_hd__and2_1
X_09610_ _09610_/A _09610_/B _09610_/C _09717_/A vssd1 vssd1 vccd1 vccd1 _09611_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_55_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06753_ _06804_/A _06806_/A vssd1 vssd1 vccd1 vccd1 _06756_/A sky130_fd_sc_hd__nand2_1
X_09541_ _09542_/A _09542_/B _09542_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__a21oi_1
X_05704_ _08188_/A vssd1 vssd1 vccd1 vccd1 _05704_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09472_ _10066_/A _09472_/B vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__nor2_1
X_06684_ _06684_/A _06684_/B vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05635_ _10546_/Q _05635_/B vssd1 vssd1 vccd1 vccd1 _05636_/B sky130_fd_sc_hd__and2_1
X_08423_ _10833_/Q _10832_/Q vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10492__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05566_ _05566_/A _05566_/B vssd1 vssd1 vccd1 vccd1 _05687_/B sky130_fd_sc_hd__and2_1
X_08354_ _08263_/A _08349_/X _08350_/Y _08353_/X _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08354_/X sky130_fd_sc_hd__o32a_1
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07305_ _07305_/A _07305_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__xnor2_1
X_08285_ _08285_/A vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05497_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05497_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_8_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10737_/CLK sky130_fd_sc_hd__clkbuf_16
X_07236_ _07236_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07244_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07167_ _07169_/A _07167_/B vssd1 vssd1 vccd1 vccd1 _07195_/A sky130_fd_sc_hd__nand2_1
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06118_ _07848_/A _06033_/X _06117_/X vssd1 vssd1 vccd1 vccd1 _06119_/B sky130_fd_sc_hd__a21oi_1
XFILLER_133_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_65_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ _07098_/A _07098_/B vssd1 vssd1 vccd1 vccd1 _07219_/B sky130_fd_sc_hd__xnor2_1
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06049_ _10659_/Q vssd1 vssd1 vccd1 vccd1 _07981_/A sky130_fd_sc_hd__buf_2
XFILLER_59_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08373__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _09876_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09809_/B sky130_fd_sc_hd__or2_1
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09739_ _09802_/C vssd1 vssd1 vccd1 vccd1 _09930_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10483__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10514_ _06163_/X _10497_/B _10513_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10977_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _10951_/Q _10431_/X _10444_/X vssd1 vssd1 vccd1 vccd1 _10951_/D sky130_fd_sc_hd__a21o_1
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10376_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07415__A _07415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05420_ _10626_/Q _05378_/Y _05380_/Y _05461_/C _05419_/X vssd1 vssd1 vccd1 vccd1
+ _05420_/X sky130_fd_sc_hd__o221a_1
XFILLER_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05351_ _10634_/Q vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08070_ _08064_/X _08068_/X _08069_/X vssd1 vssd1 vccd1 vccd1 _10681_/D sky130_fd_sc_hd__o21a_1
X_05282_ _10650_/Q vssd1 vssd1 vccd1 vccd1 _06065_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07021_ _07021_/A _07030_/C vssd1 vssd1 vccd1 vccd1 _07421_/A sky130_fd_sc_hd__nand2_2
XFILLER_127_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ _08972_/A vssd1 vssd1 vccd1 vccd1 _08972_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07923_ _10613_/Q _07906_/X _07910_/X _07922_/Y vssd1 vssd1 vccd1 vccd1 _07924_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07854_ hold8/X _07849_/X _07850_/X _07852_/Y _07853_/X vssd1 vssd1 vccd1 vccd1 _07854_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_69_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06805_ _06805_/A _06805_/B vssd1 vssd1 vccd1 vccd1 _06818_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08107__B1 _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07785_ _07785_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _07786_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ _09524_/A _09472_/B vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__or2b_1
X_06736_ _06736_/A vssd1 vssd1 vccd1 vccd1 _07675_/A sky130_fd_sc_hd__buf_2
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06667_ _06667_/A _06671_/A vssd1 vssd1 vccd1 vccd1 _06686_/A sky130_fd_sc_hd__xnor2_1
X_09455_ _09454_/A _09454_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _09456_/C sky130_fd_sc_hd__a21o_1
X_05618_ _10552_/Q _05623_/A _10553_/Q vssd1 vssd1 vccd1 vccd1 _05619_/B sky130_fd_sc_hd__o21ai_1
X_08406_ _08397_/X _10743_/Q _08394_/X hold13/X vssd1 vssd1 vccd1 vccd1 _10725_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09386_ _09449_/A _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__and3_1
X_06598_ _06618_/A _06618_/B vssd1 vssd1 vccd1 vccd1 _06668_/A sky130_fd_sc_hd__xor2_1
X_08337_ input36/X _08248_/X _08088_/X _05574_/X _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08337_/X sky130_fd_sc_hd__o221a_1
X_05549_ _05549_/A _05636_/A vssd1 vssd1 vccd1 vccd1 _05629_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10836__D _10836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08268_ _08268_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08268_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08291__C1 _08258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07219_ _10980_/Q _07219_/B vssd1 vssd1 vccd1 vccd1 _07249_/B sky130_fd_sc_hd__and2_1
X_08199_ _08208_/B _08061_/A _08197_/Y _08198_/Y _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08199_/X sky130_fd_sc_hd__a311o_1
XFILLER_106_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _10246_/B _10228_/A _10291_/S vssd1 vssd1 vccd1 vccd1 _10231_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10161_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__xnor2_1
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10092_ _10155_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__a21oi_1
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05962__B _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08821__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10428_ _06206_/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__a21bo_1
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10359_ _10351_/X _06806_/B _10355_/X _10926_/Q vssd1 vssd1 vccd1 vccd1 _10926_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06060__A1 _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09344__B _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07570_ _07570_/A _09920_/B _07570_/C vssd1 vssd1 vccd1 vccd1 _07571_/B sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_13_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06521_ _06521_/A _06521_/B vssd1 vssd1 vccd1 vccd1 _06522_/C sky130_fd_sc_hd__xor2_1
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ _10820_/Q _09210_/X _09212_/X _09238_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09241_/B sky130_fd_sc_hd__a32o_1
XFILLER_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05323__B1 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06452_ _06626_/A _06568_/B _06451_/C vssd1 vssd1 vccd1 vccd1 _06453_/B sky130_fd_sc_hd__a21oi_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clock _10981_/CLK vssd1 vssd1 vccd1 vccd1 _10976_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05403_ _10649_/Q vssd1 vssd1 vccd1 vccd1 _05405_/A sky130_fd_sc_hd__clkinv_2
X_09171_ _05883_/A _09123_/X _09203_/A _09170_/X vssd1 vssd1 vccd1 vccd1 _09171_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09065__A1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06383_ _06872_/A _06872_/B _06383_/C vssd1 vssd1 vccd1 vccd1 _06874_/A sky130_fd_sc_hd__and3_1
X_08122_ _08114_/X _08130_/B _08116_/Y _08121_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08122_/X sky130_fd_sc_hd__o311a_1
XFILLER_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05334_ _10672_/Q vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08812__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ _09403_/A vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__clkbuf_4
X_07004_ _07211_/A vssd1 vssd1 vccd1 vccd1 _07188_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10836_/CLK sky130_fd_sc_hd__clkbuf_16
X_08955_ _10963_/Q vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08328__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _07906_/A vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08879__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08886_ _08814_/X _08883_/Y _08884_/X _08885_/X vssd1 vssd1 vccd1 vccd1 _10824_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_57_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ _07827_/X _05462_/B _07823_/X _07836_/Y vssd1 vssd1 vccd1 vccd1 _10622_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_26_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10945_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07768_ _07768_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07769_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09270__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10438__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06719_ _06719_/A _06719_/B _06719_/C vssd1 vssd1 vccd1 vccd1 _06720_/B sky130_fd_sc_hd__and3_1
X_09507_ _09507_/A _09676_/C vssd1 vssd1 vccd1 vccd1 _09508_/B sky130_fd_sc_hd__xnor2_4
XFILLER_37_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07699_ _09690_/A _09690_/B _07698_/X vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__o21ai_4
XFILLER_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _09438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09056__A1 _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ _10889_/Q _10905_/Q vssd1 vssd1 vccd1 vccd1 _09369_/X sky130_fd_sc_hd__and2b_1
XFILLER_40_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08031__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10213_ _10950_/Q _10934_/Q vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06042__B2 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05973__A _10432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10144_ _10144_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input42_A io_wbs_m2s_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09531__A2 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10977_ _10978_/CLK _10977_/D vssd1 vssd1 vccd1 vccd1 _10977_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05883__A _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09355__A _10905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07781__A1 _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05952_ _10583_/Q vssd1 vssd1 vccd1 vccd1 _06019_/A sky130_fd_sc_hd__buf_2
X_08740_ _08740_/A _08740_/B _08740_/C vssd1 vssd1 vccd1 vccd1 _08740_/X sky130_fd_sc_hd__and3_1
XANTENNA__07781__B2 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05883_ _05883_/A _10659_/Q _05891_/A vssd1 vssd1 vccd1 vccd1 _05883_/X sky130_fd_sc_hd__or3_1
X_08671_ _08671_/A vssd1 vssd1 vccd1 vccd1 _08830_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07622_ _07622_/A _07622_/B vssd1 vssd1 vccd1 vccd1 _07623_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08089__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07553_ _07430_/A _07430_/B _07429_/A vssd1 vssd1 vccd1 vccd1 _07558_/B sky130_fd_sc_hd__o21a_1
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07484_ _07509_/A _07025_/Y _07483_/X vssd1 vssd1 vccd1 vccd1 _07485_/B sky130_fd_sc_hd__o21a_1
X_06504_ _06517_/A vssd1 vssd1 vccd1 vccd1 _06758_/A sky130_fd_sc_hd__clkbuf_2
X_09223_ _09228_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__and2_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06435_ _06435_/A vssd1 vssd1 vccd1 vccd1 _06486_/A sky130_fd_sc_hd__clkinv_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09154_ _09154_/A vssd1 vssd1 vccd1 vccd1 _09202_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08105_ _08105_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__nor2_1
X_06366_ _10978_/Q _06459_/B vssd1 vssd1 vccd1 vccd1 _06917_/A sky130_fd_sc_hd__nand2_4
XFILLER_135_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05317_ _08352_/A _05827_/A vssd1 vssd1 vccd1 vccd1 _05318_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _10937_/Q _09008_/X _08947_/A _10953_/Q vssd1 vssd1 vccd1 vccd1 _09085_/X
+ sky130_fd_sc_hd__a22o_1
X_06297_ _10921_/Q _09356_/A _06416_/A _06302_/B vssd1 vssd1 vccd1 vccd1 _06730_/A
+ sky130_fd_sc_hd__a31oi_2
X_08036_ _08236_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08074_/A sky130_fd_sc_hd__nor2_2
XFILLER_103_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07772__A1 _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _09921_/B _09922_/B _09377_/X vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__o21ai_1
XFILLER_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08938_ _08938_/A vssd1 vssd1 vccd1 vccd1 _10833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ _08814_/X _08866_/X _08867_/Y _08868_/X vssd1 vssd1 vccd1 vccd1 _10822_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10900_ _10920_/CLK _10900_/D vssd1 vssd1 vccd1 vccd1 _10900_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09204__S _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10831_ _10832_/CLK _10831_/D vssd1 vssd1 vccd1 vccd1 _10831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06129__A _10432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10762_ _10833_/CLK _10762_/D vssd1 vssd1 vccd1 vccd1 _10762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10693_ _10845_/CLK _10693_/D vssd1 vssd1 vccd1 vccd1 _10693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09201__A1 _09112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06799__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10127_ _10087_/A _10087_/B _10090_/A vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__o21a_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10058_ _10487_/A _10123_/B _10057_/C vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06311__B _10909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05829__B2 _08032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06220_ _10602_/Q _06223_/B vssd1 vssd1 vccd1 vccd1 _06220_/X sky130_fd_sc_hd__or2_1
XFILLER_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06151_ _06151_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06151_/Y sky130_fd_sc_hd__nand2_1
X_06082_ _06082_/A _06082_/B _06082_/C _06081_/X vssd1 vssd1 vccd1 vccd1 _06082_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06254__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09910_ _09910_/A _10049_/C vssd1 vssd1 vccd1 vccd1 _09911_/B sky130_fd_sc_hd__nand2_1
XFILLER_113_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10338__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09841_ _09841_/A _09841_/B vssd1 vssd1 vccd1 vccd1 _09842_/B sky130_fd_sc_hd__nor2_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09772_ _09844_/B _09772_/B vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__and2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _07083_/A _07061_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _06997_/C sky130_fd_sc_hd__or3_1
X_05935_ _10702_/Q _05935_/B vssd1 vssd1 vccd1 vccd1 _05935_/X sky130_fd_sc_hd__or2_1
XFILLER_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08723_ _08919_/B vssd1 vssd1 vccd1 vccd1 _08918_/B sky130_fd_sc_hd__buf_2
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05866_ _05350_/B _05854_/B _05865_/Y vssd1 vssd1 vccd1 vccd1 _05866_/X sky130_fd_sc_hd__o21a_1
XFILLER_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08654_ _09016_/A _09126_/A vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__nor2_1
X_05797_ _08160_/A _05694_/Y _05712_/Y _08146_/A _05713_/X vssd1 vssd1 vccd1 vccd1
+ _05798_/B sky130_fd_sc_hd__o221a_1
X_08585_ _10781_/Q _10780_/Q _08585_/C vssd1 vssd1 vccd1 vccd1 _08586_/B sky130_fd_sc_hd__and3_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07605_ _07708_/A _07605_/B vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__xor2_2
XFILLER_26_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07536_ _07617_/B _07618_/B vssd1 vssd1 vccd1 vccd1 _07536_/X sky130_fd_sc_hd__or2_1
XFILLER_22_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09206_ _08815_/A _09168_/X _09203_/X _09205_/X vssd1 vssd1 vccd1 vccd1 _09207_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07467_ _07746_/A _07469_/B _07466_/Y vssd1 vssd1 vccd1 vccd1 _07499_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08164__A _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08219__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06418_ _10921_/Q _07061_/A vssd1 vssd1 vccd1 vccd1 _06418_/Y sky130_fd_sc_hd__nand2_1
X_07398_ _07728_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07753_/A sky130_fd_sc_hd__nand2_2
X_09137_ _05461_/C _09136_/X _06212_/B _08150_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09137_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10844__D _10844_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06349_ _06436_/A _06568_/B vssd1 vssd1 vccd1 vccd1 _06457_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06245__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ _10968_/Q vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08019_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08019_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10814_ _10814_/CLK _10814_/D vssd1 vssd1 vccd1 vccd1 _10814_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10745_ _10855_/CLK _10745_/D vssd1 vssd1 vccd1 vccd1 _10745_/Q sky130_fd_sc_hd__dfxtp_1
X_10676_ _10676_/CLK _10676_/D vssd1 vssd1 vccd1 vccd1 _10676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10109__A _10109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08521__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07418__A _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07736__A1 _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05720_ _08082_/A _05536_/B _05737_/B _08082_/B vssd1 vssd1 vccd1 vccd1 _05794_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08161__A1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05651_ _05652_/A _05652_/B _05652_/C vssd1 vssd1 vccd1 vccd1 _05651_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_63_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08370_ _10251_/S vssd1 vssd1 vccd1 vccd1 _08547_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05582_ _05769_/A _05582_/B vssd1 vssd1 vccd1 vccd1 _05583_/B sky130_fd_sc_hd__and2_1
X_07321_ _07560_/A _07394_/A _07151_/C vssd1 vssd1 vccd1 vccd1 _07322_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07252_ _07513_/A _07516_/A vssd1 vssd1 vccd1 vccd1 _07514_/A sky130_fd_sc_hd__or2_1
XFILLER_117_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06203_ _10598_/Q vssd1 vssd1 vccd1 vccd1 _06204_/A sky130_fd_sc_hd__inv_2
X_07183_ _07183_/A _07183_/B vssd1 vssd1 vccd1 vccd1 _07208_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06134_ _06134_/A _06145_/B vssd1 vssd1 vccd1 vccd1 _06134_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07975__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06065_ _06065_/A vssd1 vssd1 vccd1 vccd1 _06065_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_99_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__xnor2_2
XFILLER_86_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09755_/A _09755_/B _09755_/C vssd1 vssd1 vccd1 vccd1 _09755_/X sky130_fd_sc_hd__and3_1
X_06967_ _07112_/A vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__clkbuf_4
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05918_ _08095_/A _05906_/X _05909_/Y _05718_/A _05917_/X vssd1 vssd1 vccd1 vccd1
+ _05918_/X sky130_fd_sc_hd__o221a_1
X_08706_ _10531_/A _08672_/X _08674_/X _08701_/A vssd1 vssd1 vccd1 vccd1 _08706_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_73_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09686_ _09686_/A _09686_/B _09686_/C vssd1 vssd1 vccd1 vccd1 _09686_/X sky130_fd_sc_hd__or3_1
X_06898_ _06930_/A _06930_/B vssd1 vssd1 vccd1 vccd1 _06936_/A sky130_fd_sc_hd__xor2_4
XANTENNA__10839__D _10839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05849_ _10667_/Q _10666_/Q _10665_/Q _05872_/A vssd1 vssd1 vccd1 vccd1 _05863_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08637_ _08638_/B _08638_/C _08636_/Y vssd1 vssd1 vccd1 vccd1 _10794_/D sky130_fd_sc_hd__o21a_1
XANTENNA__07998__A _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08568_ _08568_/A vssd1 vssd1 vccd1 vccd1 _10775_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_clock_A _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08499_ _08498_/X _08496_/X _08494_/X _10748_/Q vssd1 vssd1 vccd1 vccd1 _10748_/D
+ sky130_fd_sc_hd__a22o_1
X_07519_ _09303_/B _07519_/B vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__or2_1
X_10530_ _07732_/A _10522_/X _10528_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10982_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10262__A2 _10115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10461_ _10957_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or2_1
XFILLER_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06126__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09718__A _09930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06142__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05981__A _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08143__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08143__B2 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10728_ _10839_/CLK _10728_/D vssd1 vssd1 vccd1 vccd1 _10728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10659_ _10694_/CLK _10659_/D vssd1 vssd1 vccd1 vccd1 _10659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07870_ _07906_/A vssd1 vssd1 vccd1 vccd1 _07870_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_95_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06821_ _06821_/A _06821_/B vssd1 vssd1 vccd1 vccd1 _06823_/B sky130_fd_sc_hd__xor2_1
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06752_ _06752_/A _06752_/B _06752_/C _06746_/A vssd1 vssd1 vccd1 vccd1 _06806_/A
+ sky130_fd_sc_hd__or4b_1
X_09540_ _09458_/A _09599_/A _09696_/A vssd1 vssd1 vccd1 vccd1 _09542_/C sky130_fd_sc_hd__nand3b_1
XFILLER_37_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08134__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05703_ _10693_/Q vssd1 vssd1 vccd1 vccd1 _08188_/A sky130_fd_sc_hd__clkbuf_2
X_09471_ _09471_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09472_/B sky130_fd_sc_hd__and2_1
XFILLER_36_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08422_ _10763_/Q _10764_/Q _08421_/Y vssd1 vssd1 vccd1 vccd1 _08424_/A sky130_fd_sc_hd__o21ai_2
XFILLER_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06683_ _06945_/A _06945_/B _06948_/A vssd1 vssd1 vccd1 vccd1 _06943_/C sky130_fd_sc_hd__or3_1
XFILLER_36_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05634_ _10685_/Q vssd1 vssd1 vccd1 vccd1 _06037_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05565_ _10570_/Q _05576_/A _10571_/Q vssd1 vssd1 vccd1 vccd1 _05566_/B sky130_fd_sc_hd__o21ai_1
X_08353_ _08037_/A _06115_/B _08351_/Y _08352_/Y vssd1 vssd1 vccd1 vccd1 _08353_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08284_ _08284_/A _08284_/B vssd1 vssd1 vccd1 vccd1 _10702_/D sky130_fd_sc_hd__nor2_1
X_07304_ _07289_/A _07304_/B vssd1 vssd1 vccd1 vccd1 _07305_/A sky130_fd_sc_hd__and2b_1
X_05496_ _05380_/Y _05489_/X _05495_/X _05461_/C vssd1 vssd1 vccd1 vccd1 _10550_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07235_ _07515_/A _07235_/B _07235_/C vssd1 vssd1 vccd1 vccd1 _07237_/B sky130_fd_sc_hd__and3b_1
X_07166_ _07166_/A _07166_/B vssd1 vssd1 vccd1 vccd1 _07334_/A sky130_fd_sc_hd__nand2_1
X_06117_ _08065_/B _08258_/A _06117_/C _06117_/D vssd1 vssd1 vccd1 vccd1 _06117_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_106_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07097_ _10913_/Q _07102_/A vssd1 vssd1 vccd1 vccd1 _07098_/B sky130_fd_sc_hd__nand2_1
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06048_ _10710_/Q _08032_/A _06045_/X _06047_/X vssd1 vssd1 vccd1 vccd1 _06071_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09273__A _09273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ input23/X _07987_/X _07998_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10664_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09807_ _09807_/A _09856_/C vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10180__A1 _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09738_ _09919_/B vssd1 vssd1 vccd1 vccd1 _10129_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10212__A _10934_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09669_ _09731_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09671_/B sky130_fd_sc_hd__or2_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06137__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10513_ _10513_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10513_/X sky130_fd_sc_hd__or2_1
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08352__A _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05976__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _05958_/X _10440_/B _05977_/X vssd1 vssd1 vccd1 vccd1 _10444_/X sky130_fd_sc_hd__a21o_1
XFILLER_40_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10375_ _10932_/Q _10379_/B vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__and2_1
XFILLER_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10171__A1 _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10122__A _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07431__A _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05350_ _10667_/Q _05350_/B vssd1 vssd1 vccd1 vccd1 _05350_/X sky130_fd_sc_hd__xor2_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05281_ _10575_/Q vssd1 vssd1 vccd1 vccd1 _05454_/A sky130_fd_sc_hd__inv_2
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07020_ _07021_/A _07020_/B vssd1 vssd1 vccd1 vccd1 _07509_/A sky130_fd_sc_hd__nand2_2
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08971_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _08972_/A sky130_fd_sc_hd__nand2_1
X_07922_ _07922_/A vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__clkinv_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07853_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07853_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09093__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06804_ _06804_/A vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__buf_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07784_ _10510_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07785_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06118__B1 _06117_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09523_ _10131_/A vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__clkbuf_2
X_06735_ _06735_/A _06735_/B vssd1 vssd1 vccd1 vccd1 _06746_/A sky130_fd_sc_hd__xor2_4
XFILLER_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06666_ _06666_/A _06666_/B vssd1 vssd1 vccd1 vccd1 _06667_/A sky130_fd_sc_hd__nand2_1
X_09454_ _09454_/A _09454_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__nand3_1
X_05617_ _10552_/Q _05623_/A vssd1 vssd1 vccd1 vccd1 _05617_/X sky130_fd_sc_hd__xor2_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08405_ _08408_/A _10759_/Q vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__or2_1
X_09385_ _09810_/A _09383_/A _09417_/A vssd1 vssd1 vccd1 vccd1 _09533_/C sky130_fd_sc_hd__a21o_1
XFILLER_24_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08336_ _05574_/X _08339_/C _08335_/Y vssd1 vssd1 vccd1 vccd1 _08336_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06597_ _06549_/A _06597_/B _06597_/C vssd1 vssd1 vccd1 vccd1 _06618_/B sky130_fd_sc_hd__nand3b_1
XFILLER_138_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05548_ _10546_/Q _05635_/B vssd1 vssd1 vccd1 vccd1 _05636_/A sky130_fd_sc_hd__nor2_1
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08267_ _08267_/A _08267_/B vssd1 vssd1 vccd1 vccd1 _08267_/Y sky130_fd_sc_hd__nand2_1
X_05479_ _05479_/A vssd1 vssd1 vccd1 vccd1 _05489_/A sky130_fd_sc_hd__clkbuf_2
X_08198_ _08198_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08198_/Y sky130_fd_sc_hd__nor2_1
X_07218_ _07222_/A _07215_/B _07216_/B _10979_/Q vssd1 vssd1 vccd1 vccd1 _07218_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10852__D _10852_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _07511_/A _07327_/A _07149_/C vssd1 vssd1 vccd1 vccd1 _07150_/B sky130_fd_sc_hd__and3b_1
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10207__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10091_ _10155_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10121_/S sky130_fd_sc_hd__and3_1
XFILLER_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10427_ _10946_/Q _10427_/B vssd1 vssd1 vccd1 vccd1 _10427_/X sky130_fd_sc_hd__and2_1
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10117__A _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _10351_/X _06752_/A _10355_/X _10925_/Q vssd1 vssd1 vccd1 vccd1 _10925_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10289_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10289_/X sky130_fd_sc_hd__or2_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_7_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06520_ _06532_/A _06523_/B _06523_/C vssd1 vssd1 vccd1 vccd1 _06520_/X sky130_fd_sc_hd__a21o_1
X_06451_ _06456_/A _06568_/B _06451_/C vssd1 vssd1 vccd1 vccd1 _06453_/A sky130_fd_sc_hd__and3_1
XFILLER_22_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05323__A1 _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05402_ _10618_/Q _05483_/A vssd1 vssd1 vccd1 vccd1 _05402_/X sky130_fd_sc_hd__or2_1
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09170_ _05460_/D _09136_/X _09148_/X _08180_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09170_/X sky130_fd_sc_hd__a221o_1
X_06382_ _06394_/A _06382_/B vssd1 vssd1 vccd1 vccd1 _06383_/C sky130_fd_sc_hd__or2_1
X_08121_ _08132_/B _08061_/A _08117_/Y _08119_/Y _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08121_/X sky130_fd_sc_hd__a311o_1
X_05333_ _10640_/Q vssd1 vssd1 vccd1 vccd1 _07903_/A sky130_fd_sc_hd__clkbuf_2
X_08052_ _08052_/A vssd1 vssd1 vccd1 vccd1 _08052_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08812__A2 _08672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07003_ _10981_/Q vssd1 vssd1 vccd1 vccd1 _07211_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08954_ _09098_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _10474_/B sky130_fd_sc_hd__nor2_2
XANTENNA__08328__A1 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _07916_/A _07905_/B vssd1 vssd1 vccd1 vccd1 _10640_/D sky130_fd_sc_hd__nor2_1
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08885_ input33/X _08819_/X _08820_/X _10824_/Q _10412_/A vssd1 vssd1 vccd1 vccd1
+ _08885_/X sky130_fd_sc_hd__o221a_1
XFILLER_84_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10135__B2 _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07836_ _06165_/A _07828_/X _07829_/X _07835_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07836_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07767_ _10506_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _07768_/B sky130_fd_sc_hd__nand2_1
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09506_ _09506_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09676_/C sky130_fd_sc_hd__nor2_2
X_06718_ _06718_/A _06718_/B vssd1 vssd1 vccd1 vccd1 _06720_/A sky130_fd_sc_hd__nand2_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07698_ _07698_/A _07698_/B vssd1 vssd1 vccd1 vccd1 _07698_/X sky130_fd_sc_hd__or2_1
XFILLER_80_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10847__D _10847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09437_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__or2_1
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06649_ _06663_/A _06692_/A _06692_/B _06622_/B vssd1 vssd1 vccd1 vccd1 _06650_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09676_/A _09546_/A _09546_/B _09367_/Y _09356_/A vssd1 vssd1 vccd1 vccd1
+ _09607_/A sky130_fd_sc_hd__a32o_1
XFILLER_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08319_ _08324_/B _08253_/X _08317_/Y _08318_/Y vssd1 vssd1 vccd1 vccd1 _08319_/X
+ sky130_fd_sc_hd__a31o_1
X_09299_ _10343_/A _09299_/B vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__and2_1
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06134__B _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10212_ _10934_/Q _10950_/Q vssd1 vssd1 vccd1 vccd1 _10226_/B sky130_fd_sc_hd__or2b_1
XANTENNA__06042__A2 _08021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10143_ _10143_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10144_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input35_A io_wbs_m2s_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06150__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__nor2_1
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10429__A2 _10727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10976_/CLK _10976_/D vssd1 vssd1 vccd1 vccd1 _10976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05951_ _05717_/X _05788_/X _05809_/X _05950_/Y vssd1 vssd1 vccd1 vccd1 _10540_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05882_ _10658_/Q _05895_/A vssd1 vssd1 vccd1 vccd1 _05891_/A sky130_fd_sc_hd__or2_1
XFILLER_94_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08670_ _08670_/A _08670_/B _08670_/C vssd1 vssd1 vccd1 vccd1 _08670_/X sky130_fd_sc_hd__and3_1
XANTENNA__06995__A _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08730__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07621_ _07621_/A _07702_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__xnor2_2
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07552_ _07448_/A _07448_/B _07447_/A vssd1 vssd1 vccd1 vccd1 _07583_/B sky130_fd_sc_hd__o21ba_1
X_06503_ _06503_/A _06503_/B vssd1 vssd1 vccd1 vccd1 _06503_/Y sky130_fd_sc_hd__nor2_1
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07483_ _07442_/X _07728_/B _07729_/B _07715_/C vssd1 vssd1 vccd1 vccd1 _07483_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09222_ _10817_/Q _09210_/X _09212_/X _09221_/X _09203_/X vssd1 vssd1 vccd1 vccd1
+ _09223_/B sky130_fd_sc_hd__a32o_1
X_06434_ _06434_/A _06434_/B vssd1 vssd1 vccd1 vccd1 _06435_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08246__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09153_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _10844_/D sky130_fd_sc_hd__nor2_4
X_06365_ _07682_/B _06365_/B _06451_/C _06367_/A vssd1 vssd1 vccd1 vccd1 _06872_/B
+ sky130_fd_sc_hd__or4b_1
X_05316_ _08034_/A _05318_/A vssd1 vssd1 vccd1 vccd1 _05525_/B sky130_fd_sc_hd__xnor2_4
X_08104_ _08105_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _08104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09084_ _09908_/A vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__clkbuf_4
X_06296_ _10922_/Q _10905_/Q vssd1 vssd1 vccd1 vccd1 _06302_/B sky130_fd_sc_hd__and2_1
X_08035_ input40/X _07985_/B _08034_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10679_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09986_ _09925_/A _09924_/B _10131_/A vssd1 vssd1 vccd1 vccd1 _09990_/A sky130_fd_sc_hd__o21ai_1
XFILLER_103_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08937_ _10832_/Q _10529_/A vssd1 vssd1 vccd1 vccd1 _08938_/A sky130_fd_sc_hd__and2_1
X_08868_ input31/X _08819_/X _08820_/X _10822_/Q _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08868_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07819_ _06255_/X _09020_/A _06257_/X hold20/X vssd1 vssd1 vccd1 vccd1 _10618_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08799_ _06206_/X _08785_/X _08786_/X _10814_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08799_/X sky130_fd_sc_hd__o221a_1
X_10830_ _10830_/CLK _10830_/D vssd1 vssd1 vccd1 vccd1 _10830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05314__A _10677_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ _10955_/CLK _10761_/D vssd1 vssd1 vccd1 vccd1 _10761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10692_ _10845_/CLK _10692_/D vssd1 vssd1 vccd1 vccd1 _10692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06248__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05968__B input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_56_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10347__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10126_ _10126_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10057_ _10057_/A _10123_/B _10057_/C vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__and3_1
XFILLER_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ _10960_/CLK _10959_/D vssd1 vssd1 vccd1 vccd1 _10959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_10_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10791_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08535__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08779__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06150_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06170_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09440__A2 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06081_ _08282_/A _05851_/A _08198_/A _08196_/A _06080_/X vssd1 vssd1 vccd1 vccd1
+ _06081_/X sky130_fd_sc_hd__o221a_1
XANTENNA__06254__A2 _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10803_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09840_ _09974_/A _09839_/B _09839_/C vssd1 vssd1 vccd1 vccd1 _09841_/B sky130_fd_sc_hd__a21oi_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09771_ _09771_/A _09771_/B _09771_/C vssd1 vssd1 vccd1 vccd1 _09772_/B sky130_fd_sc_hd__or3_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _07066_/A _07056_/A _10901_/Q _07475_/B vssd1 vssd1 vccd1 vccd1 _07060_/B
+ sky130_fd_sc_hd__or4_1
X_05934_ _08251_/B _05863_/X _05867_/X _05932_/X _05933_/X vssd1 vssd1 vccd1 vccd1
+ _05934_/X sky130_fd_sc_hd__o221a_1
X_08722_ _08902_/B vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05865_ _05358_/A _05823_/A _10666_/Q vssd1 vssd1 vccd1 vccd1 _05865_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08653_ _08651_/Y _08649_/C _08652_/X vssd1 vssd1 vccd1 vccd1 _10798_/D sky130_fd_sc_hd__a21oi_1
XFILLER_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05796_ _05788_/B _05794_/Y _05795_/Y vssd1 vssd1 vccd1 vccd1 _05796_/X sky130_fd_sc_hd__o21a_1
X_08584_ _10780_/Q _08585_/C _08583_/Y vssd1 vssd1 vccd1 vccd1 _10780_/D sky130_fd_sc_hd__o21a_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06190__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07604_ _07604_/A _07604_/B vssd1 vssd1 vccd1 vccd1 _07605_/B sky130_fd_sc_hd__xor2_4
X_07535_ _07535_/A _07535_/B vssd1 vssd1 vccd1 vccd1 _07618_/B sky130_fd_sc_hd__nor2_1
X_07466_ _07466_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07466_/Y sky130_fd_sc_hd__nand2_1
X_09205_ _07998_/A _09204_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__mux2_1
X_06417_ _09356_/A vssd1 vssd1 vccd1 vccd1 _07061_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07397_ _07397_/A _07397_/B vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__xnor2_2
XFILLER_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09136_ _09136_/A vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06348_ _06547_/C vssd1 vssd1 vccd1 vccd1 _06568_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09067_ _07727_/A _08965_/Y _09036_/X _09063_/X _09066_/X vssd1 vssd1 vccd1 vccd1
+ _09067_/X sky130_fd_sc_hd__a221o_1
X_06279_ _06558_/B _06558_/C vssd1 vssd1 vccd1 vccd1 _06338_/A sky130_fd_sc_hd__and2_1
X_08018_ _08018_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08018_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08180__A _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _09969_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__xnor2_2
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09215__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06181__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10813_ _10813_/CLK _10813_/D vssd1 vssd1 vccd1 vccd1 _10813_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10744_ _10781_/CLK _10744_/D vssd1 vssd1 vccd1 vccd1 _10744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10675_ _10676_/CLK _10675_/D vssd1 vssd1 vccd1 vccd1 _10675_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10109_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10162_/B sky130_fd_sc_hd__xor2_1
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08161__A2 _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05650_ _10683_/Q vssd1 vssd1 vccd1 vccd1 _05718_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05581_ _10567_/Q _05582_/B vssd1 vssd1 vccd1 vccd1 _05681_/B sky130_fd_sc_hd__nor2_1
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07320_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07488_/B sky130_fd_sc_hd__nor2_1
X_07251_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06202_ input21/X vssd1 vssd1 vccd1 vccd1 _06202_/X sky130_fd_sc_hd__clkbuf_4
X_07182_ _07183_/A _07183_/B vssd1 vssd1 vccd1 vccd1 _07280_/B sky130_fd_sc_hd__and2_1
X_06133_ _06149_/A vssd1 vssd1 vccd1 vccd1 _06145_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_132_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06064_ _05767_/Y _10675_/Q _06050_/X _09104_/A vssd1 vssd1 vccd1 vccd1 _06069_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08924__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09823_ _10876_/Q _09572_/X _09822_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10876_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _09754_/A _09754_/B vssd1 vssd1 vccd1 vccd1 _09755_/C sky130_fd_sc_hd__xnor2_1
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06966_ _06966_/A _06966_/B vssd1 vssd1 vccd1 vccd1 _07708_/A sky130_fd_sc_hd__xnor2_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05917_ _05718_/A _05909_/Y _05911_/Y _05719_/A _05916_/X vssd1 vssd1 vccd1 vccd1
+ _05917_/X sky130_fd_sc_hd__a221o_1
X_08705_ _08808_/A _08705_/B _08725_/A vssd1 vssd1 vccd1 vccd1 _08705_/X sky130_fd_sc_hd__or3_1
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09685_ _09689_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09686_/C sky130_fd_sc_hd__xnor2_1
XFILLER_27_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06897_ _06894_/A _06894_/B _06899_/A _06899_/B vssd1 vssd1 vccd1 vccd1 _06930_/B
+ sky130_fd_sc_hd__a22oi_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05848_ _06052_/A _05848_/B _05886_/B vssd1 vssd1 vccd1 vccd1 _05872_/A sky130_fd_sc_hd__or3_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _08638_/B _08638_/C _08592_/A vssd1 vssd1 vccd1 vccd1 _08636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05779_ _08355_/A _10571_/Q _10572_/Q _05778_/Y vssd1 vssd1 vccd1 vccd1 _05785_/B
+ sky130_fd_sc_hd__o22a_1
X_08567_ _08432_/Y _08565_/X _08567_/C _08567_/D vssd1 vssd1 vccd1 vccd1 _08568_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08175__A _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08498_ _10785_/Q vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07518_ _07573_/A _07394_/X _07327_/X _07021_/A vssd1 vssd1 vccd1 vccd1 _07519_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07449_ _07562_/C _07573_/C _07373_/A vssd1 vssd1 vccd1 vccd1 _07551_/B sky130_fd_sc_hd__o21ai_1
XFILLER_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ _10472_/B vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09119_ _10500_/B vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10391_ _10533_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10391_/X sky130_fd_sc_hd__a21bo_1
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08143__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06154__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08300__C1 _08258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10727_ _10737_/CLK _10727_/D vssd1 vssd1 vccd1 vccd1 _10727_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10658_ _10694_/CLK _10658_/D vssd1 vssd1 vccd1 vccd1 _10658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10589_ _10813_/CLK _10589_/D vssd1 vssd1 vccd1 vccd1 _10589_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06090__B1 _10579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06820_ _07779_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _06821_/B sky130_fd_sc_hd__xor2_2
XFILLER_95_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ _06748_/X _06772_/A _06771_/B vssd1 vssd1 vccd1 vccd1 _06779_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05702_ _05702_/A _10556_/Q vssd1 vssd1 vccd1 vccd1 _05702_/X sky130_fd_sc_hd__and2_1
X_09470_ _09520_/A _09470_/B vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__and2_1
X_06682_ _06947_/A _06947_/B vssd1 vssd1 vccd1 vccd1 _06948_/A sky130_fd_sc_hd__or2_1
X_08421_ _10763_/Q _10764_/Q _10765_/Q vssd1 vssd1 vccd1 vccd1 _08421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05633_ _10686_/Q vssd1 vssd1 vccd1 vccd1 _05726_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05564_ _05564_/A _05566_/A vssd1 vssd1 vccd1 vccd1 _05564_/Y sky130_fd_sc_hd__xnor2_2
X_08352_ _08352_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08352_/Y sky130_fd_sc_hd__nor2_1
X_08283_ _08274_/Y _08248_/X _08157_/A _08281_/X _08282_/X vssd1 vssd1 vccd1 vccd1
+ _08284_/B sky130_fd_sc_hd__o221a_1
X_05495_ _05495_/A vssd1 vssd1 vccd1 vccd1 _05495_/X sky130_fd_sc_hd__clkbuf_2
X_07303_ _07307_/A _07307_/B vssd1 vssd1 vccd1 vccd1 _07349_/C sky130_fd_sc_hd__nor2_1
X_07234_ _10981_/Q _07382_/A vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__and2_1
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07165_ _07196_/A vssd1 vssd1 vccd1 vccd1 _07184_/A sky130_fd_sc_hd__inv_2
X_06116_ _08062_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _06117_/D sky130_fd_sc_hd__or2_2
X_07096_ _07363_/C _07096_/B vssd1 vssd1 vccd1 vccd1 _07355_/A sky130_fd_sc_hd__and2_1
X_06047_ _08209_/A _05702_/A _10704_/Q _08018_/A vssd1 vssd1 vccd1 vccd1 _06047_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_120_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07998_ _07998_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _07998_/X sky130_fd_sc_hd__or2_1
XFILLER_87_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09806_ _09807_/A _09856_/C vssd1 vssd1 vccd1 vccd1 _09876_/A sky130_fd_sc_hd__and2_1
XFILLER_47_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09737_ _09737_/A vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__clkbuf_2
X_06949_ _06591_/Y _06949_/B vssd1 vssd1 vccd1 vccd1 _06950_/A sky130_fd_sc_hd__and2b_1
XFILLER_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__and2_1
XFILLER_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08619_ _08617_/X _08649_/A _08619_/C vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__and3b_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09599_ _09599_/A _09599_/B vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09086__A0 _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05322__A _10677_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08833__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ _05982_/A _10497_/B _10510_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10976_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10443_ _06147_/X _10431_/X _10440_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10950_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10374_ _10365_/X _10712_/Q _10368_/X _10372_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10931_/D sky130_fd_sc_hd__o221a_1
XANTENNA__06153__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05992__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 _10857_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05280_ _10575_/Q vssd1 vssd1 vccd1 vccd1 _05910_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__05886__B _05886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08970_ _07715_/C _08943_/X _08967_/Y _08969_/Y vssd1 vssd1 vccd1 vccd1 _08970_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07921_ _08284_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _10644_/D sky130_fd_sc_hd__nor2_1
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07852_ _10876_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06803_ _07682_/A vssd1 vssd1 vccd1 vccd1 _07780_/C sky130_fd_sc_hd__buf_2
Xinput1 io_ba_match vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07783_ _10513_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07785_/A sky130_fd_sc_hd__nand2_1
X_09522_ _09563_/B _09522_/B vssd1 vssd1 vccd1 vccd1 _09625_/A sky130_fd_sc_hd__and2_2
X_06734_ _06734_/A _06734_/B vssd1 vssd1 vccd1 vccd1 _06735_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ _09390_/A _09488_/A _10964_/Q vssd1 vssd1 vccd1 vccd1 _09454_/C sky130_fd_sc_hd__and3b_1
X_06665_ _06700_/B _06665_/B vssd1 vssd1 vccd1 vccd1 _06903_/A sky130_fd_sc_hd__xnor2_2
XFILLER_24_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05616_ _10691_/Q vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__clkbuf_2
X_08404_ _08397_/X hold6/X _08394_/X _08403_/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__o211a_1
X_09384_ _09417_/A _09810_/A _09424_/A vssd1 vssd1 vccd1 vccd1 _09533_/B sky130_fd_sc_hd__nand3_2
X_08335_ _05574_/X _08339_/C _08092_/A vssd1 vssd1 vccd1 vccd1 _08335_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06238__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06596_ _06599_/A _06599_/B vssd1 vssd1 vccd1 vccd1 _06597_/C sky130_fd_sc_hd__or2_1
X_05547_ _05547_/A _05637_/B vssd1 vssd1 vccd1 vccd1 _05635_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08266_ _08267_/A _08277_/C vssd1 vssd1 vccd1 vccd1 _08266_/Y sky130_fd_sc_hd__nor2_1
X_05478_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05495_/A sky130_fd_sc_hd__clkbuf_2
X_08197_ _08191_/A _08191_/B _05877_/X vssd1 vssd1 vccd1 vccd1 _08197_/Y sky130_fd_sc_hd__o21ai_1
X_07217_ _07250_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _07217_/Y sky130_fd_sc_hd__nor2_1
X_07148_ _07148_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07152_/B sky130_fd_sc_hd__or2_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06054__B1 _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07079_ _07163_/B _07312_/A _07149_/C vssd1 vssd1 vccd1 vccd1 _07298_/A sky130_fd_sc_hd__or3b_1
XFILLER_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10090_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10091_/C sky130_fd_sc_hd__and2_1
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05317__A _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10426_ _10408_/X _10726_/Q _10424_/X _10425_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10945_/D sky130_fd_sc_hd__o221a_1
XANTENNA__10117__B _10117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10357_ _09634_/A _06746_/A _08494_/X _10924_/Q vssd1 vssd1 vccd1 vccd1 _10924_/D
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10265_/A _10287_/C _10287_/D vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__a21bo_1
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06450_ _06468_/A _06450_/B vssd1 vssd1 vccd1 vccd1 _06477_/A sky130_fd_sc_hd__xnor2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05401_ _05401_/A _05406_/A vssd1 vssd1 vccd1 vccd1 _05483_/A sky130_fd_sc_hd__xnor2_1
XFILLER_92_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06381_ _06895_/A _06895_/B _06381_/C vssd1 vssd1 vccd1 vccd1 _06382_/B sky130_fd_sc_hd__and3_1
X_08120_ _08236_/A vssd1 vssd1 vccd1 vccd1 _08120_/X sky130_fd_sc_hd__buf_2
X_05332_ _08021_/A _05844_/B vssd1 vssd1 vccd1 vccd1 _05332_/Y sky130_fd_sc_hd__xnor2_1
X_08051_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08052_/A sky130_fd_sc_hd__buf_2
XFILLER_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07002_ _07562_/C _07573_/C vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__xor2_1
XANTENNA__06036__B1 _05405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08953_ _10914_/Q _10931_/Q _09008_/A vssd1 vssd1 vccd1 vccd1 _08953_/X sky130_fd_sc_hd__mux2_1
X_07904_ _10608_/Q _07888_/X _07892_/X _07903_/Y vssd1 vssd1 vccd1 vccd1 _07905_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08884_ _08883_/A _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08884_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__10043__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07835_ hold12/X _07845_/B vssd1 vssd1 vccd1 vccd1 _07835_/Y sky130_fd_sc_hd__nand2_1
X_07766_ _10504_/A _07766_/B vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09505_ _07066_/A _10887_/Q vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__and2b_1
XFILLER_25_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06717_ _06717_/A _06717_/B vssd1 vssd1 vccd1 vccd1 _06718_/A sky130_fd_sc_hd__nand2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09477_/B vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07697_ _07637_/A _07637_/B _07696_/X vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__o21a_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06648_ _06648_/A _06648_/B vssd1 vssd1 vccd1 vccd1 _06650_/B sky130_fd_sc_hd__xor2_1
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09367_ _10888_/Q vssd1 vssd1 vccd1 vccd1 _09367_/Y sky130_fd_sc_hd__inv_2
X_06579_ _06581_/A _06581_/C _06581_/B vssd1 vssd1 vccd1 vccd1 _06579_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ _08318_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08318_/Y sky130_fd_sc_hd__nor2_1
X_09298_ _10830_/Q _09274_/X _09275_/X _09297_/X _09127_/X vssd1 vssd1 vccd1 vccd1
+ _09299_/B sky130_fd_sc_hd__a32o_1
X_08249_ input26/X _08248_/X _08088_/X _08243_/A _08394_/A vssd1 vssd1 vccd1 vccd1
+ _08249_/X sky130_fd_sc_hd__o221a_1
XFILLER_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10218__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10211_ _10209_/Y _10210_/X _07747_/A _09406_/X vssd1 vssd1 vccd1 vccd1 _10900_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10142_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_121_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10073_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10074_/B sky130_fd_sc_hd__nor2_1
XFILLER_121_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07961__S _07983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input28_A io_wbs_m2s_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10975_ _10976_/CLK _10975_/D vssd1 vssd1 vccd1 vccd1 _10975_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_52_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05510__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08007__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10409_ _10427_/B vssd1 vssd1 vccd1 vccd1 _10424_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05950_ _05528_/X _05826_/X _05949_/X vssd1 vssd1 vccd1 vccd1 _05950_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_66_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05881_ _06039_/A _10656_/Q _05900_/A vssd1 vssd1 vccd1 vccd1 _05895_/A sky130_fd_sc_hd__or3_1
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_66_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07620_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07702_/B sky130_fd_sc_hd__xnor2_4
XFILLER_53_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07551_ _07450_/A _07551_/B vssd1 vssd1 vccd1 vccd1 _07585_/A sky130_fd_sc_hd__and2b_2
X_06502_ _06561_/B _06502_/B _06502_/C _06506_/B vssd1 vssd1 vccd1 vccd1 _06503_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07482_ _07482_/A _07482_/B vssd1 vssd1 vccd1 vccd1 _07485_/A sky130_fd_sc_hd__nor2_2
X_09221_ _08235_/A _09220_/X _09226_/S vssd1 vssd1 vccd1 vccd1 _09221_/X sky130_fd_sc_hd__mux2_1
X_06433_ _06645_/A _06433_/B vssd1 vssd1 vccd1 vccd1 _06434_/B sky130_fd_sc_hd__or2_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09152_ _09112_/X _09147_/Y _09151_/X vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09099__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06364_ _06719_/A _06460_/B vssd1 vssd1 vccd1 vccd1 _06367_/A sky130_fd_sc_hd__nand2_1
X_08103_ _08117_/B _08102_/Y _06117_/D vssd1 vssd1 vccd1 vccd1 _08103_/Y sky130_fd_sc_hd__a21oi_1
X_05315_ _08352_/A _05827_/A vssd1 vssd1 vccd1 vccd1 _05318_/A sky130_fd_sc_hd__or2_2
XFILLER_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09083_ _09764_/A vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06295_ _10922_/Q _10905_/Q vssd1 vssd1 vccd1 vccd1 _06416_/A sky130_fd_sc_hd__or2_1
X_08034_ _08034_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09985_ _09985_/A _10046_/A vssd1 vssd1 vccd1 vccd1 _10021_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08936_ _08936_/A vssd1 vssd1 vccd1 vccd1 _10832_/D sky130_fd_sc_hd__clkbuf_1
X_08867_ _08866_/A _08866_/B _08870_/D vssd1 vssd1 vccd1 vccd1 _08867_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07818_ _06145_/A _06258_/X _07807_/X _07817_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ hold20/A sky130_fd_sc_hd__o221ai_4
XFILLER_17_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08798_ _08803_/D _08798_/B vssd1 vssd1 vccd1 vccd1 _08798_/X sky130_fd_sc_hd__xor2_1
XFILLER_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10858__D _10858_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07749_ _09420_/A _07748_/A _07475_/C _07589_/B _07393_/Y vssd1 vssd1 vccd1 vccd1
+ _07750_/B sky130_fd_sc_hd__a311o_1
XFILLER_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ _10955_/CLK _10760_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10691_ _10845_/CLK _10691_/D vssd1 vssd1 vccd1 vccd1 _10691_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07810__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09419_ _09336_/A _09336_/B _09333_/A vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__a21o_1
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05968__C input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06145__B _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10044__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_6_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10935_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _09940_/B _10077_/A _10077_/B _10078_/A vssd1 vssd1 vccd1 vccd1 _10126_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10056_ _10123_/A _10122_/B _10056_/C vssd1 vssd1 vccd1 vccd1 _10057_/C sky130_fd_sc_hd__and3_1
XFILLER_48_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07704__B _09898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08088__A _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ _10958_/CLK _10958_/D vssd1 vssd1 vccd1 vccd1 _10958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10889_ _10889_/CLK _10889_/D vssd1 vssd1 vccd1 vccd1 _10889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06080_ _05744_/Y _07998_/A _07979_/A _05709_/Y vssd1 vssd1 vccd1 vccd1 _06080_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09770_ _09771_/A _09771_/B _09771_/C vssd1 vssd1 vccd1 vccd1 _09844_/B sky130_fd_sc_hd__o21ai_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06982_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__or2_4
X_05933_ _05859_/Y _05857_/B _08251_/A vssd1 vssd1 vccd1 vccd1 _05933_/X sky130_fd_sc_hd__a21o_1
X_08721_ _08888_/B vssd1 vssd1 vccd1 vccd1 _08902_/B sky130_fd_sc_hd__clkbuf_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _10798_/Q _10797_/Q _08648_/B _08592_/A vssd1 vssd1 vccd1 vccd1 _08652_/X
+ sky130_fd_sc_hd__a31o_1
X_05864_ _10698_/Q vssd1 vssd1 vccd1 vccd1 _08233_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07603_ _07603_/A _07711_/B vssd1 vssd1 vccd1 vccd1 _07604_/B sky130_fd_sc_hd__xnor2_4
X_05795_ _05732_/D _05734_/X _05732_/C vssd1 vssd1 vccd1 vccd1 _05795_/Y sky130_fd_sc_hd__a21oi_1
X_08583_ _08583_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _08583_/Y sky130_fd_sc_hd__nor2_1
X_07534_ _07534_/A _07534_/B _07534_/C vssd1 vssd1 vccd1 vccd1 _07535_/B sky130_fd_sc_hd__nor3_1
XFILLER_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ _07466_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07469_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08219__A1 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _08218_/A _07875_/A _09250_/A vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06416_ _06416_/A _06416_/B vssd1 vssd1 vccd1 vccd1 _06420_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07396_ _07396_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07397_/B sky130_fd_sc_hd__xnor2_2
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09135_ _09113_/X _09134_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09135_/Y sky130_fd_sc_hd__o21ai_1
X_06347_ _06561_/C vssd1 vssd1 vccd1 vccd1 _06547_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09066_ _05482_/X _08972_/A _08974_/A _09065_/X vssd1 vssd1 vccd1 vccd1 _09066_/X
+ sky130_fd_sc_hd__o211a_1
X_06278_ _10915_/Q _07102_/A vssd1 vssd1 vccd1 vccd1 _06558_/C sky130_fd_sc_hd__or2_1
XFILLER_135_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08017_ input31/X _08015_/X _08016_/X _08006_/X vssd1 vssd1 vccd1 vccd1 _10671_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ _10878_/Q _09572_/X _09967_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10878_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08919_ _10829_/Q _08919_/B vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__or2_1
XFILLER_92_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09899_ _09899_/A _09899_/B vssd1 vssd1 vccd1 vccd1 _09964_/A sky130_fd_sc_hd__xnor2_2
XFILLER_84_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10812_ _10819_/CLK _10812_/D vssd1 vssd1 vccd1 vccd1 _10812_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10743_ _10768_/CLK _10743_/D vssd1 vssd1 vccd1 vccd1 _10743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08355__B _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10674_ _10676_/CLK _10674_/D vssd1 vssd1 vccd1 vccd1 _10674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05995__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10108_ _09961_/A _10037_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _10109_/B sky130_fd_sc_hd__o21ai_1
XFILLER_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10039_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10141__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05580_ _05582_/B _05580_/B vssd1 vssd1 vccd1 vccd1 _05580_/X sky130_fd_sc_hd__and2_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07250_ _07250_/A _07250_/B vssd1 vssd1 vccd1 vccd1 _07515_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06201_ _06195_/X _06183_/X _06197_/Y _06200_/X vssd1 vssd1 vccd1 vccd1 _10597_/D
+ sky130_fd_sc_hd__o211a_1
X_07181_ _07229_/A _07398_/B _07181_/C vssd1 vssd1 vccd1 vccd1 _07183_/B sky130_fd_sc_hd__and3_1
XFILLER_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06132_ _10584_/Q vssd1 vssd1 vccd1 vccd1 _06134_/A sky130_fd_sc_hd__inv_2
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06063_ _05767_/Y _10675_/Q _08298_/A _05782_/Y vssd1 vssd1 vccd1 vccd1 _06063_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_99_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09822_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09753_ _09753_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09754_/B sky130_fd_sc_hd__xnor2_1
X_08704_ _08709_/A _08704_/B _08704_/C vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__nor3_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _07609_/A _07615_/A _06962_/X _07624_/A vssd1 vssd1 vccd1 vccd1 _06966_/B
+ sky130_fd_sc_hd__a31oi_4
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05916_ _05719_/A _05911_/Y _05913_/Y _08082_/C _05915_/X vssd1 vssd1 vccd1 vccd1
+ _05916_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09684_ _09684_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09685_/B sky130_fd_sc_hd__xnor2_2
XFILLER_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06896_ _06896_/A _06896_/B vssd1 vssd1 vccd1 vccd1 _06899_/B sky130_fd_sc_hd__nor2_4
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05847_ _10670_/Q vssd1 vssd1 vccd1 vccd1 _05851_/A sky130_fd_sc_hd__buf_2
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08635_ _08635_/A vssd1 vssd1 vccd1 vccd1 _10793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08566_ _10775_/Q _08578_/C vssd1 vssd1 vccd1 vccd1 _08567_/C sky130_fd_sc_hd__or2_1
XFILLER_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05778_ _10711_/Q vssd1 vssd1 vccd1 vccd1 _05778_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07517_ _07517_/A vssd1 vssd1 vccd1 vccd1 _09303_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08497_ _10784_/Q _08496_/X _08494_/X hold28/A vssd1 vssd1 vccd1 vccd1 _10747_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_71_clock _10985_/CLK vssd1 vssd1 vccd1 vccd1 _10842_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07448_ _07448_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07450_/A sky130_fd_sc_hd__xnor2_1
X_07379_ _07474_/B _07459_/B _07748_/B vssd1 vssd1 vccd1 vccd1 _07381_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09118_ _09118_/A vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _10936_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10390_/X sky130_fd_sc_hd__and2_1
X_09049_ _10934_/Q _10394_/C _10430_/B _10950_/Q vssd1 vssd1 vccd1 vccd1 _09049_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09226__S _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10652_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_73_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10486__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A io_wbs_m2s_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_39_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10854_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _10737_/CLK _10726_/D vssd1 vssd1 vccd1 vccd1 _10726_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_1_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10657_ _10657_/CLK _10657_/D vssd1 vssd1 vccd1 vccd1 _10657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10588_ _10813_/CLK _10588_/D vssd1 vssd1 vccd1 vccd1 _10588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06750_ _06758_/A _06776_/A vssd1 vssd1 vccd1 vccd1 _06771_/B sky130_fd_sc_hd__and2_1
XANTENNA__07164__B _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05701_ _08206_/A vssd1 vssd1 vccd1 vccd1 _05702_/A sky130_fd_sc_hd__inv_2
X_06681_ _06681_/A _06681_/B vssd1 vssd1 vccd1 vccd1 _06947_/B sky130_fd_sc_hd__or2_1
X_05632_ _10547_/Q _05636_/A vssd1 vssd1 vccd1 vccd1 _05632_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08420_ _06143_/X _08419_/B _08419_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10729_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05563_ _10570_/Q _10571_/Q _05576_/A vssd1 vssd1 vccd1 vccd1 _05566_/A sky130_fd_sc_hd__or3_1
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08282_ _08282_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08282_/X sky130_fd_sc_hd__or2_1
X_05494_ _05383_/X _05489_/X _05490_/X _05461_/D vssd1 vssd1 vccd1 vccd1 _10549_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_07302_ _07302_/A _07302_/B vssd1 vssd1 vccd1 vccd1 _07307_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07233_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07236_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07164_ _07166_/A _07164_/B vssd1 vssd1 vccd1 vccd1 _07196_/A sky130_fd_sc_hd__nand2_2
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06115_ _06115_/A _06115_/B vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07095_ _07284_/A _07095_/B vssd1 vssd1 vccd1 vccd1 _07096_/B sky130_fd_sc_hd__nand2_1
XFILLER_121_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06046_ _10663_/Q vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__buf_2
XFILLER_113_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input2_A io_qei_ch_a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07997_ _06206_/X _07987_/X _07996_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10663_/D
+ sky130_fd_sc_hd__o211a_1
X_09805_ _09805_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09856_/C sky130_fd_sc_hd__and2_1
XFILLER_101_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09736_ _09931_/A _09736_/B _09737_/A _09802_/C vssd1 vssd1 vccd1 vccd1 _09870_/A
+ sky130_fd_sc_hd__and4_1
X_06948_ _06948_/A _06948_/B vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__and2_1
XFILLER_67_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10468__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09667_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__nor2_1
X_08618_ _08600_/X _08597_/B _08623_/D _10789_/Q vssd1 vssd1 vccd1 vccd1 _08619_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06879_ _06881_/A _06881_/B _06878_/Y vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__o21a_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09560_/A _09560_/B _09597_/X vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__o21ai_1
X_08549_ _08549_/A vssd1 vssd1 vccd1 vccd1 _10770_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05647__A1 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10511_ _10529_/A vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10442_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10373_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09745__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09480__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05513__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ _10854_/CLK _10709_/D vssd1 vssd1 vccd1 vccd1 _10709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06063__A1 _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07920_ _10612_/Q _07906_/X _07910_/X _07919_/Y vssd1 vssd1 vccd1 vccd1 _07921_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_clkbuf_leaf_47_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07851_ _10577_/Q vssd1 vssd1 vccd1 vccd1 _07866_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput2 io_qei_ch_a vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07782_ _07782_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__xnor2_1
X_06802_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _06821_/A sky130_fd_sc_hd__xor2_2
X_09521_ _09520_/B _09520_/C _09520_/A vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__o21ai_1
X_06733_ _06752_/B _06752_/C vssd1 vssd1 vccd1 vccd1 _06745_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06118__A2 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__and2_1
X_06664_ _06695_/A _06695_/B _06661_/A vssd1 vssd1 vccd1 vccd1 _06665_/B sky130_fd_sc_hd__a21oi_2
XFILLER_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05615_ _10555_/Q _05664_/A vssd1 vssd1 vccd1 vccd1 _05615_/Y sky130_fd_sc_hd__xnor2_1
X_08403_ _08408_/A _10758_/Q vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__or2_1
XFILLER_51_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _09383_/A vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06595_ _06607_/B _06607_/C _06607_/A vssd1 vssd1 vccd1 vccd1 _06599_/B sky130_fd_sc_hd__a21boi_1
X_08334_ _08027_/A _08058_/X _08333_/X _06011_/X vssd1 vssd1 vccd1 vccd1 _08334_/X
+ sky130_fd_sc_hd__o211a_1
X_05546_ _05652_/A _05546_/B vssd1 vssd1 vccd1 vccd1 _05637_/B sky130_fd_sc_hd__or2_1
XFILLER_51_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05477_ _05643_/A vssd1 vssd1 vccd1 vccd1 _05912_/B sky130_fd_sc_hd__buf_2
X_08265_ _08267_/A _08277_/C vssd1 vssd1 vccd1 vccd1 _08276_/B sky130_fd_sc_hd__and2_1
X_08196_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08196_/X sky130_fd_sc_hd__and2_1
X_07216_ _07222_/A _07216_/B vssd1 vssd1 vccd1 vccd1 _07217_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07147_ _07147_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07309_/B sky130_fd_sc_hd__xor2_1
XFILLER_126_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07078_ _07167_/B vssd1 vssd1 vccd1 vccd1 _07163_/B sky130_fd_sc_hd__clkinv_2
X_06029_ _10412_/A _08157_/A _10351_/A _10578_/Q vssd1 vssd1 vccd1 vccd1 _06029_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10504__A _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08200__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _09599_/A _09760_/B _09903_/A _09805_/A vssd1 vssd1 vccd1 vccd1 _09719_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08644__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10425_ _06202_/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__a21bo_1
XFILLER_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10356_ _10351_/X _06752_/B _10355_/X _10923_/Q vssd1 vssd1 vccd1 vccd1 _10923_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10287_ _10287_/A _10287_/B _10287_/C _10287_/D vssd1 vssd1 vccd1 vccd1 _10289_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08819__A _08819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B2 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05400_ _05400_/A _05400_/B vssd1 vssd1 vccd1 vccd1 _05485_/A sky130_fd_sc_hd__xnor2_2
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06380_ _06896_/A _06381_/C vssd1 vssd1 vccd1 vccd1 _06394_/A sky130_fd_sc_hd__nor2_1
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05331_ _10673_/Q vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__09369__B _10905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08050_ _10369_/A _08971_/B _08416_/A _10583_/Q vssd1 vssd1 vccd1 vccd1 _08124_/A
+ sky130_fd_sc_hd__a31o_2
X_07001_ _07574_/A _07439_/A vssd1 vssd1 vccd1 vccd1 _07573_/C sky130_fd_sc_hd__nand2_2
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _10341_/B _09016_/B vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__nor2_1
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07903_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07903_/Y sky130_fd_sc_hd__clkinv_2
X_08883_ _08883_/A _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08883_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_69_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07834_ _07827_/X _05462_/C _07823_/X _07833_/Y vssd1 vssd1 vccd1 vccd1 _10621_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07765_ _10504_/A _07767_/B _06860_/B _06859_/A vssd1 vssd1 vccd1 vccd1 _07769_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07696_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _07696_/X sky130_fd_sc_hd__or2b_1
X_06716_ _06876_/B _06876_/A vssd1 vssd1 vccd1 vccd1 _07794_/A sky130_fd_sc_hd__or2b_1
X_09504_ _09676_/B _09444_/A _09444_/B _09361_/A vssd1 vssd1 vccd1 vccd1 _09507_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ _09471_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09477_/B sky130_fd_sc_hd__xnor2_2
X_06647_ _06647_/A _06647_/B vssd1 vssd1 vccd1 vccd1 _06648_/B sky130_fd_sc_hd__or2_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08249__C1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06578_ _06578_/A _06578_/B _06578_/C vssd1 vssd1 vccd1 vccd1 _06581_/B sky130_fd_sc_hd__and3_1
X_09366_ _09676_/B _09444_/A _09444_/B _09361_/A _09506_/B vssd1 vssd1 vccd1 vccd1
+ _09546_/B sky130_fd_sc_hd__a311o_1
X_05529_ _10572_/Q vssd1 vssd1 vccd1 vccd1 _05564_/A sky130_fd_sc_hd__inv_2
X_08317_ _08317_/A _08317_/B vssd1 vssd1 vccd1 vccd1 _08317_/Y sky130_fd_sc_hd__nand2_1
X_09297_ _10679_/Q _09296_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08248_ _08248_/A vssd1 vssd1 vccd1 vccd1 _08248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08179_ _08191_/B _08178_/X _06117_/D vssd1 vssd1 vccd1 vccd1 _08179_/Y sky130_fd_sc_hd__a21oi_1
X_10210_ _10202_/X _10203_/X _10208_/X _09480_/X vssd1 vssd1 vccd1 vccd1 _10210_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09295__A _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07808__A _07849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _10484_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05328__A _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__and2_1
XFILLER_87_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08724__B1 _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10974_ _10976_/CLK _10974_/D vssd1 vssd1 vccd1 vccd1 _10974_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10408_ _10408_/A vssd1 vssd1 vccd1 vccd1 _10408_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_125_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10339_ _10337_/Y _10338_/X _07539_/A _10192_/X vssd1 vssd1 vccd1 vccd1 _10913_/D
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05880_ _10655_/Q _10654_/Q _06038_/A _05906_/A vssd1 vssd1 vccd1 vccd1 _05900_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_93_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07550_ _07743_/B _07550_/B vssd1 vssd1 vccd1 vccd1 _07586_/A sky130_fd_sc_hd__or2_2
XFILLER_19_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06501_ _06517_/A _06489_/B _06506_/B _06758_/B vssd1 vssd1 vccd1 vccd1 _06503_/A
+ sky130_fd_sc_hd__a22oi_1
X_09220_ _08233_/A _07882_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__mux2_1
X_07481_ _07489_/A _07481_/B vssd1 vssd1 vccd1 vccd1 _07482_/B sky130_fd_sc_hd__and2_1
XFILLER_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08284__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06432_ _06645_/A _06433_/B vssd1 vssd1 vccd1 vccd1 _06434_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09151_ _10809_/Q _08985_/X _08988_/X _10722_/Q _09150_/X vssd1 vssd1 vccd1 vccd1
+ _09151_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10964__D _10964_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06363_ _06576_/B vssd1 vssd1 vccd1 vccd1 _06460_/B sky130_fd_sc_hd__clkbuf_2
X_08102_ _08098_/A _08098_/B _05728_/X vssd1 vssd1 vccd1 vccd1 _08102_/Y sky130_fd_sc_hd__o21ai_1
X_05314_ _10677_/Q _10676_/Q _05831_/B vssd1 vssd1 vccd1 vccd1 _05827_/A sky130_fd_sc_hd__or3_1
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09082_ _10969_/Q vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08033_ input39/X _07985_/B _08032_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06294_ _10904_/Q vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_115_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06251__B _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09984_ _09918_/A _09918_/B _09916_/A vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__a21oi_1
X_08935_ _08935_/A _10831_/Q vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__and2_1
XANTENNA__08706__B1 _08674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08182__A1 _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ _08866_/A _08866_/B _08870_/D vssd1 vssd1 vccd1 vccd1 _08866_/X sky130_fd_sc_hd__and3_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08797_ _10813_/Q _08815_/B _08792_/Y vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__a21bo_1
X_07817_ _10868_/Q _07824_/B vssd1 vssd1 vccd1 vccd1 _07817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07748_ _07748_/A _07748_/B vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07679_ _09303_/B _07249_/B _07519_/B vssd1 vssd1 vccd1 vccd1 _07680_/B sky130_fd_sc_hd__a21bo_1
X_10690_ _10845_/CLK _10690_/D vssd1 vssd1 vccd1 vccd1 _10690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09418_ _09418_/A vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__08237__A2 _08061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ _07013_/A _10891_/Q vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__and2b_1
XFILLER_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06248__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input40_A io_wbs_m2s_data[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10124_ _10124_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10055_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10091_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08369__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10957_ _10958_/CLK _10957_/D vssd1 vssd1 vccd1 vccd1 _10957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10888_ _10889_/CLK _10888_/D vssd1 vssd1 vccd1 vccd1 _10888_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_129_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _07098_/A _07102_/A vssd1 vssd1 vccd1 vccd1 _07747_/B sky130_fd_sc_hd__or2_2
X_05932_ _08224_/A _05870_/X _05866_/X _08233_/A _05931_/X vssd1 vssd1 vccd1 vccd1
+ _05932_/X sky130_fd_sc_hd__o221a_1
X_08720_ _08840_/B vssd1 vssd1 vccd1 vccd1 _08888_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05863_ _05863_/A _05863_/B vssd1 vssd1 vccd1 vccd1 _05863_/X sky130_fd_sc_hd__and2_1
XFILLER_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08651_ _10798_/Q vssd1 vssd1 vccd1 vccd1 _08651_/Y sky130_fd_sc_hd__inv_2
X_07602_ _07502_/A _07502_/B _07455_/A vssd1 vssd1 vccd1 vccd1 _07711_/B sky130_fd_sc_hd__o21ai_2
XFILLER_26_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05794_ _05794_/A _05794_/B vssd1 vssd1 vccd1 vccd1 _05794_/Y sky130_fd_sc_hd__nor2_1
X_08582_ _10780_/Q _08585_/C vssd1 vssd1 vccd1 vccd1 _08583_/B sky130_fd_sc_hd__and2_1
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07533_ _07623_/A _07622_/B vssd1 vssd1 vccd1 vccd1 _07617_/B sky130_fd_sc_hd__or2_1
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07464_ _07464_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _07466_/B sky130_fd_sc_hd__nor2_1
X_09203_ _09203_/A vssd1 vssd1 vccd1 vccd1 _09203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06415_ _10922_/Q _07083_/A vssd1 vssd1 vccd1 vccd1 _06416_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08219__A2 _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05788__D _05802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _09114_/X _09133_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__o21a_1
XFILLER_50_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07395_ _07393_/Y _07394_/X _07386_/B vssd1 vssd1 vccd1 vccd1 _07594_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__07978__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06346_ _06346_/A _06346_/B vssd1 vssd1 vccd1 vccd1 _06561_/C sky130_fd_sc_hd__nand2_1
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09065_ _06038_/X _08995_/X _09064_/X _08981_/A vssd1 vssd1 vccd1 vccd1 _09065_/X
+ sky130_fd_sc_hd__a211o_1
X_06277_ _10898_/Q vssd1 vssd1 vccd1 vccd1 _07102_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08016_ _08289_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08016_/X sky130_fd_sc_hd__or2_1
XFILLER_89_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09967_/Y sky130_fd_sc_hd__xnor2_1
X_08918_ _10829_/Q _08918_/B vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07805__B _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__xnor2_1
X_08849_ _08846_/X _08848_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10819_/D sky130_fd_sc_hd__a21oi_1
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10811_ _10811_/CLK _10811_/D vssd1 vssd1 vccd1 vccd1 _10811_/Q sky130_fd_sc_hd__dfxtp_1
X_10742_ _10791_/CLK _10742_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ _10673_/CLK _10673_/D vssd1 vssd1 vccd1 vccd1 _10673_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09407__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06172__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10107_ _10107_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__xor2_4
X_10038_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09930__B _09930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06200_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06200_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07180_ _07197_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07181_/C sky130_fd_sc_hd__nand2_1
XFILLER_118_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06131_ _06204_/B vssd1 vssd1 vccd1 vccd1 _06131_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06062_ _08282_/A _05851_/A _05388_/A _05726_/A _06061_/X vssd1 vssd1 vccd1 vccd1
+ _06062_/X sky130_fd_sc_hd__a221o_1
XFILLER_117_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07906__A _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _09754_/A _09754_/B _09757_/B vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__o21ba_1
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09752_ _09684_/A _09683_/B _09961_/A vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08703_ _08709_/A _08704_/B _08704_/C vssd1 vssd1 vccd1 vccd1 _08705_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _07662_/A vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__buf_2
X_05915_ _05408_/Y _05912_/B _05813_/X _05914_/X vssd1 vssd1 vccd1 vccd1 _05915_/X
+ sky130_fd_sc_hd__a31o_1
X_09683_ _10066_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__nor2_1
X_06895_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _06896_/B sky130_fd_sc_hd__nor2_1
X_05846_ _10671_/Q vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__buf_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08737__A _08837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_5_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10955_/CLK sky130_fd_sc_hd__clkbuf_16
X_08634_ _08638_/C _08634_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _08635_/A sky130_fd_sc_hd__and3b_1
X_05777_ _06113_/A _10570_/Q _10569_/Q _05766_/Y vssd1 vssd1 vccd1 vccd1 _05785_/A
+ sky130_fd_sc_hd__o22a_1
X_08565_ _10251_/S _10775_/Q _08565_/C vssd1 vssd1 vccd1 vccd1 _08565_/X sky130_fd_sc_hd__and3_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07516_ _07516_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__and2_1
XFILLER_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06257__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08496_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08496_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07447_ _07447_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07448_/B sky130_fd_sc_hd__or2_1
XFILLER_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07378_ _07728_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07378_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08073__B1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ _10939_/Q _09008_/X _09116_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09117_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06329_ _10913_/Q vssd1 vssd1 vccd1 vccd1 _07112_/A sky130_fd_sc_hd__buf_2
XFILLER_136_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09048_ _10369_/B vssd1 vssd1 vccd1 vccd1 _10394_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_124_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06167__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _10737_/CLK _10725_/D vssd1 vssd1 vccd1 vccd1 _10725_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10656_ _10657_/CLK _10656_/D vssd1 vssd1 vccd1 vccd1 _10656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10587_ _10813_/CLK _10587_/D vssd1 vssd1 vccd1 vccd1 _10587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07726__A _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05700_ _10695_/Q vssd1 vssd1 vccd1 vccd1 _08206_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06680_ _06680_/A _06680_/B vssd1 vssd1 vccd1 vccd1 _06681_/B sky130_fd_sc_hd__and2_1
X_05631_ _10687_/Q _05631_/B vssd1 vssd1 vccd1 vccd1 _05631_/X sky130_fd_sc_hd__or2_1
XANTENNA__08557__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08350_ _08350_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08350_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05562_ _10569_/Q _10568_/Q _05769_/A _05582_/B vssd1 vssd1 vccd1 vccd1 _05576_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA_clkbuf_leaf_43_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07301_ _07301_/A _07344_/A vssd1 vssd1 vccd1 vccd1 _07302_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08281_ _08263_/X _08276_/Y _08295_/C _08280_/X _08062_/X vssd1 vssd1 vccd1 vccd1
+ _08281_/X sky130_fd_sc_hd__o32a_1
X_05493_ _05385_/Y _05489_/X _05490_/X _05462_/A vssd1 vssd1 vccd1 vccd1 _10548_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07232_ _07232_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07163_ _07415_/A _07163_/B _07186_/C vssd1 vssd1 vccd1 vccd1 _07193_/A sky130_fd_sc_hd__or3_1
X_06114_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _06115_/B sky130_fd_sc_hd__or2_1
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10401__A2 _10719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07094_ _07284_/A _07095_/B vssd1 vssd1 vccd1 vccd1 _07363_/C sky130_fd_sc_hd__or2_1
X_06045_ _06045_/A _06045_/B vssd1 vssd1 vccd1 vccd1 _06045_/X sky130_fd_sc_hd__or2_1
XANTENNA__06081__A2 _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _09870_/B _09804_/B vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__and2b_1
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07996_ _08209_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _07996_/X sky130_fd_sc_hd__or2_1
XFILLER_86_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09735_ _09735_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09802_/C sky130_fd_sc_hd__xor2_1
X_06947_ _06947_/A _06947_/B vssd1 vssd1 vccd1 vccd1 _06948_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09666_ _09621_/A _09621_/B _09624_/A vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08617_ _10789_/Q _08617_/B _08623_/D vssd1 vssd1 vccd1 vccd1 _08617_/X sky130_fd_sc_hd__and3_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06878_ _06878_/A _06878_/B vssd1 vssd1 vccd1 vccd1 _06878_/Y sky130_fd_sc_hd__nand2_1
X_05829_ _05318_/A _05831_/C _05827_/Y _08032_/A vssd1 vssd1 vccd1 vccd1 _05829_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09597_ _09597_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__or2_1
X_08548_ _08580_/B _08548_/B _08553_/B vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__and3_1
XFILLER_70_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08479_ _10780_/Q _10743_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10510_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__or2_1
X_10441_ _10441_/A vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__buf_2
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10372_ _06124_/A _10371_/X _10408_/A vssd1 vssd1 vccd1 vccd1 _10372_/X sky130_fd_sc_hd__a21bo_1
XFILLER_136_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ _10854_/CLK _10708_/D vssd1 vssd1 vccd1 vccd1 _10708_/Q sky130_fd_sc_hd__dfxtp_1
X_10639_ _10830_/CLK _10639_/D vssd1 vssd1 vccd1 vccd1 _10639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06063__A2 _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07850_ _07850_/A vssd1 vssd1 vccd1 vccd1 _07850_/X sky130_fd_sc_hd__buf_4
XFILLER_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07012__A1 _06997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07781_ _10502_/A _06857_/B _07780_/X _07635_/A vssd1 vssd1 vccd1 vccd1 _07782_/B
+ sky130_fd_sc_hd__a22o_1
X_06801_ _10510_/A _06842_/A vssd1 vssd1 vccd1 vccd1 _07774_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_70_clock _10985_/CLK vssd1 vssd1 vccd1 vccd1 _10986_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09520_ _09520_/A _09520_/B _09520_/C vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__or3_1
X_06732_ _06732_/A _06732_/B vssd1 vssd1 vccd1 vccd1 _06752_/C sky130_fd_sc_hd__nand2_1
Xinput3 io_qei_ch_b vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_6
XFILLER_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10967__D _10967_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06663_ _06663_/A _06663_/B vssd1 vssd1 vccd1 vccd1 _06695_/B sky130_fd_sc_hd__xnor2_2
X_09451_ _09489_/A _09451_/B _09579_/A vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__and3_1
X_05614_ _10554_/Q _05663_/B vssd1 vssd1 vccd1 vccd1 _05664_/A sky130_fd_sc_hd__nor2_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08402_ _08397_/X _10741_/Q _08394_/X _08401_/X vssd1 vssd1 vccd1 vccd1 _10723_/D
+ sky130_fd_sc_hd__o211a_1
X_09382_ _09431_/A _09431_/B vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__xnor2_1
X_06594_ _06594_/A _06594_/B _06579_/Y vssd1 vssd1 vccd1 vccd1 _06607_/A sky130_fd_sc_hd__or3b_1
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08333_ _08333_/A _08333_/B _08038_/A vssd1 vssd1 vccd1 vccd1 _08333_/X sky130_fd_sc_hd__or3b_1
X_05545_ _05652_/B _05652_/C vssd1 vssd1 vccd1 vccd1 _05546_/B sky130_fd_sc_hd__nor2_1
X_08264_ _08277_/B vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05476_ _10616_/Q _05471_/X _05474_/Y _05475_/X vssd1 vssd1 vccd1 vccd1 _10541_/D
+ sky130_fd_sc_hd__a22o_1
X_08195_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__nor2_1
X_07215_ _07248_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07250_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07146_ _07148_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07309_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06054__A2 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clock _10857_/CLK vssd1 vssd1 vccd1 vccd1 _10654_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_106_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07077_ _07151_/A _07390_/B _07375_/A vssd1 vssd1 vccd1 vccd1 _07091_/B sky130_fd_sc_hd__a21boi_1
XFILLER_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06028_ _08489_/A vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10705_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07979_ _07979_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07979_/X sky130_fd_sc_hd__or2_1
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09718_ _09930_/B _09903_/A vssd1 vssd1 vccd1 vccd1 _09718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ _09619_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__and2b_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08082__D _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08660__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _10945_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10424_/X sky130_fd_sc_hd__and2_1
XFILLER_124_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10377__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10355_ _10355_/A vssd1 vssd1 vccd1 vccd1 _10355_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10301_/A _10300_/A vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05330_ _10641_/Q vssd1 vssd1 vccd1 vccd1 _07907_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07000_ _09920_/B _07000_/B vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__xnor2_1
XFILLER_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08951_ _09126_/A _09142_/D vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__or2_1
X_07902_ _07916_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _10639_/D sky130_fd_sc_hd__nor2_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08882_ _10824_/Q _08888_/B vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__xor2_1
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07833_ _06160_/A _07828_/X _07829_/X _07831_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07833_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07764_ _07764_/A _07764_/B vssd1 vssd1 vccd1 vccd1 _07803_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08497__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09503_ _09448_/A _09879_/B _09678_/A vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__o21ai_2
X_06715_ _06715_/A _06721_/A vssd1 vssd1 vccd1 vccd1 _06876_/A sky130_fd_sc_hd__xnor2_1
X_07695_ _07693_/A _07693_/B _09576_/A vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__a21bo_1
XFILLER_80_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09434_ _10066_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__nor2_1
X_06646_ _06646_/A _06646_/B vssd1 vssd1 vccd1 vccd1 _06647_/B sky130_fd_sc_hd__and2_1
XFILLER_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08249__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09365_ _10887_/Q _10903_/Q vssd1 vssd1 vccd1 vccd1 _09506_/B sky130_fd_sc_hd__and2b_1
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06577_ _06578_/A _06578_/B _06578_/C vssd1 vssd1 vccd1 vccd1 _06581_/C sky130_fd_sc_hd__a21oi_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05528_ _05528_/A vssd1 vssd1 vccd1 vccd1 _05528_/X sky130_fd_sc_hd__clkbuf_4
X_08316_ _08305_/A _08315_/C _08317_/A vssd1 vssd1 vccd1 vccd1 _08316_/Y sky130_fd_sc_hd__a21oi_1
X_09296_ _06115_/A _10647_/Q _09296_/S vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _08243_/A _08251_/C _08246_/Y vssd1 vssd1 vccd1 vccd1 _08247_/Y sky130_fd_sc_hd__a21oi_1
X_05459_ _05453_/A _09107_/A _09078_/A _05455_/X _05458_/X vssd1 vssd1 vccd1 vccd1
+ _05459_/X sky130_fd_sc_hd__a221o_1
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08178_ _08173_/A _08173_/B _08181_/A vssd1 vssd1 vccd1 vccd1 _08178_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08480__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10515__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07129_ _10985_/Q _07229_/B _07376_/A vssd1 vssd1 vccd1 vccd1 _07133_/B sky130_fd_sc_hd__a21boi_2
XFILLER_121_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _10482_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10071_ _10482_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__and2_1
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10973_ _10976_/CLK _10973_/D vssd1 vssd1 vccd1 vccd1 _10973_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10407_ _10389_/X _10721_/Q _10405_/X _10406_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10940_/D sky130_fd_sc_hd__o221a_1
XFILLER_112_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10338_ _10336_/X _10332_/X _10333_/Y _09480_/X vssd1 vssd1 vccd1 vccd1 _10338_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05777__B2 _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08176__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10269_ _10252_/A _10247_/A _10261_/A _10268_/Y vssd1 vssd1 vccd1 vccd1 _10287_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07518__A2 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07480_ _07480_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__xnor2_1
X_06500_ _06502_/B vssd1 vssd1 vccd1 vccd1 _06758_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08565__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06431_ _06431_/A _06431_/B vssd1 vssd1 vccd1 vccd1 _06433_/B sky130_fd_sc_hd__xor2_1
X_09150_ _07979_/A _09123_/X _09127_/X _09149_/X vssd1 vssd1 vccd1 vccd1 _09150_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06362_ _06587_/A vssd1 vssd1 vccd1 vccd1 _06576_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08101_ _08097_/X _08099_/X _08100_/X vssd1 vssd1 vccd1 vccd1 _10684_/D sky130_fd_sc_hd__o21a_1
X_05313_ _05329_/A vssd1 vssd1 vccd1 vccd1 _05831_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09081_ _08974_/X _09077_/X _09078_/Y _09036_/X _09080_/X vssd1 vssd1 vccd1 vccd1
+ _09081_/X sky130_fd_sc_hd__a32o_1
X_06293_ _06293_/A _06293_/B vssd1 vssd1 vccd1 vccd1 _06805_/A sky130_fd_sc_hd__nor2_2
X_08032_ _08032_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09396__A _09396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput50 io_wbs_m2s_we vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05768__A1 _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09983_ _09983_/A _09983_/B vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10210__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05768__B2 _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ _08934_/A vssd1 vssd1 vccd1 vccd1 _10831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08167__C1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__B2 _08701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08706__A1 _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08865_ _10822_/Q _08865_/B vssd1 vssd1 vccd1 vccd1 _08870_/D sky130_fd_sc_hd__xor2_1
XFILLER_69_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07816_ _06255_/X _08994_/A _06257_/X _07815_/Y vssd1 vssd1 vccd1 vccd1 _10617_/D
+ sky130_fd_sc_hd__o211a_1
X_08796_ _10814_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08803_/D sky130_fd_sc_hd__xor2_1
XFILLER_84_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07747_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07748_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07678_ _07678_/A _09303_/B vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__nand2_1
X_09417_ _09417_/A _09810_/A vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__or2_1
XFILLER_12_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06629_ _06800_/A _06719_/C vssd1 vssd1 vccd1 vccd1 _06630_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09348_ _10891_/Q _10907_/Q vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _09289_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09280_/A sky130_fd_sc_hd__and2_1
XFILLER_4_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09198__B2 _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__nand2_1
XFILLER_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input33_A io_wbs_m2s_data[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10054_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__or2_1
XFILLER_36_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08330__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08385__A _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ _10956_/CLK _10956_/D vssd1 vssd1 vccd1 vccd1 _10956_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05802__A _05802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10887_ _10889_/CLK _10887_/D vssd1 vssd1 vccd1 vccd1 _10887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07436__A1 _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07436__B2 _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__A _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _10899_/Q vssd1 vssd1 vccd1 vccd1 _07098_/A sky130_fd_sc_hd__clkbuf_2
X_05931_ _08218_/A _05872_/X _05870_/X _08224_/A _05930_/X vssd1 vssd1 vccd1 vccd1
+ _05931_/X sky130_fd_sc_hd__a221o_1
XFILLER_100_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05862_ _05350_/B _05854_/B _08244_/A vssd1 vssd1 vccd1 vccd1 _05863_/A sky130_fd_sc_hd__o21ai_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08650_ _08650_/A vssd1 vssd1 vccd1 vccd1 _10797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07601_ _07601_/A _07601_/B vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__xnor2_4
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05793_ _05732_/B _05741_/Y _05742_/B vssd1 vssd1 vccd1 vccd1 _05794_/B sky130_fd_sc_hd__a21oi_1
X_08581_ _08581_/A vssd1 vssd1 vccd1 vccd1 _10779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06808__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07532_ _07628_/A _07627_/B vssd1 vssd1 vccd1 vccd1 _07622_/B sky130_fd_sc_hd__or2_1
XFILLER_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07463_ _07473_/A _07463_/B vssd1 vssd1 vccd1 vccd1 _07464_/B sky130_fd_sc_hd__and2_1
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09202_ _09202_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _10849_/D sky130_fd_sc_hd__nor2_4
X_06414_ _10905_/Q vssd1 vssd1 vccd1 vccd1 _07083_/A sky130_fd_sc_hd__buf_2
X_09133_ _10940_/Q _09008_/X _09132_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09133_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_07394_ _07394_/A vssd1 vssd1 vccd1 vccd1 _07394_/X sky130_fd_sc_hd__buf_2
XFILLER_136_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06345_ _06343_/A _06736_/A _06371_/C vssd1 vssd1 vccd1 vccd1 _06346_/B sky130_fd_sc_hd__o21ai_1
X_09064_ _05462_/C _08978_/A _06129_/B _05728_/X _09179_/A vssd1 vssd1 vccd1 vccd1
+ _09064_/X sky130_fd_sc_hd__o221a_1
X_06276_ _06276_/A _06276_/B vssd1 vssd1 vccd1 vccd1 _06352_/A sky130_fd_sc_hd__nand2_1
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08015_ _08015_/A vssd1 vssd1 vccd1 vccd1 _08015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_38_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _09893_/Y _09896_/B _09894_/A vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__a21o_1
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08917_ _08814_/X _08915_/Y _08916_/X vssd1 vssd1 vccd1 vccd1 _10828_/D sky130_fd_sc_hd__o21a_1
X_09897_ _10877_/Q _09572_/X _09896_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10877_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07805__C _10117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08848_ input28/X _08672_/X _08674_/X _08847_/X vssd1 vssd1 vccd1 vccd1 _08848_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06166__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08779_ _06191_/X _08728_/X _08729_/X _08771_/A vssd1 vssd1 vccd1 vccd1 _08779_/X
+ sky130_fd_sc_hd__a22o_1
X_10810_ _10813_/CLK _10810_/D vssd1 vssd1 vccd1 vccd1 _10810_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10741_ _10791_/CLK _10741_/D vssd1 vssd1 vccd1 vccd1 _10741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10672_ _10673_/CLK _10672_/D vssd1 vssd1 vccd1 vccd1 _10672_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08933__A _08935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10106_ _10035_/A _10035_/B _10105_/X vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__a21o_2
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07715__C _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05770__A1_N _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ _10037_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06157__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10939_ _10955_/CLK _10939_/D vssd1 vssd1 vccd1 vccd1 _10939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06130_ _06149_/A vssd1 vssd1 vccd1 vccd1 _06204_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__07459__A _09304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06061_ _06061_/A _08000_/A vssd1 vssd1 vccd1 vccd1 _06061_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08909__A1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A0 _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06810__B _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09751_ _10066_/A vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06963_ _07675_/A vssd1 vssd1 vccd1 vccd1 _07662_/A sky130_fd_sc_hd__clkbuf_2
X_05914_ _10681_/Q _05913_/Y _05814_/X vssd1 vssd1 vccd1 vccd1 _05914_/X sky130_fd_sc_hd__a21bo_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08702_ _08691_/B _08693_/B _08689_/Y vssd1 vssd1 vccd1 vccd1 _08704_/C sky130_fd_sc_hd__a21o_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ _09682_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06894_ _06894_/A _06894_/B vssd1 vssd1 vccd1 vccd1 _06899_/A sky130_fd_sc_hd__xor2_4
X_05845_ _05845_/A _05941_/B vssd1 vssd1 vccd1 vccd1 _05940_/B sky130_fd_sc_hd__and2_1
XFILLER_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08633_ _08633_/A vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__buf_2
X_05776_ _08297_/A _05772_/Y _05564_/A _06115_/A _05807_/A vssd1 vssd1 vccd1 vccd1
+ _05786_/C sky130_fd_sc_hd__o221a_1
X_08564_ _10774_/Q _08559_/X _08562_/X _08563_/X vssd1 vssd1 vccd1 vccd1 _10774_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07515_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07516_/B sky130_fd_sc_hd__or2_1
XFILLER_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08495_ _10783_/Q _08491_/X _08494_/X _10746_/Q vssd1 vssd1 vccd1 vccd1 _10746_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07446_ _07714_/S _07445_/B _07445_/C vssd1 vssd1 vccd1 vccd1 _07447_/B sky130_fd_sc_hd__a21oi_1
XFILLER_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07377_ _07377_/A vssd1 vssd1 vccd1 vccd1 _07728_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09116_ _10955_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09116_/Y sky130_fd_sc_hd__nor2_1
X_06328_ _06288_/X _06851_/A _06851_/B _06850_/A vssd1 vssd1 vccd1 vccd1 _06342_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__06084__B1 _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09047_ _10432_/A _09142_/C _09142_/D _10341_/B vssd1 vssd1 vccd1 vccd1 _10369_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06259_ _10978_/Q vssd1 vssd1 vccd1 vccd1 _06436_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09949_ _09949_/A vssd1 vssd1 vccd1 vccd1 _09949_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07832__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09089__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _10737_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _10724_/Q sky130_fd_sc_hd__dfxtp_1
X_10655_ _10657_/CLK _10655_/D vssd1 vssd1 vccd1 vccd1 _10655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08064__A1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10586_ _10808_/CLK _10586_/D vssd1 vssd1 vccd1 vccd1 _10586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05527__A _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05630_ _05630_/A _05630_/B vssd1 vssd1 vccd1 vccd1 _05631_/B sky130_fd_sc_hd__and2_1
XANTENNA__05889__B1 _05886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05561_ _10566_/Q _05588_/A vssd1 vssd1 vccd1 vccd1 _05582_/B sky130_fd_sc_hd__or2_1
X_07300_ _07349_/B _07300_/B vssd1 vssd1 vccd1 vccd1 _07307_/A sky130_fd_sc_hd__or2_1
X_08280_ _05851_/A _08235_/B _08278_/Y _08279_/X vssd1 vssd1 vccd1 vccd1 _08280_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05492_ _05389_/Y _05489_/X _05490_/X _05462_/B vssd1 vssd1 vccd1 vccd1 _10547_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07231_ _07231_/A _07231_/B vssd1 vssd1 vccd1 vccd1 _07258_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08055__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09252__A0 _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ _07211_/A _07166_/B vssd1 vssd1 vccd1 vccd1 _07186_/C sky130_fd_sc_hd__nand2_1
XFILLER_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06113_ _06113_/A _08333_/A vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08055__B2 _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07093_ _07363_/B _07093_/B vssd1 vssd1 vccd1 vccd1 _07095_/B sky130_fd_sc_hd__nand2_1
XFILLER_126_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06044_ _05749_/A _10671_/Q _05408_/Y _08082_/D vssd1 vssd1 vccd1 vccd1 _06045_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_114_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10343__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09803_ _10069_/A _09802_/B _09930_/C _09932_/A vssd1 vssd1 vccd1 vccd1 _09804_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07995_ _07995_/A vssd1 vssd1 vccd1 vccd1 _08005_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _09734_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09735_/B sky130_fd_sc_hd__xnor2_2
X_06946_ _06946_/A _06948_/A vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__xnor2_2
XFILLER_28_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09665_ _09665_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__xor2_1
XFILLER_27_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06877_ _06878_/A _06878_/B vssd1 vssd1 vccd1 vccd1 _06881_/B sky130_fd_sc_hd__xnor2_2
X_05828_ _10678_/Q vssd1 vssd1 vccd1 vccd1 _08032_/A sky130_fd_sc_hd__clkinv_2
XFILLER_70_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08616_ _08614_/Y _08612_/C _08623_/D _08617_/B _08630_/A vssd1 vssd1 vccd1 vccd1
+ _10788_/D sky130_fd_sc_hd__a221oi_1
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05759_ _06061_/A vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__inv_2
X_08547_ _08547_/A _08547_/B vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08483__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08478_ _08478_/A vssd1 vssd1 vccd1 vccd1 _10742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07429_ _07429_/A _07429_/B vssd1 vssd1 vccd1 vccd1 _07430_/B sky130_fd_sc_hd__nand2_1
X_10440_ _10950_/Q _10440_/B vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__or2_1
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _10371_/A vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10253__A _10253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07562__A _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06178__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_7_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10707_ _10707_/CLK _10707_/D vssd1 vssd1 vccd1 vccd1 _10707_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10638_ _10669_/CLK _10638_/D vssd1 vssd1 vccd1 vccd1 _10638_/Q sky130_fd_sc_hd__dfxtp_1
X_10569_ _10865_/CLK _10569_/D vssd1 vssd1 vccd1 vccd1 _10569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_4_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10946_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07780_ _06855_/A _07780_/B _07780_/C vssd1 vssd1 vccd1 vccd1 _07780_/X sky130_fd_sc_hd__and3b_1
X_06800_ _06800_/A vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06731_ _06731_/A _06731_/B vssd1 vssd1 vccd1 vccd1 _06752_/B sky130_fd_sc_hd__xnor2_4
Xinput4 io_wbs_m2s_addr[0] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
X_09450_ _09555_/A _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__and3_1
XFILLER_91_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08401_ _08408_/A _10757_/Q vssd1 vssd1 vccd1 vccd1 _08401_/X sky130_fd_sc_hd__or2_1
XFILLER_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06662_ _06692_/A _06692_/B _06621_/A vssd1 vssd1 vccd1 vccd1 _06663_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05613_ _10694_/Q vssd1 vssd1 vccd1 vccd1 _05877_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09381_ _09381_/A _10897_/Q vssd1 vssd1 vccd1 vccd1 _09431_/B sky130_fd_sc_hd__xor2_4
XFILLER_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06593_ _06593_/A _06593_/B _06593_/C vssd1 vssd1 vccd1 vccd1 _06607_/C sky130_fd_sc_hd__and3_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08332_ _08332_/A _08332_/B vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__and2_1
X_05544_ _05910_/B _05737_/B _05543_/Y vssd1 vssd1 vccd1 vccd1 _05652_/C sky130_fd_sc_hd__a21oi_1
X_08263_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08263_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10983__D _10983_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05475_ _10648_/Q vssd1 vssd1 vccd1 vccd1 _05475_/X sky130_fd_sc_hd__buf_4
X_07214_ _07214_/A _07214_/B vssd1 vssd1 vccd1 vccd1 _07232_/A sky130_fd_sc_hd__and2_1
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08194_ _08190_/X _08192_/X _08193_/X vssd1 vssd1 vccd1 vccd1 _10693_/D sky130_fd_sc_hd__o21a_1
XANTENNA__08028__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07145_ _07145_/A _07145_/B vssd1 vssd1 vccd1 vccd1 _07148_/B sky130_fd_sc_hd__xnor2_1
X_07076_ _07137_/A _07076_/B vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06027_ _08201_/A _09403_/B vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__and2_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08200__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _06178_/X _07965_/X _07976_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10657_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09717_ _09717_/A vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06929_ _06937_/A _06937_/B _06928_/Y vssd1 vssd1 vccd1 vccd1 _06936_/B sky130_fd_sc_hd__a21o_1
XFILLER_90_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09648_ _09649_/B _09619_/A vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__or2b_1
XFILLER_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ _10408_/X _10725_/Q _10421_/X _10422_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10944_/D sky130_fd_sc_hd__o221a_1
XFILLER_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ _09634_/A _06732_/B _08494_/X _10922_/Q vssd1 vssd1 vccd1 vccd1 _10922_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08727__C1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10285_ _10957_/Q _10941_/Q vssd1 vssd1 vccd1 vccd1 _10300_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09758__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08950_ _09142_/A _09142_/B vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__or2_1
X_07901_ _10607_/Q _07888_/X _07892_/X _07900_/Y vssd1 vssd1 vccd1 vccd1 _07902_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _10823_/D sky130_fd_sc_hd__nor2_1
XANTENNA__09682__A _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07832_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07941__A0 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07763_ _07763_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07764_/B sky130_fd_sc_hd__xnor2_1
X_09502_ _09501_/B _09501_/C _09501_/A vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08280__A2_N _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10190__B_N _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06714_ _06722_/A _06714_/B vssd1 vssd1 vccd1 vccd1 _06721_/A sky130_fd_sc_hd__xnor2_1
X_07694_ _09575_/B _09575_/C _09575_/A vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__o21ai_1
XFILLER_37_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07930__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__nor2_1
X_06645_ _06645_/A _06645_/B vssd1 vssd1 vccd1 vccd1 _06648_/A sky130_fd_sc_hd__or2_1
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08249__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09364_ _09336_/A _09336_/B _09421_/B _09333_/A vssd1 vssd1 vccd1 vccd1 _09444_/B
+ sky130_fd_sc_hd__a211o_1
X_08315_ _08315_/A _08315_/B _08315_/C vssd1 vssd1 vccd1 vccd1 _08327_/B sky130_fd_sc_hd__and3_1
XANTENNA__05450__A _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06576_ _10974_/Q _06576_/B _06951_/A vssd1 vssd1 vccd1 vccd1 _06578_/C sky130_fd_sc_hd__and3_1
XFILLER_138_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09295_ _09295_/A vssd1 vssd1 vccd1 vccd1 _10864_/D sky130_fd_sc_hd__clkbuf_1
X_05527_ _06115_/A vssd1 vssd1 vccd1 vccd1 _05528_/A sky130_fd_sc_hd__clkbuf_2
X_08246_ _08243_/A _08251_/C _08067_/X vssd1 vssd1 vccd1 vccd1 _08246_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__05468__D1 _05467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05458_ _05455_/X _09078_/A _05283_/Y _09020_/A _05457_/X vssd1 vssd1 vccd1 vccd1
+ _05458_/X sky130_fd_sc_hd__o221a_1
XFILLER_137_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08177_ _08172_/X _08174_/X _08176_/X vssd1 vssd1 vccd1 vccd1 _10691_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05389_ _05389_/A _05389_/B vssd1 vssd1 vccd1 vccd1 _05389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07128_ _07137_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _07376_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07059_ _07560_/A _07076_/B vssd1 vssd1 vccd1 vccd1 _07357_/C sky130_fd_sc_hd__nand2_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08724__A2 _08701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10531__A _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__A_N _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10972_ _10976_/CLK _10972_/D vssd1 vssd1 vccd1 vccd1 _10972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08655__B _08989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10406_ _06178_/X _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10406_/X sky130_fd_sc_hd__a21bo_1
XFILLER_124_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06191__A input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10337_ _10332_/X _10333_/Y _10336_/X vssd1 vssd1 vccd1 vccd1 _10337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _10268_/A vssd1 vssd1 vccd1 vccd1 _10268_/Y sky130_fd_sc_hd__inv_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10441__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ _10197_/Y _10198_/Y _09757_/A vssd1 vssd1 vccd1 vccd1 _10199_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06083__A2_N _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__B _10160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clock _10857_/CLK vssd1 vssd1 vccd1 vccd1 _10657_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06430_ _06631_/A _06430_/B vssd1 vssd1 vccd1 vccd1 _06431_/B sky130_fd_sc_hd__or2_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06366__A _10978_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06085__B _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06361_ _06281_/B _06359_/Y _06360_/X vssd1 vssd1 vccd1 vccd1 _06587_/A sky130_fd_sc_hd__o21a_1
X_08100_ _10531_/A _08047_/X _08052_/X _08098_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08100_/X sky130_fd_sc_hd__o221a_1
X_05312_ _10675_/Q _05834_/A vssd1 vssd1 vccd1 vccd1 _05329_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_37_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10702_/CLK sky130_fd_sc_hd__clkbuf_16
X_09080_ _10718_/Q _09079_/X _09037_/Y _10805_/Q vssd1 vssd1 vccd1 vccd1 _09080_/X
+ sky130_fd_sc_hd__a22o_1
X_06292_ _10927_/Q _06993_/A vssd1 vssd1 vccd1 vccd1 _06293_/B sky130_fd_sc_hd__nor2_1
Xinput40 io_wbs_m2s_data[31] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_6
X_08031_ input37/X _07985_/B _08029_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10677_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 reset vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_6
XFILLER_131_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09982_ _09982_/A _09982_/B vssd1 vssd1 vccd1 vccd1 _09983_/B sky130_fd_sc_hd__xnor2_1
X_08933_ _08935_/A input2/X vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__and2_1
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08706__A2 _08672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08864_ _08881_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _10821_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10351__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08795_ _08793_/X _08794_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10813_/D sky130_fd_sc_hd__o21a_1
XFILLER_84_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07815_ _06140_/A _06258_/X _07807_/X _07814_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07815_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07746_ _07746_/A _07746_/B vssd1 vssd1 vccd1 vccd1 _07755_/A sky130_fd_sc_hd__xnor2_1
XFILLER_65_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09416_ _10964_/Q _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__and3_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07677_ _07677_/A _07677_/B vssd1 vssd1 vccd1 vccd1 _07681_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_leaf_34_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06628_ _06841_/A _06408_/B _06409_/C vssd1 vssd1 vccd1 vccd1 _06633_/A sky130_fd_sc_hd__a21boi_1
X_09347_ _09863_/A _09797_/A vssd1 vssd1 vccd1 vccd1 _09372_/A sky130_fd_sc_hd__nand2_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06559_ _06281_/B _06359_/Y _06360_/X _06558_/X _06502_/B vssd1 vssd1 vccd1 vccd1
+ _07676_/A sky130_fd_sc_hd__o2111a_1
XFILLER_138_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _10826_/Q _09274_/X _09275_/X _09277_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09279_/B sky130_fd_sc_hd__a32o_1
X_08229_ _06117_/C _08074_/A _08228_/Y _08044_/A _08000_/A vssd1 vssd1 vccd1 vccd1
+ _08229_/X sky130_fd_sc_hd__a32o_1
XANTENNA__08491__A _08514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10526__A _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09198__A2 _09136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10122_ _10491_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _10148_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input26_A io_wbs_m2s_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07570__A _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10955_ _10955_/CLK _10955_/D vssd1 vssd1 vccd1 vccd1 _10955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10886_ _10889_/CLK _10886_/D vssd1 vssd1 vccd1 vccd1 _10886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09189__A2 _09136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05930_ _08206_/A _05876_/X _05872_/X _08224_/B _05929_/X vssd1 vssd1 vccd1 vccd1
+ _05930_/X sky130_fd_sc_hd__o221a_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05861_ _10667_/Q vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08580_ _08585_/C _08580_/B _08580_/C vssd1 vssd1 vccd1 vccd1 _08581_/A sky130_fd_sc_hd__and3b_1
XFILLER_82_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07600_ _07598_/Y _07451_/B _07599_/X vssd1 vssd1 vccd1 vccd1 _07601_/B sky130_fd_sc_hd__o21a_2
XFILLER_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05792_ _05747_/X _05761_/X _05749_/X vssd1 vssd1 vccd1 vccd1 _05792_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07531_ _07633_/A _07632_/B vssd1 vssd1 vccd1 vccd1 _07627_/B sky130_fd_sc_hd__or2_1
X_07462_ _07462_/A _07462_/B vssd1 vssd1 vccd1 vccd1 _07466_/A sky130_fd_sc_hd__nor2_1
XFILLER_34_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09201_ _09112_/A _09197_/Y _09200_/X vssd1 vssd1 vccd1 vccd1 _09202_/B sky130_fd_sc_hd__a21oi_1
X_07393_ _07592_/A vssd1 vssd1 vccd1 vccd1 _07393_/Y sky130_fd_sc_hd__clkinv_4
X_06413_ _06736_/A _06732_/A vssd1 vssd1 vccd1 vccd1 _06421_/A sky130_fd_sc_hd__nor2_1
X_09132_ _10956_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09132_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06344_ _06352_/C vssd1 vssd1 vccd1 vccd1 _06736_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09063_ _10717_/Q _08999_/X _09037_/Y _10804_/Q vssd1 vssd1 vccd1 vccd1 _09063_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10346__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06275_ _06275_/A _06275_/B vssd1 vssd1 vccd1 vccd1 _06276_/B sky130_fd_sc_hd__or2_1
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08014_ input30/X _08002_/X _08013_/Y _08006_/X vssd1 vssd1 vccd1 vccd1 _10670_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07358__C _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09965_ _09965_/A _09964_/X vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__or2b_1
XFILLER_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08916_ input37/X _08819_/X _08820_/X _10828_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08916_/X sky130_fd_sc_hd__o221a_1
X_09896_ _09896_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_57_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08847_ _10819_/Q vssd1 vssd1 vccd1 vccd1 _08847_/X sky130_fd_sc_hd__clkbuf_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08778_ _08778_/A _08778_/B _08778_/C vssd1 vssd1 vccd1 vccd1 _08778_/X sky130_fd_sc_hd__and3_1
XFILLER_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07390__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07729_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07730_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08863__A1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ _10836_/CLK _10740_/D vssd1 vssd1 vccd1 vccd1 _10740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ _10673_/CLK _10671_/D vssd1 vssd1 vccd1 vccd1 _10671_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08933__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09110__A _09228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08379__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09040__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10186__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ _10033_/B _10105_/B vssd1 vssd1 vccd1 vccd1 _10105_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10036_ _09961_/B _09962_/A _09961_/A vssd1 vssd1 vccd1 vccd1 _10037_/B sky130_fd_sc_hd__a21o_1
XFILLER_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05813__A _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10938_ _10955_/CLK _10938_/D vssd1 vssd1 vccd1 vccd1 _10938_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10869_ _10889_/CLK _10869_/D vssd1 vssd1 vccd1 vccd1 _10869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06060_ _08315_/A _08023_/A _08256_/A _05751_/Y _06059_/X vssd1 vssd1 vccd1 vccd1
+ _06070_/A sky130_fd_sc_hd__o221a_1
XFILLER_117_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08790__B1 _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _09815_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__or2_1
X_06962_ _07620_/A _06962_/B vssd1 vssd1 vccd1 vccd1 _06962_/X sky130_fd_sc_hd__and2_1
X_05913_ _05913_/A _05913_/B vssd1 vssd1 vccd1 vccd1 _05913_/Y sky130_fd_sc_hd__nand2_1
X_08701_ _08701_/A _08732_/B vssd1 vssd1 vccd1 vccd1 _08704_/B sky130_fd_sc_hd__nor2_1
X_09681_ _09681_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__xor2_2
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08632_ _08600_/X _08642_/D _10793_/Q vssd1 vssd1 vccd1 vccd1 _08634_/B sky130_fd_sc_hd__a21o_1
X_06893_ _06893_/A _06893_/B vssd1 vssd1 vccd1 vccd1 _06894_/B sky130_fd_sc_hd__xor2_4
X_05844_ _05844_/A _05844_/B _05844_/C vssd1 vssd1 vccd1 vccd1 _05941_/B sky130_fd_sc_hd__or3_1
XFILLER_94_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06819__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05775_ _06113_/A _10570_/Q _10571_/Q _08355_/A vssd1 vssd1 vccd1 vccd1 _05807_/A
+ sky130_fd_sc_hd__a22oi_1
X_08563_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08563_/X sky130_fd_sc_hd__buf_4
XANTENNA__10986__D _10986_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08494_ _10355_/A vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__buf_2
X_07514_ _07514_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__and2_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07445_ _07714_/S _07445_/B _07445_/C vssd1 vssd1 vccd1 vccd1 _07447_/A sky130_fd_sc_hd__and3_1
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07376_ _07376_/A vssd1 vssd1 vccd1 vccd1 _07459_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _09194_/B vssd1 vssd1 vccd1 vccd1 _09164_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06327_ _10929_/Q _10912_/Q vssd1 vssd1 vccd1 vccd1 _06850_/A sky130_fd_sc_hd__and2_1
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06084__B2 _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06258_ _07849_/A vssd1 vssd1 vccd1 vccd1 _06258_/X sky130_fd_sc_hd__buf_4
X_09046_ _09930_/B vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_123_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09022__A1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06189_ _06189_/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10168__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08781__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09948_ _09810_/B _09744_/B _09769_/B _10493_/A vssd1 vssd1 vccd1 vccd1 _09949_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09879_ _10129_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10274__B_N _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10798_/CLK _10723_/D vssd1 vssd1 vccd1 vccd1 _10723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10654_ _10654_/CLK _10654_/D vssd1 vssd1 vccd1 vccd1 _10654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08064__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10585_ _10813_/CLK _10585_/D vssd1 vssd1 vccd1 vccd1 _10585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_3_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10019_ _10089_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__and2_1
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05560_ _10565_/Q _10564_/Q _05593_/A vssd1 vssd1 vccd1 vccd1 _05588_/A sky130_fd_sc_hd__or3_1
XFILLER_91_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05491_ _05393_/B _05489_/X _05490_/X _05462_/C vssd1 vssd1 vccd1 vccd1 _10546_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07230_ _07231_/A _07231_/B vssd1 vssd1 vccd1 vccd1 _07230_/X sky130_fd_sc_hd__and2_1
XFILLER_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07161_ _10982_/Q vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__clkinv_2
X_06112_ _08339_/B _08332_/B vssd1 vssd1 vccd1 vccd1 _08333_/A sky130_fd_sc_hd__nor2_1
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07092_ _07402_/A _07091_/B _07091_/C vssd1 vssd1 vccd1 vccd1 _07093_/B sky130_fd_sc_hd__o21ai_1
X_06043_ _10680_/Q vssd1 vssd1 vccd1 vccd1 _08082_/D sky130_fd_sc_hd__buf_2
XFILLER_113_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09802_ _09931_/A _09802_/B _09802_/C _09932_/A vssd1 vssd1 vccd1 vccd1 _09870_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_115_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07994_ _06202_/X _07987_/X _07991_/Y _07993_/X vssd1 vssd1 vccd1 vccd1 _10662_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09733_ _09371_/B _09733_/B vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__and2b_1
X_06945_ _06945_/A _06945_/B vssd1 vssd1 vccd1 vccd1 _06946_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09664_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09728_/B sky130_fd_sc_hd__xor2_1
XFILLER_28_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06876_ _06876_/A _06876_/B vssd1 vssd1 vccd1 vccd1 _06878_/B sky130_fd_sc_hd__xnor2_1
X_05827_ _05827_/A _05831_/C vssd1 vssd1 vccd1 vccd1 _05827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08615_ _10788_/Q _10787_/Q _10786_/Q _10785_/Q vssd1 vssd1 vccd1 vccd1 _08623_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09595_ _09593_/Y _09595_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__and2b_1
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05758_ _08224_/A vssd1 vssd1 vccd1 vccd1 _06061_/A sky130_fd_sc_hd__clkbuf_4
X_08546_ _10769_/Q _08543_/B _10770_/Q vssd1 vssd1 vccd1 vccd1 _08548_/B sky130_fd_sc_hd__a21o_1
X_05689_ _05528_/X _05564_/Y _05687_/B _08350_/A _05688_/X vssd1 vssd1 vccd1 vccd1
+ _05689_/X sky130_fd_sc_hd__a221o_1
X_08477_ _08477_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08478_/A sky130_fd_sc_hd__or2_1
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07428_ _07428_/A _07428_/B _07428_/C vssd1 vssd1 vccd1 vccd1 _07429_/B sky130_fd_sc_hd__nand3_1
XFILLER_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07359_ _07359_/A _07359_/B vssd1 vssd1 vccd1 vccd1 _07407_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ _10399_/A vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09029_ _09716_/A vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__buf_2
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08939__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06459__A _10977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10706_ _10854_/CLK _10706_/D vssd1 vssd1 vccd1 vccd1 _10706_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09482__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10637_ _10669_/CLK _10637_/D vssd1 vssd1 vccd1 vccd1 _10637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10568_ _10865_/CLK _10568_/D vssd1 vssd1 vccd1 vccd1 _10568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08993__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ _06124_/X _10496_/X _10497_/Y _10498_/X vssd1 vssd1 vccd1 vccd1 _10971_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 io_wbs_m2s_addr[10] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
X_06730_ _06730_/A _06730_/B _06730_/C vssd1 vssd1 vccd1 vccd1 _06731_/A sky130_fd_sc_hd__nand3_2
XANTENNA__10193__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06661_ _06661_/A _06661_/B vssd1 vssd1 vccd1 vccd1 _06695_/A sky130_fd_sc_hd__nor2_1
X_05612_ _05612_/A _05612_/B vssd1 vssd1 vccd1 vccd1 _05612_/X sky130_fd_sc_hd__and2_1
X_08400_ _08397_/X _10740_/Q _08394_/X _08399_/X vssd1 vssd1 vccd1 vccd1 _10722_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09380_ _09338_/X _10065_/C _10063_/B _10062_/A vssd1 vssd1 vccd1 vccd1 _09431_/A
+ sky130_fd_sc_hd__a31o_2
X_06592_ _06949_/B _06952_/A _06591_/Y vssd1 vssd1 vccd1 vccd1 _06593_/C sky130_fd_sc_hd__a21o_1
X_08331_ _08157_/X _08326_/X _08329_/Y _08330_/X vssd1 vssd1 vccd1 vccd1 _10707_/D
+ sky130_fd_sc_hd__o31a_1
X_05543_ _05454_/A _10543_/Q _05641_/A vssd1 vssd1 vccd1 vccd1 _05543_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09399__B _09399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08262_ _08262_/A vssd1 vssd1 vccd1 vccd1 _10700_/D sky130_fd_sc_hd__clkbuf_1
X_05474_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05474_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07213_ _07186_/A _07125_/A _07222_/B _07211_/A vssd1 vssd1 vccd1 vccd1 _07214_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08193_ _06195_/X _08164_/X _08165_/X _08191_/A _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08193_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08028__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07144_ _07144_/A _07144_/B vssd1 vssd1 vccd1 vccd1 _07148_/A sky130_fd_sc_hd__and2_1
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07075_ _07377_/A _07151_/A _07076_/B _07390_/B vssd1 vssd1 vccd1 vccd1 _07402_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06026_ _10581_/Q _10582_/Q vssd1 vssd1 vccd1 vccd1 _09403_/B sky130_fd_sc_hd__and2b_2
XFILLER_114_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07977_ _07977_/A vssd1 vssd1 vccd1 vccd1 _07977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09716_ _09716_/A _09760_/B vssd1 vssd1 vccd1 vccd1 _09716_/Y sky130_fd_sc_hd__nand2_1
X_06928_ _06928_/A _06928_/B vssd1 vssd1 vccd1 vccd1 _06928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06859_ _06859_/A _06859_/B vssd1 vssd1 vccd1 vccd1 _06860_/B sky130_fd_sc_hd__nor2_1
X_09647_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__xnor2_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08494__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09563_/A _09563_/B _09564_/A vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__a21oi_1
XFILLER_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08529_ _06008_/A _10394_/B _08418_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _08529_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10529__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10422_ input20/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__a21bo_1
XFILLER_137_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08660__C _08989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ _10351_/X _06412_/A _10346_/X _10921_/Q vssd1 vssd1 vccd1 vccd1 _10921_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10284_ _10941_/Q _10957_/Q vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_29_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10174__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07900_ _07900_/A vssd1 vssd1 vccd1 vccd1 _07900_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_97_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08880_ _08814_/A _08891_/A _08878_/X _08879_/Y vssd1 vssd1 vccd1 vccd1 _08881_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07831_ hold11/X _07845_/B vssd1 vssd1 vccd1 vccd1 _07831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07941__A1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09501_ _09501_/A _09501_/B _09501_/C vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__nand3_1
XFILLER_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07762_ _06871_/A _06871_/B _07761_/X vssd1 vssd1 vccd1 vccd1 _07763_/B sky130_fd_sc_hd__o21a_1
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06713_ _06719_/B _06635_/B _06634_/A vssd1 vssd1 vccd1 vccd1 _06714_/B sky130_fd_sc_hd__o21a_1
X_07693_ _07693_/A _07693_/B vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08939__D_N input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ _09432_/A vssd1 vssd1 vccd1 vccd1 _10066_/A sky130_fd_sc_hd__clkbuf_2
X_06644_ _06841_/A _06408_/B _06408_/C vssd1 vssd1 vccd1 vccd1 _06645_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06575_ _10973_/Q _06575_/B vssd1 vssd1 vccd1 vccd1 _06951_/A sky130_fd_sc_hd__nand2_1
X_09363_ _09420_/A _10885_/Q vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__nor2_1
X_08314_ input34/X vssd1 vssd1 vccd1 vccd1 _08314_/Y sky130_fd_sc_hd__inv_2
X_05526_ _10711_/Q vssd1 vssd1 vccd1 vccd1 _06115_/A sky130_fd_sc_hd__buf_2
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _10343_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__and2_2
X_08245_ _06105_/B _08058_/X _08243_/Y _08244_/Y _08062_/X vssd1 vssd1 vccd1 vccd1
+ _08245_/Y sky130_fd_sc_hd__a311oi_1
XFILLER_119_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05457_ _09020_/A _05283_/Y _05286_/B _08994_/A vssd1 vssd1 vccd1 vccd1 _05457_/X
+ sky130_fd_sc_hd__a211o_1
X_08176_ _06187_/X _08164_/X _08165_/X _05692_/A _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08176_/X sky130_fd_sc_hd__o221a_1
XFILLER_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05388_ _05388_/A _05392_/A vssd1 vssd1 vccd1 vccd1 _05389_/B sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_2_3_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07658__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07127_ _07748_/B _07147_/A vssd1 vssd1 vccd1 vccd1 _07133_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07058_ _07197_/B vssd1 vssd1 vccd1 vccd1 _07076_/B sky130_fd_sc_hd__clkbuf_2
X_06009_ _10579_/Q vssd1 vssd1 vccd1 vccd1 _08236_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_30_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07393__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10971_ _10978_/CLK _10971_/D vssd1 vssd1 vccd1 vccd1 _10971_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08893__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clock clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10962_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07999__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06120__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07568__A _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10940_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10405_/X sky130_fd_sc_hd__and2_1
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10336_ _10291_/S _10324_/A _10334_/Y _10335_/Y _10334_/A vssd1 vssd1 vccd1 vccd1
+ _10336_/X sky130_fd_sc_hd__o32a_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10267_ _10266_/X _10259_/X _10257_/B vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__a21o_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08176__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10198_ _10198_/A _10198_/B vssd1 vssd1 vccd1 vccd1 _10198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08100__A1 _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06360_ _06360_/A _09302_/B _06736_/A vssd1 vssd1 vccd1 vccd1 _06360_/X sky130_fd_sc_hd__or3_1
X_05311_ _10674_/Q _10673_/Q _05844_/B vssd1 vssd1 vccd1 vccd1 _05834_/A sky130_fd_sc_hd__or3_2
X_06291_ _10910_/Q vssd1 vssd1 vccd1 vccd1 _06993_/A sky130_fd_sc_hd__clkbuf_4
Xinput30 io_wbs_m2s_data[22] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_4
X_08030_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08030_/X sky130_fd_sc_hd__buf_4
Xinput41 io_wbs_m2s_data[3] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09981_ _09907_/A _09907_/B _09911_/A vssd1 vssd1 vccd1 vccd1 _09982_/B sky130_fd_sc_hd__o21a_1
XFILLER_115_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08932_ _08929_/Y _08930_/X _08931_/X vssd1 vssd1 vccd1 vccd1 _10830_/D sky130_fd_sc_hd__o21a_1
XFILLER_130_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08167__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08863_ _08658_/X _08860_/X _08866_/B _08862_/X vssd1 vssd1 vccd1 vccd1 _08864_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08794_ _06202_/X _08728_/X _08729_/X _10813_/Q vssd1 vssd1 vccd1 vccd1 _08794_/X
+ sky130_fd_sc_hd__a22o_1
X_07814_ hold24/X _07824_/B vssd1 vssd1 vccd1 vccd1 _07814_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07745_ _07745_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07746_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09415_ _09443_/B _09487_/A _09411_/A _09449_/A _10964_/Q vssd1 vssd1 vccd1 vccd1
+ _09454_/A sky130_fd_sc_hd__o2111a_2
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07677_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06627_ _06841_/A _06627_/B vssd1 vssd1 vccd1 vccd1 _06719_/B sky130_fd_sc_hd__nand2_2
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06558_ _10972_/Q _06558_/B _06558_/C vssd1 vssd1 vccd1 vccd1 _06558_/X sky130_fd_sc_hd__and3_1
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _08025_/A _09276_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__mux2_1
X_05509_ _05350_/X _05503_/X _05506_/X _07885_/A vssd1 vssd1 vccd1 vccd1 _10560_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_06489_ _06600_/A _06489_/B vssd1 vssd1 vccd1 vccd1 _06541_/C sky130_fd_sc_hd__nand2_2
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08228_ _08228_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_126_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08159_ _08158_/X _08160_/B _08058_/A vssd1 vssd1 vccd1 vccd1 _08159_/X sky130_fd_sc_hd__a21bo_1
XFILLER_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10121_ _10120_/X _10101_/A _10121_/S vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ _10052_/A _10051_/A vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10280__B1_N _10253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input19_A io_wbs_m2s_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07851__A _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08330__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__B2 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10954_ _10955_/CLK _10954_/D vssd1 vssd1 vccd1 vccd1 _10954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10885_ _10984_/CLK _10885_/D vssd1 vssd1 vccd1 vccd1 _10885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10319_ _10317_/X _10318_/Y _10329_/S vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__mux2_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05860_ _08251_/A _05859_/Y _05857_/B _05858_/Y _10701_/Q vssd1 vssd1 vccd1 vccd1
+ _05860_/X sky130_fd_sc_hd__a32o_1
XFILLER_66_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05791_ _05791_/A _05791_/B vssd1 vssd1 vccd1 vccd1 _05791_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _07638_/B _07639_/A vssd1 vssd1 vccd1 vccd1 _07632_/B sky130_fd_sc_hd__or2b_1
XFILLER_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07461_ _07461_/A _07461_/B _07471_/A vssd1 vssd1 vccd1 vccd1 _07462_/B sky130_fd_sc_hd__nor3_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09200_ _10814_/Q _09168_/X _09079_/X _10727_/Q _09199_/X vssd1 vssd1 vccd1 vccd1
+ _09200_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06412_ _06412_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06732_/A sky130_fd_sc_hd__nor2_1
X_07392_ _07391_/A _07163_/B _07588_/A vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__o21ai_2
XFILLER_22_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09131_ _09153_/A _09131_/B vssd1 vssd1 vccd1 vccd1 _10842_/D sky130_fd_sc_hd__nor2_4
X_06343_ _06343_/A _06371_/C _06352_/C vssd1 vssd1 vccd1 vccd1 _06346_/A sky130_fd_sc_hd__or3_1
X_09062_ _09056_/X _09061_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10838_/D sky130_fd_sc_hd__o21a_2
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06274_ _06305_/A _06274_/B vssd1 vssd1 vccd1 vccd1 _06371_/A sky130_fd_sc_hd__xor2_4
XFILLER_128_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _08013_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09964_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__or2_1
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08915_ _08921_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _08915_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09895_ _09820_/B _09822_/B _09820_/A vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__o21bai_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _08844_/A _08844_/B _08845_/Y _08814_/A vssd1 vssd1 vccd1 vccd1 _08846_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08778_/C sky130_fd_sc_hd__nand2_1
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05989_ input51/X vssd1 vssd1 vccd1 vccd1 _08462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08312__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _07728_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07730_/A sky130_fd_sc_hd__nand2_1
XFILLER_41_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07659_ _07659_/A _07659_/B vssd1 vssd1 vccd1 vccd1 _07688_/B sky130_fd_sc_hd__xor2_2
XFILLER_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10670_ _10673_/CLK _10670_/D vssd1 vssd1 vccd1 vccd1 _10670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09329_ _09329_/A _09329_/B vssd1 vssd1 vccd1 vccd1 _09400_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10537__A _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clock _10857_/CLK vssd1 vssd1 vccd1 vccd1 _10841_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10186__A1 _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10104_ _10104_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__xnor2_4
XFILLER_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10035_ _10035_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_36_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10700_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08551__A1 _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10937_ _10955_/CLK _10937_/D vssd1 vssd1 vccd1 vccd1 _10937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10868_ _10889_/CLK _10868_/D vssd1 vssd1 vccd1 vccd1 _10868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09301__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10799_ _10803_/CLK _10799_/D vssd1 vssd1 vccd1 vccd1 _10799_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09803__A1 _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10413__A2 _10722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07475__B _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06250__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06961_ _07625_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _06962_/B sky130_fd_sc_hd__and2_1
X_05912_ _10648_/Q _05912_/B vssd1 vssd1 vccd1 vccd1 _05913_/B sky130_fd_sc_hd__xor2_1
X_08700_ _10803_/Q vssd1 vssd1 vccd1 vccd1 _08701_/A sky130_fd_sc_hd__buf_2
X_09680_ _09867_/B _09737_/A vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__nand2_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08631_ _10793_/Q _10792_/Q _08631_/C vssd1 vssd1 vccd1 vccd1 _08638_/C sky130_fd_sc_hd__and3_1
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06892_ _06902_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _06894_/A sky130_fd_sc_hd__xor2_4
X_05843_ _05844_/B _05844_/C _05844_/A vssd1 vssd1 vccd1 vccd1 _05845_/A sky130_fd_sc_hd__o21ai_1
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05774_ _10710_/Q vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__inv_2
X_08562_ _08531_/X _08565_/C _10774_/Q _08531_/A vssd1 vssd1 vccd1 vccd1 _08562_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08493_ _08633_/A vssd1 vssd1 vccd1 vccd1 _10355_/A sky130_fd_sc_hd__buf_2
X_07513_ _07513_/A _07516_/A vssd1 vssd1 vccd1 vccd1 _07514_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07444_ _07717_/A _07444_/B vssd1 vssd1 vccd1 vccd1 _07445_/C sky130_fd_sc_hd__nor2_1
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07375_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10404__A2 _10720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ _09114_/A vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06326_ _10928_/Q _10911_/Q _06805_/A _06805_/B _06293_/A vssd1 vssd1 vccd1 vccd1
+ _06851_/B sky130_fd_sc_hd__a221o_1
XFILLER_136_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06257_ _08557_/A vssd1 vssd1 vccd1 vccd1 _06257_/X sky130_fd_sc_hd__clkbuf_2
X_09045_ _09599_/A vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06188_ _10595_/Q vssd1 vssd1 vccd1 vccd1 _06189_/A sky130_fd_sc_hd__inv_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10168__A1 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09947_ _10129_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _10023_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09878_ _09953_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09882_/A sky130_fd_sc_hd__xor2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08829_ _08841_/A _08841_/B _08827_/X _08828_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08829_/X sky130_fd_sc_hd__o311a_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10798_/CLK _10722_/D vssd1 vssd1 vccd1 vccd1 _10722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06745__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10653_ _10654_/CLK _10653_/D vssd1 vssd1 vccd1 vccd1 _10653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ _10808_/CLK _10584_/D vssd1 vssd1 vccd1 vccd1 _10584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _10017_/A _10017_/B _10016_/Y vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__o21bai_1
XFILLER_64_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05490_ _05490_/A vssd1 vssd1 vccd1 vccd1 _05490_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10177__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07160_ _07280_/A _07159_/X vssd1 vssd1 vccd1 vccd1 _07200_/A sky130_fd_sc_hd__or2b_1
X_06111_ _10707_/Q _08324_/B vssd1 vssd1 vccd1 vccd1 _08332_/B sky130_fd_sc_hd__or2_1
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ _07402_/A _07091_/B _07091_/C vssd1 vssd1 vccd1 vccd1 _07363_/B sky130_fd_sc_hd__or3_1
X_06042_ _10705_/Q _08021_/A _05475_/X _05736_/A vssd1 vssd1 vccd1 vccd1 _06045_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08763__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09801_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__inv_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07993_ _08563_/A vssd1 vssd1 vccd1 vccd1 _07993_/X sky130_fd_sc_hd__clkbuf_2
X_09732_ _09432_/A _09679_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__o21a_1
XFILLER_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06944_ _06944_/A _06944_/B vssd1 vssd1 vccd1 vccd1 _07645_/A sky130_fd_sc_hd__nand2_2
XFILLER_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06875_ _06875_/A _06875_/B vssd1 vssd1 vccd1 vccd1 _06878_/A sky130_fd_sc_hd__xnor2_2
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ _09661_/X _09663_/B vssd1 vssd1 vccd1 vccd1 _09779_/B sky130_fd_sc_hd__and2b_1
X_05826_ _05525_/B _08034_/A _05831_/C vssd1 vssd1 vccd1 vccd1 _05826_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05453__B _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08614_ _10788_/Q vssd1 vssd1 vccd1 vccd1 _08614_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09594_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09595_/B sky130_fd_sc_hd__nand2_1
X_08545_ _08545_/A vssd1 vssd1 vccd1 vccd1 _10769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05757_ _08242_/A _05752_/Y _10559_/Q _08232_/A vssd1 vssd1 vccd1 vccd1 _05765_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05688_ _05570_/X _05571_/X _05686_/X _05687_/X vssd1 vssd1 vccd1 vccd1 _05688_/X
+ sky130_fd_sc_hd__o211a_1
X_08476_ _10779_/Q hold6/A _08476_/S vssd1 vssd1 vccd1 vccd1 _08477_/B sky130_fd_sc_hd__mux2_1
XFILLER_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ _07428_/A _07428_/B _07428_/C vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__a21o_1
XFILLER_10_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07358_ _07070_/A _07398_/B _07562_/A vssd1 vssd1 vccd1 vccd1 _07359_/B sky130_fd_sc_hd__and3b_1
XFILLER_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06309_ _06734_/A _06309_/B vssd1 vssd1 vccd1 vccd1 _06731_/B sky130_fd_sc_hd__nand2_2
X_07289_ _07289_/A _07305_/B _07304_/B vssd1 vssd1 vccd1 vccd1 _07289_/X sky130_fd_sc_hd__or3b_1
XFILLER_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09028_ _09805_/A vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08754__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08939__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10705_ _10705_/CLK _10705_/D vssd1 vssd1 vccd1 vccd1 _10705_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10636_ _10826_/CLK _10636_/D vssd1 vssd1 vccd1 vccd1 _10636_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06048__A2 _08032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ _10865_/CLK _10567_/D vssd1 vssd1 vccd1 vccd1 _10567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10498_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput6 io_wbs_m2s_addr[11] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09170__B2 _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ _06660_/A _06660_/B vssd1 vssd1 vccd1 vccd1 _06661_/B sky130_fd_sc_hd__nor2_1
X_05611_ _10555_/Q _05663_/A _05663_/B _10556_/Q vssd1 vssd1 vccd1 vccd1 _05612_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_52_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06591_ _06591_/A _06591_/B vssd1 vssd1 vccd1 vccd1 _06591_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ input35/X _08248_/X _08088_/X _08324_/A _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08330_/X sky130_fd_sc_hd__o221a_1
X_05542_ _05482_/X _05741_/B _05541_/X vssd1 vssd1 vccd1 vccd1 _05641_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08261_ _08259_/X _08261_/B vssd1 vssd1 vccd1 vccd1 _08262_/A sky130_fd_sc_hd__and2b_1
X_05473_ _05479_/A vssd1 vssd1 vccd1 vccd1 _05517_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07212_ _07415_/A _07244_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07214_/A sky130_fd_sc_hd__or3b_1
X_08192_ _06117_/C _08074_/X _08191_/Y _08044_/A _07988_/A vssd1 vssd1 vccd1 vccd1
+ _08192_/X sky130_fd_sc_hd__a32o_1
XFILLER_118_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ _10985_/Q _07327_/A _07490_/A vssd1 vssd1 vccd1 vccd1 _07144_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__08105__A _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07074_ _07186_/B vssd1 vssd1 vccd1 vccd1 _07390_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06025_ _08096_/A vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__buf_4
XFILLER_105_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07976_ _07976_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07976_/X sky130_fd_sc_hd__or2_1
XFILLER_101_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _09780_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__xnor2_1
X_06927_ _06938_/A _06938_/B _06926_/X vssd1 vssd1 vccd1 vccd1 _06937_/B sky130_fd_sc_hd__a21o_1
XFILLER_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09161__B2 _10723_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09646_ _09695_/B _09646_/B vssd1 vssd1 vccd1 vccd1 _09647_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06858_ _07780_/C _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06859_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05809_ _05787_/B _05791_/Y _05792_/Y _05802_/Y _05808_/X vssd1 vssd1 vccd1 vccd1
+ _05809_/X sky130_fd_sc_hd__a311o_1
XFILLER_55_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ _06741_/A _06834_/B _06788_/X vssd1 vssd1 vccd1 vccd1 _06832_/A sky130_fd_sc_hd__o21ai_2
X_09577_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09623_/A sky130_fd_sc_hd__nor2_1
XFILLER_42_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08528_ _10765_/Q _08419_/B _08527_/X vssd1 vssd1 vccd1 vccd1 _10765_/D sky130_fd_sc_hd__a21o_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08121__C1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08459_ _10774_/Q _10737_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ _10944_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__and2_1
XFILLER_137_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08015__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10352_ _10351_/X _06387_/B _10346_/X _10920_/Q vssd1 vssd1 vccd1 vccd1 _10920_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10981__CLK _10981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10283_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10283_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10534__A1 _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input49_A io_wbs_m2s_stb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10619_ _10652_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _10619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08966__A1 _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10525__A1 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07830_ _10577_/Q vssd1 vssd1 vccd1 vccd1 _07845_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07761_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07761_/X sky130_fd_sc_hd__or2_1
XANTENNA__10704__CLK _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06712_ _06718_/B _06712_/B vssd1 vssd1 vccd1 vccd1 _06722_/A sky130_fd_sc_hd__and2_1
X_09500_ _09542_/B _09499_/B _09499_/C vssd1 vssd1 vccd1 vccd1 _09501_/C sky130_fd_sc_hd__a21o_1
XFILLER_37_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07692_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09575_/C sky130_fd_sc_hd__and2b_1
XFILLER_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _09431_/A _09431_/B vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__xor2_4
X_06643_ _06643_/A _06643_/B vssd1 vssd1 vccd1 vccd1 _06702_/B sky130_fd_sc_hd__xor2_4
X_06574_ _06585_/A _06585_/B _06573_/C vssd1 vssd1 vccd1 vccd1 _06578_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _09420_/A _10885_/Q vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__nand2_1
X_05525_ _05525_/A _05525_/B vssd1 vssd1 vccd1 vccd1 _10572_/D sky130_fd_sc_hd__nor2_1
X_08313_ _09154_/A vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__buf_6
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07457__A1 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09293_ _10829_/Q _09274_/X _09275_/X _09292_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09294_/B sky130_fd_sc_hd__a32o_1
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08244_ _08244_/A _08306_/B vssd1 vssd1 vccd1 vccd1 _08244_/Y sky130_fd_sc_hd__nor2_1
X_05456_ _10618_/Q vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__06843__A _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08175_ _08175_/A vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__buf_2
X_05387_ _10622_/Q vssd1 vssd1 vccd1 vccd1 _05462_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07126_ _10985_/Q _07474_/B vssd1 vssd1 vccd1 vccd1 _07147_/A sky130_fd_sc_hd__nand2_1
XFILLER_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07057_ _07166_/B vssd1 vssd1 vccd1 vccd1 _07197_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06008_ _06008_/A vssd1 vssd1 vccd1 vccd1 _06008_/X sky130_fd_sc_hd__buf_4
XANTENNA__10516__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05943__A1 _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07959_ _08443_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07960_/A sky130_fd_sc_hd__or2_1
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10970_ _10970_/CLK _10970_/D vssd1 vssd1 vccd1 vccd1 _10970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09629_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__and2_1
XFILLER_71_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08645__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06120__A1 _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07849__A _07849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10275__A _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10404_ _10389_/X _10720_/Q _10402_/X _10403_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10939_/D sky130_fd_sc_hd__o221a_1
XFILLER_109_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10335_ _10324_/A _10327_/A _10279_/S vssd1 vssd1 vccd1 vccd1 _10335_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10266_ _10938_/Q _10954_/Q vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2b_1
XANTENNA__10507__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10197_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_120_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09125__B2 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09304__A _09304_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05310_ _05336_/A vssd1 vssd1 vccd1 vccd1 _05844_/B sky130_fd_sc_hd__clkbuf_2
X_06290_ _10927_/Q _10910_/Q vssd1 vssd1 vccd1 vccd1 _06293_/A sky130_fd_sc_hd__and2_1
XFILLER_30_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput31 io_wbs_m2s_data[23] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_4
Xinput20 io_wbs_m2s_data[13] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
XFILLER_128_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05279__A _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput42 io_wbs_m2s_data[4] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_4
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09980_ _09980_/A _09980_/B vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__xnor2_1
XFILLER_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ input40/X _08819_/X _08820_/X _10830_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08931_/X sky130_fd_sc_hd__o221a_1
X_08862_ input30/X _08830_/A _08831_/A _10821_/Q vssd1 vssd1 vccd1 vccd1 _08862_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07813_ _06255_/X _10616_/Q _06257_/X _07812_/Y vssd1 vssd1 vccd1 vccd1 _10616_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08793_ _08803_/C _08790_/X _08791_/X _08792_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08793_/X sky130_fd_sc_hd__o311a_1
XFILLER_53_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07744_ _07744_/A _07744_/B vssd1 vssd1 vccd1 vccd1 _07745_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07675_ _07675_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _07677_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09414_ _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09487_/A sky130_fd_sc_hd__and2_1
X_06626_ _06626_/A vssd1 vssd1 vccd1 vccd1 _06841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09345_ _09344_/B _10892_/Q vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__and2b_1
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06557_ _06561_/B _07675_/B vssd1 vssd1 vccd1 vccd1 _06587_/C sky130_fd_sc_hd__and2_1
XFILLER_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09276_ _08324_/A _07914_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09276_/X sky130_fd_sc_hd__mux2_1
X_05508_ _05353_/X _05503_/X _05506_/X _07882_/A vssd1 vssd1 vccd1 vccd1 _10559_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06488_ _06567_/A vssd1 vssd1 vccd1 vccd1 _06600_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08227_ _08092_/X _08232_/B _08226_/X _08096_/X vssd1 vssd1 vccd1 vccd1 _08227_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05439_ _10642_/Q vssd1 vssd1 vccd1 vccd1 _07911_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06292__B _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08158_ _08160_/A vssd1 vssd1 vccd1 vccd1 _08158_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08089_ _10528_/A _08086_/X _08088_/X _05733_/X _08166_/A vssd1 vssd1 vccd1 vccd1
+ _08090_/B sky130_fd_sc_hd__o221a_1
XFILLER_107_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07109_ _07215_/B vssd1 vssd1 vccd1 vccd1 _07125_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_121_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10120_ _10102_/A _10102_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _10120_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10051_ _10051_/A _10052_/A vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__or2b_1
XFILLER_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10953_ _10955_/CLK _10953_/D vssd1 vssd1 vccd1 vccd1 _10953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10884_ _10984_/CLK _10884_/D vssd1 vssd1 vccd1 vccd1 _10884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09291__A0 _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10318_ _10307_/A _10309_/Y _10307_/B vssd1 vssd1 vccd1 vccd1 _10318_/Y sky130_fd_sc_hd__o21bai_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ _10249_/A vssd1 vssd1 vccd1 vccd1 _10249_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05790_ _05765_/C _05789_/X _05765_/B vssd1 vssd1 vccd1 vccd1 _05791_/B sky130_fd_sc_hd__a21bo_1
XFILLER_66_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07460_ _07460_/A _07460_/B vssd1 vssd1 vccd1 vccd1 _07746_/A sky130_fd_sc_hd__xnor2_2
X_07391_ _07391_/A _07391_/B vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__nand2_1
X_06411_ _06717_/A _06411_/B vssd1 vssd1 vccd1 vccd1 _06431_/A sky130_fd_sc_hd__or2_1
XFILLER_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08085__B2 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09130_ _09112_/X _09122_/Y _09129_/X vssd1 vssd1 vccd1 vccd1 _09131_/B sky130_fd_sc_hd__a21oi_1
X_06342_ _06342_/A _06342_/B vssd1 vssd1 vccd1 vccd1 _06352_/C sky130_fd_sc_hd__xor2_2
XANTENNA_clkbuf_leaf_73_clock_A _10981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _10487_/A _10474_/B _10495_/B _10508_/A _09060_/X vssd1 vssd1 vccd1 vccd1
+ _09061_/X sky130_fd_sc_hd__a221o_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08012_ input29/X _08002_/X _08011_/X _08006_/X vssd1 vssd1 vccd1 vccd1 _10669_/D
+ sky130_fd_sc_hd__o211a_1
X_06273_ _06263_/Y _06270_/A _06276_/A _06272_/Y vssd1 vssd1 vccd1 vccd1 _06274_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08793__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_2_clock _10981_/CLK vssd1 vssd1 vccd1 vccd1 _10956_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08914_ _08927_/A _08921_/B vssd1 vssd1 vccd1 vccd1 _08915_/B sky130_fd_sc_hd__or2_1
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09894_ _09894_/A _09893_/Y vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__or2b_1
XFILLER_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08845_ _08845_/A vssd1 vssd1 vccd1 vccd1 _08845_/Y sky130_fd_sc_hd__inv_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08776_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08778_/B sky130_fd_sc_hd__or2_1
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05472__A _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05988_ _09078_/A _05975_/X _05987_/Y _05977_/X vssd1 vssd1 vccd1 vccd1 _10575_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_85_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07727_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08848__B1 _08674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07658_ _07670_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07659_/B sky130_fd_sc_hd__nand2_1
XFILLER_41_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07589_ _07589_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07593_/A sky130_fd_sc_hd__xnor2_2
X_06609_ _06758_/A vssd1 vssd1 vccd1 vccd1 _06856_/A sky130_fd_sc_hd__clkbuf_2
X_09328_ _09312_/X _09325_/Y _09402_/B _09327_/X vssd1 vssd1 vccd1 vccd1 _10867_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08076__B2 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06087__B1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _09259_/A _09259_/B vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__and2_1
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ _10029_/A _10029_/B _10022_/A vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__09328__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input31_A io_wbs_m2s_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10034_ _09955_/A _09955_/B _09960_/A vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10936_ _10955_/CLK _10936_/D vssd1 vssd1 vccd1 vccd1 _10936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _10889_/CLK _10867_/D vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dfxtp_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10798_/CLK _10798_/D vssd1 vssd1 vccd1 vccd1 _10798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09029__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06960_ _07630_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__and2b_1
X_05911_ _05911_/A _05911_/B vssd1 vssd1 vccd1 vccd1 _05911_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_67_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06891_ _06891_/A _06891_/B vssd1 vssd1 vccd1 vccd1 _06930_/A sky130_fd_sc_hd__xnor2_4
X_05842_ _10673_/Q vssd1 vssd1 vccd1 vccd1 _05844_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08630_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _10792_/D sky130_fd_sc_hd__nor2_1
XFILLER_94_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05773_ _10709_/Q vssd1 vssd1 vccd1 vccd1 _06113_/A sky130_fd_sc_hd__clkinv_2
X_08561_ _10773_/Q _08559_/B _08560_/X _08030_/X vssd1 vssd1 vccd1 vccd1 _10773_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08492_ input51/X _09403_/B vssd1 vssd1 vccd1 vccd1 _08633_/A sky130_fd_sc_hd__nor2_1
X_07512_ _07522_/B _07512_/B vssd1 vssd1 vccd1 vccd1 _07657_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07443_ _07715_/C _07726_/B _07732_/B _07442_/X vssd1 vssd1 vccd1 vccd1 _07444_/B
+ sky130_fd_sc_hd__a22oi_1
X_09113_ _09113_/A vssd1 vssd1 vccd1 vccd1 _09113_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ _07374_/A _07374_/B vssd1 vssd1 vccd1 vccd1 _07456_/A sky130_fd_sc_hd__xor2_1
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06325_ _06734_/B _06318_/X _06735_/A _06322_/X _06324_/X vssd1 vssd1 vccd1 vccd1
+ _06805_/B sky130_fd_sc_hd__o311ai_4
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06256_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08557_/A sky130_fd_sc_hd__buf_2
X_09044_ _09489_/A vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10373__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06187_ input18/X vssd1 vssd1 vccd1 vccd1 _06187_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08230__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__B2 _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09946_ _10031_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07682__A _07682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _09943_/B _09877_/B vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__or2_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08828_ _08841_/B _08827_/X _08841_/A vssd1 vssd1 vccd1 vccd1 _08828_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08759_ _08759_/A _08759_/B vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__and2_1
XFILLER_61_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10737_/CLK _10721_/D vssd1 vssd1 vccd1 vccd1 _10721_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08018__A _08018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09246__A0 _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10652_ _10652_/CLK _10652_/D vssd1 vssd1 vccd1 vccd1 _10652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _10652_/CLK _10583_/D vssd1 vssd1 vccd1 vccd1 _10583_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10283__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_clock_A _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07592__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10017_ _10017_/A _10017_/B _10016_/Y vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09312__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10919_ _10980_/CLK _10919_/D vssd1 vssd1 vccd1 vccd1 _10919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06110_ _10706_/Q _08317_/B vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__or2_1
XANTENNA__07767__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ _07359_/A _07090_/B vssd1 vssd1 vccd1 vccd1 _07091_/C sky130_fd_sc_hd__or2_1
XFILLER_133_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06041_ _08105_/A _06038_/X _06040_/X vssd1 vssd1 vccd1 vccd1 _06071_/A sky130_fd_sc_hd__o21ai_1
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07992_ _10441_/A vssd1 vssd1 vccd1 vccd1 _08563_/A sky130_fd_sc_hd__buf_2
X_09800_ _09867_/B _09937_/A vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08598__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ _09731_/A _09731_/B vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__xnor2_2
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06943_ _06943_/A _06943_/B _06943_/C vssd1 vssd1 vccd1 vccd1 _06944_/B sky130_fd_sc_hd__nand3_1
XFILLER_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06874_ _06874_/A _06874_/B vssd1 vssd1 vccd1 vccd1 _06881_/A sky130_fd_sc_hd__or2_2
X_09662_ _09662_/A _09662_/B _09660_/Y vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__or3b_1
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05825_ _05844_/C vssd1 vssd1 vccd1 vccd1 _05831_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_08613_ _08613_/A vssd1 vssd1 vccd1 vccd1 _10787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09593_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05756_ _05756_/A vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__clkbuf_2
X_08544_ _08580_/B _08544_/B _08544_/C vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__and3_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05687_ _08350_/A _05687_/B vssd1 vssd1 vccd1 vccd1 _05687_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_20_clock _10857_/CLK vssd1 vssd1 vccd1 vccd1 _10839_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10368__A _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ _08475_/A vssd1 vssd1 vccd1 vccd1 _10741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07426_ _07426_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07428_/C sky130_fd_sc_hd__xnor2_1
XFILLER_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07357_ _07377_/A _07390_/B _07357_/C vssd1 vssd1 vccd1 vccd1 _07360_/A sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_35_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10707_/CLK sky130_fd_sc_hd__clkbuf_16
X_06308_ _10923_/Q _10906_/Q vssd1 vssd1 vccd1 vccd1 _06309_/B sky130_fd_sc_hd__or2_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09027_ _09555_/A vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__clkbuf_2
X_07288_ _07302_/A _07344_/A _07279_/B vssd1 vssd1 vccd1 vccd1 _07304_/B sky130_fd_sc_hd__o21ai_1
X_06239_ _06253_/B vssd1 vssd1 vccd1 vccd1 _06249_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_105_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09340__A_N _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08939__C _08939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09929_ _09929_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _10704_/CLK _10704_/D vssd1 vssd1 vccd1 vccd1 _10704_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10635_ _10814_/CLK _10635_/D vssd1 vssd1 vccd1 vccd1 _10635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07587__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10566_ _10865_/CLK _10566_/D vssd1 vssd1 vccd1 vccd1 _10566_/Q sky130_fd_sc_hd__dfxtp_1
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10497_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 io_wbs_m2s_addr[1] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_4
XFILLER_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05610_ _05610_/A _05610_/B vssd1 vssd1 vccd1 vccd1 _05610_/X sky130_fd_sc_hd__and2_1
XFILLER_25_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06590_ _06951_/A _06951_/B vssd1 vssd1 vccd1 vccd1 _06952_/A sky130_fd_sc_hd__nor2_1
X_05541_ _05643_/A _05539_/Y _05540_/X vssd1 vssd1 vccd1 vccd1 _05541_/X sky130_fd_sc_hd__a21o_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08260_ input28/X _08212_/X _08124_/X _05598_/X _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08261_/B sky130_fd_sc_hd__o221a_1
X_05472_ _05490_/A _05472_/B vssd1 vssd1 vccd1 vccd1 _05479_/A sky130_fd_sc_hd__or2_1
XANTENNA__08881__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08191_ _08191_/A _08191_/B vssd1 vssd1 vccd1 vccd1 _08191_/Y sky130_fd_sc_hd__xnor2_1
X_07211_ _07211_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07244_/A sky130_fd_sc_hd__nand2_1
X_07142_ _10986_/Q _07142_/B vssd1 vssd1 vccd1 vccd1 _07490_/A sky130_fd_sc_hd__nand2_2
XANTENNA__08433__A1 _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07073_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07377_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06024_ _06024_/A vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07944__A0 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ _06172_/X _07965_/X _07974_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10656_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09217__A _09228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09714_ _09553_/A _09656_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09715_/B sky130_fd_sc_hd__a21oi_1
X_06926_ _06925_/B _06926_/B vssd1 vssd1 vccd1 vccd1 _06926_/X sky130_fd_sc_hd__and2b_1
XFILLER_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06857_ _07682_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06859_/A sky130_fd_sc_hd__and3_1
X_09645_ _09596_/A _09595_/B _09593_/Y vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05808_ _05785_/B _05807_/Y _05528_/A _05564_/A vssd1 vssd1 vccd1 vccd1 _05808_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_70_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _10506_/A _07784_/B _07773_/B _06900_/A vssd1 vssd1 vccd1 vccd1 _06788_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09576_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__nand2_1
X_05739_ _08132_/A _05739_/B vssd1 vssd1 vccd1 vccd1 _05742_/C sky130_fd_sc_hd__nor2_1
X_08527_ _06124_/A _10394_/B _08418_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _08527_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_70_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06295__B _10905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08458_ _08476_/S vssd1 vssd1 vccd1 vccd1 _08473_/S sky130_fd_sc_hd__buf_2
XFILLER_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07409_ _07540_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07410_/B sky130_fd_sc_hd__xor2_1
XFILLER_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10420_ _10408_/X _10724_/Q _10418_/X _10419_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10943_/D sky130_fd_sc_hd__o221a_1
X_08389_ _08383_/X _10736_/Q _08380_/X _08388_/X vssd1 vssd1 vccd1 vccd1 _10718_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ _10351_/A vssd1 vssd1 vccd1 vccd1 _10351_/X sky130_fd_sc_hd__clkbuf_2
X_10282_ _07013_/A _10253_/A _10281_/Y _08563_/X vssd1 vssd1 vccd1 vccd1 _10907_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09127__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05410__A1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09688__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07870__A _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08360__B1 _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06910__B2 _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06910__A1 _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10618_ _10652_/CLK _10618_/D vssd1 vssd1 vccd1 vccd1 _10618_/Q sky130_fd_sc_hd__dfxtp_1
X_10549_ _10657_/CLK _10549_/D vssd1 vssd1 vccd1 vccd1 _10549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09128__C1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ _06393_/A _06393_/B _07801_/A vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__a21o_1
XFILLER_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06711_ _06711_/A _06711_/B vssd1 vssd1 vccd1 vccd1 _06712_/B sky130_fd_sc_hd__or2_1
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07691_ _09483_/A _09483_/B _07654_/A vssd1 vssd1 vccd1 vccd1 _09532_/B sky130_fd_sc_hd__o21ai_2
X_09430_ _09430_/A _09430_/B vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__xnor2_2
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06901__A1 _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06642_ _06642_/A _06642_/B vssd1 vssd1 vccd1 vccd1 _06885_/A sky130_fd_sc_hd__nor2_2
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06573_ _06585_/A _06585_/B _06573_/C vssd1 vssd1 vccd1 vccd1 _06578_/A sky130_fd_sc_hd__nand3_1
X_09361_ _09361_/A _09361_/B vssd1 vssd1 vccd1 vccd1 _09676_/B sky130_fd_sc_hd__nor2_2
X_08312_ _08157_/X _08307_/X _08309_/Y _08311_/X vssd1 vssd1 vccd1 vccd1 _10705_/D
+ sky130_fd_sc_hd__o31a_1
X_09292_ _08352_/A _09291_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09292_/X sky130_fd_sc_hd__mux2_1
X_05524_ _10647_/Q vssd1 vssd1 vccd1 vccd1 _05525_/A sky130_fd_sc_hd__inv_2
X_08243_ _08243_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _08243_/Y sky130_fd_sc_hd__nand2_1
X_05455_ _10619_/Q vssd1 vssd1 vccd1 vccd1 _05455_/X sky130_fd_sc_hd__clkbuf_2
X_08174_ _06117_/C _08074_/X _08173_/Y _08044_/X _07981_/A vssd1 vssd1 vccd1 vccd1
+ _08174_/X sky130_fd_sc_hd__a32o_1
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05386_ _10623_/Q vssd1 vssd1 vccd1 vccd1 _05462_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07125_ _07125_/A vssd1 vssd1 vccd1 vccd1 _07474_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07056_ _07056_/A _07056_/B vssd1 vssd1 vccd1 vccd1 _07166_/B sky130_fd_sc_hd__xor2_2
XFILLER_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06007_ input27/X vssd1 vssd1 vccd1 vccd1 _06008_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_68_clock_A _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07958_ _10535_/A _08119_/A _07983_/A vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08786__A _08820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ _07889_/A vssd1 vssd1 vccd1 vccd1 _07889_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_56_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06909_ _09302_/B _06367_/A _06368_/B vssd1 vssd1 vccd1 vccd1 _06914_/A sky130_fd_sc_hd__o21a_2
XFILLER_55_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09628_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _09516_/A _09516_/C _09516_/B vssd1 vssd1 vccd1 vccd1 _09560_/B sky130_fd_sc_hd__a21boi_4
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10403_ _06172_/X _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__a21bo_1
XFILLER_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07865__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10334_ _10334_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10334_/Y sky130_fd_sc_hd__nor2_1
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__nor2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10196_ _10196_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__nor2_1
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09291__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09125__A2 _09136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10230__S _10291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10443__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09320__A _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput21 io_wbs_m2s_data[14] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_4
Xinput10 io_wbs_m2s_addr[4] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_4
Xinput32 io_wbs_m2s_data[24] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput43 io_wbs_m2s_data[5] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_4
XANTENNA__09061__A1 _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09061__B2 _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08930_ _08920_/A _08927_/X _08928_/X _08814_/A vssd1 vssd1 vccd1 vccd1 _08930_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_123_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08861_ _08870_/C _08861_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07812_ _06134_/A _06258_/X _07807_/X _07809_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07812_/Y sky130_fd_sc_hd__o221ai_4
X_08792_ _08790_/X _08791_/X _08803_/C vssd1 vssd1 vccd1 vccd1 _08792_/Y sky130_fd_sc_hd__o21ai_1
X_07743_ _07743_/A _07743_/B _07743_/C vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__or3_1
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07674_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05689__A1 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06625_ _06643_/A _06643_/B vssd1 vssd1 vccd1 vccd1 _06641_/B sky130_fd_sc_hd__nor2_1
X_09413_ _09494_/B _09413_/B vssd1 vssd1 vccd1 vccd1 _09429_/A sky130_fd_sc_hd__or2_1
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06854__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ _10892_/Q _09344_/B vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__and2b_1
X_06556_ _10971_/Q _06575_/B vssd1 vssd1 vccd1 vccd1 _07675_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05507_ _05358_/X _05503_/X _05506_/X _07878_/A vssd1 vssd1 vccd1 vccd1 _10558_/D
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09230__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09275_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06487_ _10973_/Q vssd1 vssd1 vccd1 vccd1 _06567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08226_ _08216_/X _08208_/A _08207_/B _06061_/A vssd1 vssd1 vccd1 vccd1 _08226_/X
+ sky130_fd_sc_hd__a31o_1
X_05438_ _07907_/A _05332_/Y _05437_/X vssd1 vssd1 vccd1 vccd1 _05438_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08157_ _08157_/A vssd1 vssd1 vccd1 vccd1 _08157_/X sky130_fd_sc_hd__buf_2
XFILLER_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05369_ _05369_/A _05369_/B vssd1 vssd1 vccd1 vccd1 _05369_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09052__B2 _08701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07108_ _07747_/A _07108_/B vssd1 vssd1 vccd1 vccd1 _07215_/B sky130_fd_sc_hd__xnor2_2
X_08088_ _08355_/B vssd1 vssd1 vccd1 vccd1 _08088_/X sky130_fd_sc_hd__buf_2
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07039_ _07416_/A _07472_/A _07039_/C vssd1 vssd1 vccd1 vccd1 _07424_/A sky130_fd_sc_hd__and3_1
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _10050_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09405__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10952_ _10956_/CLK _10952_/D vssd1 vssd1 vccd1 vccd1 _10952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _10920_/CLK _10883_/D vssd1 vssd1 vccd1 vccd1 _10883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10425__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09286__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10317_ _10307_/A _10310_/X _10307_/B vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__o21ba_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10248_ _10224_/A _10935_/Q _10233_/X _10235_/B _10247_/Y vssd1 vssd1 vccd1 vccd1
+ _10249_/A sky130_fd_sc_hd__o311a_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10179_ _06997_/B _10174_/X _10177_/X _10890_/Q vssd1 vssd1 vccd1 vccd1 _10890_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_93_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10113__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06410_ _06626_/A _06428_/B _06872_/A vssd1 vssd1 vccd1 vccd1 _06411_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07390_ _07592_/A _07390_/B vssd1 vssd1 vccd1 vccd1 _07391_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08085__A2 _08043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10416__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06341_ _06371_/B vssd1 vssd1 vccd1 vccd1 _06343_/A sky130_fd_sc_hd__inv_2
X_09060_ _10935_/Q _10394_/C _10430_/B _10951_/Q vssd1 vssd1 vccd1 vccd1 _09060_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06272_ _10918_/Q _10901_/Q vssd1 vssd1 vccd1 vccd1 _06272_/Y sky130_fd_sc_hd__nor2_1
X_08011_ _08268_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08011_/X sky130_fd_sc_hd__or2_1
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _09962_/A _09962_/B vssd1 vssd1 vccd1 vccd1 _09964_/B sky130_fd_sc_hd__xnor2_1
XFILLER_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08913_ _10828_/Q _08919_/B vssd1 vssd1 vccd1 vccd1 _08921_/B sky130_fd_sc_hd__and2_1
XFILLER_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09893_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09893_/Y sky130_fd_sc_hd__nand2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08844_ _08844_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__or2_1
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05987_ _05992_/B _05986_/X _05993_/S vssd1 vssd1 vccd1 vccd1 _05987_/Y sky130_fd_sc_hd__a21oi_1
X_08775_ _08804_/A _08804_/B _08804_/C _08806_/A vssd1 vssd1 vccd1 vccd1 _08777_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07726_ _07726_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07734_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08848__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__B _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07657_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__nor2_1
XFILLER_41_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06608_ _06607_/A _06607_/B _06607_/C vssd1 vssd1 vccd1 vccd1 _06614_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07588_ _07588_/A _07588_/B vssd1 vssd1 vccd1 vccd1 _07589_/B sky130_fd_sc_hd__xor2_2
X_09327_ hold24/A _10283_/A vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__and2_1
X_06539_ _06532_/A _06532_/B _06538_/X vssd1 vssd1 vccd1 vccd1 _06542_/A sky130_fd_sc_hd__o21ba_1
XFILLER_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06087__B2 _05721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06087__A1 _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09258_ _08876_/A _09243_/X _09244_/X _09257_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09259_/B sky130_fd_sc_hd__a32o_1
X_08209_ _08209_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08209_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09189_ _05460_/B _09136_/A _09148_/X _05877_/X _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09189_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08023__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10102_ _10102_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10104_/A sky130_fd_sc_hd__xnor2_4
XFILLER_76_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10033_ _10105_/B _10033_/B vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__xnor2_2
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input24_A io_wbs_m2s_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10935_ _10935_/CLK _10935_/D vssd1 vssd1 vccd1 vccd1 _10935_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__05522__B1 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10866_ _10920_/CLK _10866_/D vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10797_ _10797_/CLK _10797_/D vssd1 vssd1 vccd1 vccd1 _10797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06250__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08527__B1 _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05910_ _06065_/A _05910_/B vssd1 vssd1 vccd1 vccd1 _05911_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06890_ _06932_/B _06890_/B vssd1 vssd1 vccd1 vccd1 _06935_/A sky130_fd_sc_hd__xnor2_4
X_05841_ _05337_/B _08018_/A _05844_/C vssd1 vssd1 vccd1 vccd1 _05841_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05772_ _10565_/Q vssd1 vssd1 vccd1 vccd1 _05772_/Y sky130_fd_sc_hd__inv_2
X_08560_ _08531_/X _08559_/X _10773_/Q _08531_/A vssd1 vssd1 vccd1 vccd1 _08560_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08491_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08491_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07511_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07512_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07442_ _07573_/A vssd1 vssd1 vccd1 vccd1 _07442_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07373_ _07373_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07374_/B sky130_fd_sc_hd__nand2_1
X_09112_ _09112_/A vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06324_ _06323_/Y _06317_/A _06313_/A vssd1 vssd1 vccd1 vccd1 _06324_/X sky130_fd_sc_hd__o21a_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06255_ _07848_/A vssd1 vssd1 vccd1 vccd1 _06255_/X sky130_fd_sc_hd__clkbuf_2
X_09043_ _10966_/Q vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06186_ _06182_/X _06183_/X _06185_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10594_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08124__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06241__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09945_ _09945_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__xnor2_1
XFILLER_131_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08518__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09876_ _09876_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09877_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07682__B _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08827_ _10816_/Q _08815_/A _08928_/B vssd1 vssd1 vccd1 vccd1 _08827_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08758_ _08758_/A _08758_/B vssd1 vssd1 vccd1 vccd1 _08804_/A sky130_fd_sc_hd__and2_1
XFILLER_57_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _10802_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07709_ _10045_/A _10045_/B _07708_/X vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__o21ai_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _10737_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _10720_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08018__B _08021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10651_/CLK _10651_/D vssd1 vssd1 vccd1 vccd1 _10651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10582_ _10803_/CLK _10582_/D vssd1 vssd1 vccd1 vccd1 _10582_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08034__A _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07873__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06232__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07980__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10016_ _09945_/A _09945_/B _09929_/B vssd1 vssd1 vccd1 vccd1 _10016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_1_clock _10981_/CLK vssd1 vssd1 vccd1 vccd1 _10924_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10918_ _10980_/CLK _10918_/D vssd1 vssd1 vccd1 vccd1 _10918_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08209__A _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849_ _10852_/CLK _10849_/D vssd1 vssd1 vccd1 vccd1 _10849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05568__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06040_ _05749_/A _08289_/A _07976_/A _05711_/Y vssd1 vssd1 vccd1 vccd1 _06040_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07991_ _07991_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _07991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07783__A _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09730_ _09793_/B _09730_/B vssd1 vssd1 vccd1 vccd1 _09731_/B sky130_fd_sc_hd__xnor2_1
X_06942_ _06942_/A _06942_/B vssd1 vssd1 vccd1 vccd1 _07641_/A sky130_fd_sc_hd__or2_2
XFILLER_95_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06873_ _06383_/C _06873_/B vssd1 vssd1 vccd1 vccd1 _06874_/B sky130_fd_sc_hd__and2b_1
X_09661_ _09662_/A _09662_/B _09660_/Y vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__o21ba_1
X_05824_ _05854_/B vssd1 vssd1 vccd1 vccd1 _05844_/C sky130_fd_sc_hd__clkbuf_2
X_08612_ _10355_/A _08612_/B _08612_/C vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__and3_1
X_09592_ _09640_/A _09592_/B vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__or2_1
X_05755_ _10698_/Q vssd1 vssd1 vccd1 vccd1 _05756_/A sky130_fd_sc_hd__inv_2
X_08543_ _10769_/Q _08543_/B vssd1 vssd1 vccd1 vccd1 _08544_/C sky130_fd_sc_hd__nand2_1
XFILLER_82_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05686_ _05574_/X _05576_/X _05571_/X _05570_/X _05685_/X vssd1 vssd1 vccd1 vccd1
+ _05686_/X sky130_fd_sc_hd__a221o_1
X_08474_ _08477_/A _08474_/B vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__or2_1
XFILLER_50_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07425_ _07425_/A _07425_/B vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__or2_1
X_07356_ _07560_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07406_/A sky130_fd_sc_hd__nand2_2
X_06307_ _10923_/Q _10906_/Q vssd1 vssd1 vccd1 vccd1 _06734_/A sky130_fd_sc_hd__nand2_2
XFILLER_40_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07287_ _07287_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _07305_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__05478__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06238_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06238_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09026_ _10965_/Q vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06169_ _10591_/Q vssd1 vssd1 vccd1 vccd1 _06170_/A sky130_fd_sc_hd__inv_2
XFILLER_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09928_ _10056_/C _10069_/B vssd1 vssd1 vccd1 vccd1 _09929_/B sky130_fd_sc_hd__or2_1
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09859_ _09859_/A vssd1 vssd1 vccd1 vccd1 _09859_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05941__A _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10705_/CLK _10703_/D vssd1 vssd1 vccd1 vccd1 _10703_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10634_ _10814_/CLK _10634_/D vssd1 vssd1 vccd1 vccd1 _10634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05388__A _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10565_ _10646_/CLK _10565_/D vssd1 vssd1 vccd1 vccd1 _10565_/Q sky130_fd_sc_hd__dfxtp_2
X_10496_ _10497_/B vssd1 vssd1 vccd1 vccd1 _10496_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07650__B1 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06205__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput8 io_wbs_m2s_addr[2] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_4
XANTENNA__07108__A _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05851__A _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05540_ _10574_/Q _10542_/Q vssd1 vssd1 vccd1 vccd1 _05540_/X sky130_fd_sc_hd__xor2_1
XFILLER_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05471_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05471_/X sky130_fd_sc_hd__clkbuf_4
X_08190_ _08092_/X _08196_/B _08189_/X _08096_/X vssd1 vssd1 vccd1 vccd1 _08190_/X
+ sky130_fd_sc_hd__a31o_1
X_07210_ _07210_/A _07260_/A vssd1 vssd1 vccd1 vccd1 _07275_/A sky130_fd_sc_hd__xnor2_1
XFILLER_20_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07141_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07296_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08433__A2 _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07072_ _10986_/Q vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__clkbuf_2
X_06023_ _10583_/Q _06023_/B vssd1 vssd1 vccd1 vccd1 _06024_/A sky130_fd_sc_hd__nand2_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07944__A1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07974_ _07974_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07974_/X sky130_fd_sc_hd__or2_1
XFILLER_101_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09713_ _09713_/A _09713_/B vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07018__A _07229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06925_ _06926_/B _06925_/B vssd1 vssd1 vccd1 vccd1 _06938_/B sky130_fd_sc_hd__xnor2_2
X_09644_ _09644_/A _09769_/C vssd1 vssd1 vccd1 vccd1 _09695_/B sky130_fd_sc_hd__xor2_1
X_06856_ _06856_/A _07766_/B _06856_/C vssd1 vssd1 vccd1 vccd1 _06857_/C sky130_fd_sc_hd__and3_1
XFILLER_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05807_ _05807_/A _05807_/B vssd1 vssd1 vccd1 vccd1 _05807_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06857__A _07682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ _10506_/A _07773_/B vssd1 vssd1 vccd1 vccd1 _06834_/B sky130_fd_sc_hd__nand2_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09575_ _09575_/A _09575_/B _09575_/C vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__or3_1
XFILLER_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05738_ _08130_/A vssd1 vssd1 vccd1 vccd1 _08132_/A sky130_fd_sc_hd__clkbuf_2
X_08526_ _08526_/A vssd1 vssd1 vccd1 vccd1 _10764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05669_ _10695_/Q _05612_/X _05610_/X _08224_/B _05668_/X vssd1 vssd1 vccd1 vccd1
+ _05669_/X sky130_fd_sc_hd__a221o_1
X_08457_ _08457_/A vssd1 vssd1 vccd1 vccd1 _10736_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_64_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07408_ _07543_/A _07361_/B _07407_/X vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__a21bo_1
X_08388_ _08395_/A _10752_/Q vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__or2_1
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07339_ _07528_/B _07339_/B vssd1 vssd1 vccd1 vccd1 _07526_/A sky130_fd_sc_hd__nand2_1
X_10350_ _09312_/X _06371_/A _10346_/X _10919_/Q vssd1 vssd1 vccd1 vccd1 _10919_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09009_ _10948_/Q _10432_/C _09008_/X _10932_/Q vssd1 vssd1 vccd1 vccd1 _09009_/X
+ sky130_fd_sc_hd__a22o_1
X_10281_ _10276_/Y _10279_/X _10280_/Y vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_105_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09408__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09385__B1 _09417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05410__A2 _10616_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09688__A1 _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08663__A2 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10617_ _10652_/CLK _10617_/D vssd1 vssd1 vccd1 vccd1 _10617_/Q sky130_fd_sc_hd__dfxtp_1
X_10548_ _10657_/CLK _10548_/D vssd1 vssd1 vccd1 vccd1 _10548_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06007__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05846__A _10671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10479_ _06124_/X _10475_/X _10478_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10963_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06710_ _06711_/A _06711_/B vssd1 vssd1 vccd1 vccd1 _06718_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_34_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10710_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07690_ _07687_/A _07687_/B _07688_/B _09442_/A vssd1 vssd1 vccd1 vccd1 _09483_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06641_ _06641_/A _06641_/B _06641_/C vssd1 vssd1 vccd1 vccd1 _06642_/B sky130_fd_sc_hd__nor3_1
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06572_ _06571_/A _06571_/C _06571_/B vssd1 vssd1 vccd1 vccd1 _06594_/B sky130_fd_sc_hd__a21oi_1
XFILLER_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09360_ _10902_/Q _10886_/Q vssd1 vssd1 vccd1 vccd1 _09361_/B sky130_fd_sc_hd__and2b_1
X_08311_ input33/X _08248_/X _08088_/X _08305_/A _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08311_/X sky130_fd_sc_hd__o221a_1
X_05523_ _05318_/X _05517_/X _05471_/X _07925_/A vssd1 vssd1 vccd1 vccd1 _10571_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09291_ _08351_/A _07925_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_49_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10823_/CLK sky130_fd_sc_hd__clkbuf_16
X_08242_ _08242_/A vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05454_ _05454_/A vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__buf_2
X_08173_ _08173_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08173_/Y sky130_fd_sc_hd__xnor2_1
X_05385_ _10655_/Q _05389_/A vssd1 vssd1 vccd1 vccd1 _05385_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_137_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07124_ _07137_/A _07229_/B vssd1 vssd1 vccd1 vccd1 _07748_/B sky130_fd_sc_hd__nand2_2
XFILLER_134_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07055_ _07113_/A _07475_/B _07112_/A vssd1 vssd1 vccd1 vccd1 _07056_/B sky130_fd_sc_hd__o21a_1
X_06006_ _06006_/A vssd1 vssd1 vccd1 vccd1 _10578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__A _09228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ _08445_/A vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07971__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06908_ _06928_/A _06928_/B vssd1 vssd1 vccd1 vccd1 _06937_/A sky130_fd_sc_hd__xor2_4
X_07888_ _07906_/A vssd1 vssd1 vccd1 vccd1 _07888_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06839_ _06839_/A _06839_/B vssd1 vssd1 vccd1 vccd1 _06840_/B sky130_fd_sc_hd__nand2_1
X_09627_ _09682_/A _09627_/B vssd1 vssd1 vccd1 vccd1 _09629_/B sky130_fd_sc_hd__xor2_2
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09558_ _09597_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__xnor2_2
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08509_ _10177_/A vssd1 vssd1 vccd1 vccd1 _08509_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10437__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05459__A2 _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09489_ _09489_/A _09555_/A _09642_/A _09492_/A vssd1 vssd1 vccd1 vccd1 _09618_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _10939_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10402_/X sky130_fd_sc_hd__and2_1
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10333_ _10962_/Q _10946_/Q vssd1 vssd1 vccd1 vccd1 _10333_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10264_ _10955_/Q _10939_/Q vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__and2b_1
XFILLER_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10195_ _10932_/Q _10948_/Q vssd1 vssd1 vccd1 vccd1 _10196_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07881__A _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput11 io_wbs_m2s_addr[5] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_4
Xinput22 io_wbs_m2s_data[15] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_4
Xinput33 io_wbs_m2s_data[25] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_4
Xinput44 io_wbs_m2s_data[6] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10482__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _08870_/C _08861_/B vssd1 vssd1 vccd1 vccd1 _08860_/X sky130_fd_sc_hd__or2_1
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07811_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07811_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_111_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08791_ _08778_/B _08803_/B vssd1 vssd1 vccd1 vccd1 _08791_/X sky130_fd_sc_hd__and2b_1
XFILLER_65_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07742_ _07406_/A _07544_/A _07753_/A vssd1 vssd1 vccd1 vccd1 _07743_/C sky130_fd_sc_hd__a21oi_1
XFILLER_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06200__A _07977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07673_ _07673_/A _07673_/B vssd1 vssd1 vccd1 vccd1 _07674_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06624_ _06624_/A _06650_/A _06624_/C vssd1 vssd1 vccd1 vccd1 _06643_/B sky130_fd_sc_hd__and3_2
XFILLER_16_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09412_ _09489_/A _09536_/B _09579_/A _10965_/Q vssd1 vssd1 vccd1 vccd1 _09413_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09343_ _09343_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06555_ _06555_/A _06555_/B vssd1 vssd1 vccd1 vccd1 _06585_/A sky130_fd_sc_hd__xnor2_2
X_05506_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05506_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09274_ _09274_/A vssd1 vssd1 vccd1 vccd1 _09274_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06486_ _06486_/A _06486_/B vssd1 vssd1 vccd1 vccd1 _06643_/A sky130_fd_sc_hd__xnor2_4
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08225_ _08233_/B vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__inv_2
X_05437_ _10641_/Q _05332_/Y _05337_/X _05436_/X vssd1 vssd1 vccd1 vccd1 _05437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08156_ _08156_/A vssd1 vssd1 vccd1 vccd1 _10689_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05368_ _10660_/Q _05886_/A _10661_/Q vssd1 vssd1 vccd1 vccd1 _05369_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07966__A _08414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07107_ _10913_/Q _07747_/B vssd1 vssd1 vccd1 vccd1 _07108_/B sky130_fd_sc_hd__nand2_1
X_08087_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__buf_2
X_05299_ _05374_/A vssd1 vssd1 vccd1 vccd1 _05886_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10392__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _07428_/B _07038_/B vssd1 vssd1 vccd1 vccd1 _07051_/A sky130_fd_sc_hd__and2_1
XFILLER_121_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08990_/C sky130_fd_sc_hd__nand2_1
XFILLER_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10951_ _10978_/CLK _10951_/D vssd1 vssd1 vccd1 vccd1 _10951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10882_ _10982_/CLK _10882_/D vssd1 vssd1 vccd1 vccd1 _10882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10316_ _10316_/A _10316_/B vssd1 vssd1 vccd1 vccd1 _10320_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10247_ _10247_/A vssd1 vssd1 vccd1 vccd1 _10247_/Y sky130_fd_sc_hd__inv_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10178_ _07083_/A _10174_/X _10177_/X _10889_/Q vssd1 vssd1 vccd1 vccd1 _10889_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06340_ _06459_/B vssd1 vssd1 vccd1 vccd1 _07682_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06271_ _06275_/A _06275_/B vssd1 vssd1 vccd1 vccd1 _06276_/A sky130_fd_sc_hd__nand2_1
X_08010_ input28/X _08002_/X _08009_/Y _08006_/X vssd1 vssd1 vccd1 vccd1 _10668_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09961_ _09961_/A _09961_/B vssd1 vssd1 vccd1 vccd1 _09962_/B sky130_fd_sc_hd__nor2_1
X_08912_ _10828_/Q _08918_/B vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09892_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__nor2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08843_ _08871_/A _08873_/A vssd1 vssd1 vccd1 vccd1 _08844_/B sky130_fd_sc_hd__nor2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05986_ input44/X input43/X vssd1 vssd1 vccd1 vccd1 _05986_/X sky130_fd_sc_hd__or2_1
X_08774_ _10810_/Q _10809_/Q _10808_/Q _08748_/X _08801_/B vssd1 vssd1 vccd1 vccd1
+ _08806_/A sky130_fd_sc_hd__o41a_1
XFILLER_57_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07725_ _07726_/A _07732_/B _07577_/B _07576_/A vssd1 vssd1 vccd1 vccd1 _07735_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08848__A2 _08672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07656_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__and2_1
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06607_ _06607_/A _06607_/B _06607_/C vssd1 vssd1 vccd1 vccd1 _06614_/A sky130_fd_sc_hd__nand3_1
X_07587_ _07592_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07588_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10407__A2 _10721_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09326_ _09326_/A _09326_/B vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__or2_1
X_06538_ _06533_/A _06538_/B vssd1 vssd1 vccd1 vccd1 _06538_/X sky130_fd_sc_hd__and2b_1
X_09257_ _08298_/A _09256_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09257_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08208_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08208_/Y sky130_fd_sc_hd__nand2_1
X_06469_ _06448_/B _06469_/B vssd1 vssd1 vccd1 vccd1 _06470_/B sky130_fd_sc_hd__and2b_1
XFILLER_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ _09113_/A _09187_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08139_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__and2_1
XFILLER_122_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10101_ _10101_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__and2_1
XFILLER_130_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10032_ _10030_/X _09952_/B _10031_/X vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__o21a_1
XFILLER_49_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input17_A io_wbs_m2s_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _10955_/CLK _10934_/D vssd1 vssd1 vccd1 vccd1 _10934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10865_ _10865_/CLK _10865_/D vssd1 vssd1 vccd1 vccd1 _10865_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10796_ _10978_/CLK _10796_/D vssd1 vssd1 vccd1 vccd1 _10796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09297__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07027__A1 _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06015__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05840_ _08298_/A vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__inv_2
XFILLER_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05771_ _05771_/A vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _07510_/A _07510_/B vssd1 vssd1 vccd1 vccd1 _07633_/A sky130_fd_sc_hd__nor2_1
X_08490_ _10181_/A vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__buf_2
XFILLER_35_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07441_ _07574_/A vssd1 vssd1 vccd1 vccd1 _07715_/C sky130_fd_sc_hd__clkbuf_4
X_07372_ _07373_/A _07374_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07454_/B sky130_fd_sc_hd__and3_1
X_09111_ _09111_/A vssd1 vssd1 vccd1 vccd1 _10841_/D sky130_fd_sc_hd__clkbuf_1
X_06323_ _10926_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _06323_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06254_ input40/X _06145_/B _06253_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10615_/D
+ sky130_fd_sc_hd__o211a_1
X_09042_ _07732_/A _08965_/Y _09036_/X _09038_/X _09041_/X vssd1 vssd1 vccd1 vccd1
+ _09042_/X sky130_fd_sc_hd__a221o_1
X_06185_ hold8/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09944_ _10012_/A _09944_/B vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__or2_1
XANTENNA__09236__A _09236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A io_wbs_m2s_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _09876_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09943_/B sky130_fd_sc_hd__and2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09191__B2 _10726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08826_ _08817_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__and2b_1
XFILLER_58_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08757_ _10809_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08758_/B sky130_fd_sc_hd__or2_1
X_05969_ _08414_/A _08939_/C vssd1 vssd1 vccd1 vccd1 _06126_/D sky130_fd_sc_hd__or2_1
XFILLER_72_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _08688_/A vssd1 vssd1 vccd1 vccd1 _08688_/X sky130_fd_sc_hd__buf_2
X_07708_ _07708_/A _07605_/B vssd1 vssd1 vccd1 vccd1 _07708_/X sky130_fd_sc_hd__or2b_1
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07639_ _07639_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _07693_/A sky130_fd_sc_hd__xor2_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10650_ _10651_/CLK _10650_/D vssd1 vssd1 vccd1 vccd1 _10650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09309_ _09313_/B _09310_/C _09396_/A vssd1 vssd1 vccd1 vccd1 _09309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10581_ _10803_/CLK _10581_/D vssd1 vssd1 vccd1 vccd1 _10581_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08315__A _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08034__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09182__B2 _10725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10017_/B sky130_fd_sc_hd__and2_1
XFILLER_49_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10917_ _10980_/CLK _10917_/D vssd1 vssd1 vccd1 vccd1 _10917_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08209__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10848_ _10848_/CLK _10848_/D vssd1 vssd1 vccd1 vccd1 _10848_/Q sky130_fd_sc_hd__dfxtp_1
X_10779_ _10781_/CLK _10779_/D vssd1 vssd1 vccd1 vccd1 _10779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08996__A1 _05721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07990_ _08015_/A vssd1 vssd1 vccd1 vccd1 _08021_/B sky130_fd_sc_hd__buf_2
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06941_ _06941_/A _06941_/B _06944_/A vssd1 vssd1 vccd1 vccd1 _06942_/B sky130_fd_sc_hd__and3_1
X_09660_ _09713_/A _09713_/B vssd1 vssd1 vccd1 vccd1 _09660_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08611_ _10787_/Q _08611_/B vssd1 vssd1 vccd1 vccd1 _08612_/C sky130_fd_sc_hd__nand2_1
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06872_ _06872_/A _06872_/B vssd1 vssd1 vccd1 vccd1 _06873_/B sky130_fd_sc_hd__nand2_1
X_05823_ _05823_/A vssd1 vssd1 vccd1 vccd1 _05854_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09591_ _09590_/B _09591_/B vssd1 vssd1 vccd1 vccd1 _09592_/B sky130_fd_sc_hd__and2b_1
X_05754_ _05751_/Y _10561_/Q _05752_/Y _08242_/A vssd1 vssd1 vccd1 vccd1 _05765_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10857__CLK _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ _10769_/Q _08543_/B vssd1 vssd1 vccd1 vccd1 _08544_/B sky130_fd_sc_hd__or2_1
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08473_ _10778_/Q _10741_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08474_/B sky130_fd_sc_hd__mux2_1
XFILLER_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05685_ _05679_/X _05683_/X _05576_/X _08339_/B _05684_/X vssd1 vssd1 vccd1 vccd1
+ _05685_/X sky130_fd_sc_hd__o221a_1
XANTENNA__08119__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08684__B1 _08674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07424_ _07424_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _07425_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07355_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07366_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05759__A _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07286_ _07286_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _07287_/B sky130_fd_sc_hd__nor2_1
X_06306_ _06263_/Y _06270_/A _06276_/A _06305_/X _06272_/Y vssd1 vssd1 vccd1 vccd1
+ _06730_/C sky130_fd_sc_hd__a311o_1
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06237_ input32/X _06225_/X _06236_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10608_/D
+ sky130_fd_sc_hd__o211a_1
X_09025_ _10714_/Q _08990_/C _09024_/X vssd1 vssd1 vccd1 vccd1 _09025_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07974__A _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06168_ _10537_/A vssd1 vssd1 vccd1 vccd1 _06168_/X sky130_fd_sc_hd__buf_6
XFILLER_2_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06099_ _10689_/Q _08150_/B vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__or2_1
XFILLER_132_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09927_ _10056_/C _10069_/B vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__nand2_1
XFILLER_49_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_60_clock_A _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09858_ _10076_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__nand2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _08804_/Y _08806_/Y _08801_/X _08802_/Y vssd1 vssd1 vccd1 vccd1 _08817_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09789_ _09848_/B _09789_/B vssd1 vssd1 vccd1 vccd1 _09827_/B sky130_fd_sc_hd__and2_2
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08029__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10702_ _10702_/CLK _10702_/D vssd1 vssd1 vccd1 vccd1 _10702_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__B1 _08674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _10811_/CLK _10633_/D vssd1 vssd1 vccd1 vccd1 _10633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10564_ _10646_/CLK _10564_/D vssd1 vssd1 vccd1 vccd1 _10564_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10495_ _10495_/A _10495_/B vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__nand2_2
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 io_wbs_m2s_addr[3] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_49_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09323__B _09323_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05470_ _05470_/A _05470_/B vssd1 vssd1 vccd1 vccd1 _05513_/A sky130_fd_sc_hd__nor2_4
XANTENNA__06141__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06963__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10485__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A1 _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ _07151_/A _07474_/B _07147_/B _07139_/X vssd1 vssd1 vccd1 vccd1 _07295_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_118_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07071_ _07357_/C _07283_/B vssd1 vssd1 vccd1 vccd1 _07284_/A sky130_fd_sc_hd__or2_1
XFILLER_114_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06022_ _08837_/A vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07973_ _08027_/B vssd1 vssd1 vccd1 vccd1 _07988_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09712_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__or2_1
XFILLER_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06924_ _06914_/A _06914_/B _06923_/X vssd1 vssd1 vccd1 vccd1 _06925_/B sky130_fd_sc_hd__a21oi_2
XFILLER_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09643_ _09764_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09769_/C sky130_fd_sc_hd__nand2_1
X_06855_ _06855_/A _06855_/B vssd1 vssd1 vccd1 vccd1 _06857_/B sky130_fd_sc_hd__xnor2_1
X_05806_ _05768_/X _05805_/X _05785_/A vssd1 vssd1 vccd1 vccd1 _05807_/B sky130_fd_sc_hd__o21ai_1
XFILLER_83_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09574_ _09570_/A _09574_/B vssd1 vssd1 vccd1 vccd1 _09631_/B sky130_fd_sc_hd__and2b_1
XFILLER_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08525_ _10763_/Q _10529_/A vssd1 vssd1 vccd1 vccd1 _08526_/A sky130_fd_sc_hd__and2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06786_ _06786_/A vssd1 vssd1 vccd1 vccd1 _07773_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08121__A2 _08061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05737_ _08082_/B _05737_/B vssd1 vssd1 vccd1 vccd1 _05742_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05668_ _05877_/A _05615_/Y _05612_/X _10695_/Q _05667_/X vssd1 vssd1 vccd1 vccd1
+ _05668_/X sky130_fd_sc_hd__o221a_1
X_08456_ _08460_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__or2_1
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08387_ _08383_/X _10735_/Q _08380_/X _08386_/X vssd1 vssd1 vccd1 vccd1 _10717_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07407_ _07407_/A _07360_/A vssd1 vssd1 vccd1 vccd1 _07407_/X sky130_fd_sc_hd__or2b_1
XFILLER_137_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05599_ _10561_/Q _05602_/A vssd1 vssd1 vccd1 vccd1 _05599_/X sky130_fd_sc_hd__xor2_1
X_07338_ _07338_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07339_/B sky130_fd_sc_hd__or2_1
XFILLER_137_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07269_ _07269_/A _07269_/B _07514_/A vssd1 vssd1 vccd1 vccd1 _07270_/B sky130_fd_sc_hd__and3_1
XFILLER_105_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _09008_/A vssd1 vssd1 vccd1 vccd1 _09008_/X sky130_fd_sc_hd__clkbuf_2
X_10280_ _10276_/Y _10279_/X _10253_/A vssd1 vssd1 vccd1 vccd1 _10280_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_132_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_0_clock _10981_/CLK vssd1 vssd1 vccd1 vccd1 _10930_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__05946__B2 _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09137__B2 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08345__C1 _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05952__A _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10616_ _10803_/CLK _10616_/D vssd1 vssd1 vccd1 vccd1 _10616_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10547_ _10654_/CLK _10547_/D vssd1 vssd1 vccd1 vccd1 _10547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10478_ _10478_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10478_/X sky130_fd_sc_hd__or2_1
XFILLER_108_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06023__A _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09128__A1 _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07780__C _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06640_ _06641_/A _06641_/B _06641_/C vssd1 vssd1 vccd1 vccd1 _06642_/A sky130_fd_sc_hd__o21a_1
XFILLER_37_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06571_ _06571_/A _06571_/B _06571_/C vssd1 vssd1 vccd1 vccd1 _06594_/A sky130_fd_sc_hd__and3_1
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09290_ _09290_/A vssd1 vssd1 vccd1 vccd1 _10863_/D sky130_fd_sc_hd__clkbuf_1
X_05522_ _05324_/X _05517_/X _05471_/X _07922_/A vssd1 vssd1 vccd1 vccd1 _10570_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_08310_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08310_/X sky130_fd_sc_hd__buf_2
XFILLER_33_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _08241_/A vssd1 vssd1 vccd1 vccd1 _10698_/D sky130_fd_sc_hd__clkbuf_1
X_05453_ _05453_/A _09107_/A vssd1 vssd1 vccd1 vccd1 _05453_/X sky130_fd_sc_hd__or2_1
XFILLER_60_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08172_ _08092_/X _08181_/B _08171_/X _08096_/X vssd1 vssd1 vccd1 vccd1 _08172_/X
+ sky130_fd_sc_hd__a31o_1
X_05384_ _10624_/Q vssd1 vssd1 vccd1 vccd1 _05461_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07123_ _07144_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07134_/A sky130_fd_sc_hd__xnor2_2
XFILLER_134_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07054_ _07151_/A vssd1 vssd1 vccd1 vccd1 _07560_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06005_ _08483_/A _06005_/B vssd1 vssd1 vccd1 vccd1 _06006_/A sky130_fd_sc_hd__and2_1
XFILLER_88_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07956_ _07956_/A vssd1 vssd1 vccd1 vccd1 _10653_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07971__B _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09244__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06907_ _06904_/X _06922_/B _06906_/X vssd1 vssd1 vccd1 vccd1 _06928_/B sky130_fd_sc_hd__a21oi_4
X_07887_ _07898_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _10635_/D sky130_fd_sc_hd__nor2_1
XFILLER_56_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09626_ _09626_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09627_/B sky130_fd_sc_hd__nand2_1
X_06838_ _06839_/A _06839_/B vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__or2_1
XFILLER_55_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06769_ _06769_/A vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09898__B _09898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09557_ _09652_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__or2_1
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08508_ _10790_/Q _08506_/X _08502_/X _10753_/Q vssd1 vssd1 vccd1 vccd1 _10753_/D
+ sky130_fd_sc_hd__a22o_1
X_09488_ _09488_/A vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08439_ _08443_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08440_/A sky130_fd_sc_hd__or2_1
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10401_ _10389_/X _10719_/Q _10398_/X _10400_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10938_/D sky130_fd_sc_hd__o221a_1
X_10332_ _10962_/Q _10946_/Q vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__or2_1
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _10939_/Q _10955_/Q vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__and2b_1
XFILLER_3_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A io_wbs_m2s_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _10948_/Q _10932_/Q vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__and2b_1
XFILLER_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09154__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06018__A _06023_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 io_wbs_m2s_addr[6] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput45 io_wbs_m2s_data[7] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_4
Xinput34 io_wbs_m2s_data[26] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_4
Xinput23 io_wbs_m2s_data[16] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_6
XFILLER_116_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07810_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07874_/A sky130_fd_sc_hd__clkbuf_4
X_08790_ _10812_/Q _08771_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08790_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07741_ _07741_/A _07741_/B vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07672_ _07673_/A _07673_/B vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__or2_1
XFILLER_37_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09411_ _09411_/A vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06623_ _06541_/C _06542_/A _06528_/Y vssd1 vssd1 vccd1 vccd1 _06624_/C sky130_fd_sc_hd__a21o_1
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09342_ _07028_/A _10893_/Q vssd1 vssd1 vccd1 vccd1 _09343_/B sky130_fd_sc_hd__and2b_1
X_06554_ _10972_/Q _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06555_/B sky130_fd_sc_hd__and3_1
X_05505_ _05360_/X _05503_/X _05495_/X _07875_/A vssd1 vssd1 vccd1 vccd1 _10557_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ _09273_/A vssd1 vssd1 vccd1 vccd1 _10860_/D sky130_fd_sc_hd__clkbuf_1
X_06485_ _06486_/A _06486_/B vssd1 vssd1 vccd1 vccd1 _06641_/A sky130_fd_sc_hd__and2_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08224_ _08224_/A _08224_/B _08224_/C vssd1 vssd1 vccd1 vccd1 _08233_/B sky130_fd_sc_hd__and3_1
X_05436_ _07900_/A _05340_/X _05337_/B _10640_/Q _05435_/X vssd1 vssd1 vccd1 vccd1
+ _05436_/X sky130_fd_sc_hd__a221o_1
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08156_/A sky130_fd_sc_hd__and2_1
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05367_ _10629_/Q vssd1 vssd1 vccd1 vccd1 _05460_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__07966__B _08939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09239__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07106_ _07384_/A _07137_/C vssd1 vssd1 vccd1 vccd1 _07144_/A sky130_fd_sc_hd__or2_2
X_08086_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08086_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__08260__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05298_ _10659_/Q _05373_/B vssd1 vssd1 vccd1 vccd1 _05374_/A sky130_fd_sc_hd__or2_1
XFILLER_122_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07037_ _07555_/B _07037_/B vssd1 vssd1 vccd1 vccd1 _07038_/B sky130_fd_sc_hd__nand2_1
XFILLER_114_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08012__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08988_ _09079_/A vssd1 vssd1 vccd1 vccd1 _08988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07939_ _07939_/A vssd1 vssd1 vccd1 vccd1 _10648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10950_ _10956_/CLK _10950_/D vssd1 vssd1 vccd1 vccd1 _10950_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09512__A1 _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__B2 _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10881_ _10958_/CLK _10881_/D vssd1 vssd1 vccd1 vccd1 _10881_/Q sky130_fd_sc_hd__dfxtp_1
X_09609_ _09867_/A _09610_/C _09717_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09611_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__09276__A0 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08318__A _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10845_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08053__A _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10315_ _10960_/Q _10944_/Q vssd1 vssd1 vccd1 vccd1 _10316_/B sky130_fd_sc_hd__and2b_1
XFILLER_106_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07892__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10246_ _10246_/A _10246_/B _10246_/C vssd1 vssd1 vccd1 vccd1 _10247_/A sky130_fd_sc_hd__and3_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_48_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10847_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10177_ _10177_/A vssd1 vssd1 vccd1 vccd1 _10177_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_94_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08711__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09019__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06270_ _06270_/A _06270_/B vssd1 vssd1 vccd1 vccd1 _06275_/B sky130_fd_sc_hd__and2_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10493__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09960_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09962_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08911_ _08904_/B _08907_/B _08904_/A vssd1 vssd1 vccd1 vccd1 _08921_/A sky130_fd_sc_hd__o21bai_1
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09891_ _09961_/B _09891_/B vssd1 vssd1 vccd1 vccd1 _09893_/B sky130_fd_sc_hd__or2_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08842_ _10818_/Q _10817_/Q _10816_/Q _08815_/A _08840_/B vssd1 vssd1 vccd1 vccd1
+ _08873_/A sky130_fd_sc_hd__o41a_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05985_ input44/X input43/X vssd1 vssd1 vccd1 vccd1 _05992_/B sky130_fd_sc_hd__nand2_1
X_08773_ _08773_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07724_ _07724_/A _07724_/B vssd1 vssd1 vccd1 vccd1 _07740_/A sky130_fd_sc_hd__or2_1
XFILLER_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07655_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07657_/B sky130_fd_sc_hd__and2_1
XFILLER_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06606_ _06680_/A _06680_/B vssd1 vssd1 vccd1 vccd1 _06681_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07586_ _07586_/A _07586_/B vssd1 vssd1 vccd1 vccd1 _07751_/A sky130_fd_sc_hd__xnor2_4
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ _09326_/A _09326_/B vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06537_ _06621_/A _06663_/A _06536_/A vssd1 vssd1 vccd1 vccd1 _06544_/B sky130_fd_sc_hd__a21oi_1
X_09256_ _08297_/A _07903_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09256_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07977__A _07977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06468_ _06468_/A _06468_/B vssd1 vssd1 vccd1 vccd1 _06474_/A sky130_fd_sc_hd__nor2_1
X_08207_ _08208_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08207_/Y sky130_fd_sc_hd__nor2_1
X_05419_ _10625_/Q _05380_/Y _05383_/X _05461_/D _05418_/X vssd1 vssd1 vccd1 vccd1
+ _05419_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05497__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ _09114_/A _09186_/X _10500_/B vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06399_ _10975_/Q vssd1 vssd1 vccd1 vccd1 _06441_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08138_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08148_/B sky130_fd_sc_hd__nor2_1
XFILLER_107_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08069_ _06008_/A _08047_/X _08052_/X _08059_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08069_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10100_ _10100_/A _10100_/B _10100_/C vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__nand3_1
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10031_ _10031_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__or2_1
XFILLER_130_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06121__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05960__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10933_ _10946_/CLK _10933_/D vssd1 vssd1 vccd1 vccd1 _10933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10864_ _10865_/CLK _10864_/D vssd1 vssd1 vccd1 vccd1 _10864_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10728__D _10728_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10795_ _10797_/CLK _10795_/D vssd1 vssd1 vccd1 vccd1 _10795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_55_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output78_A _10836_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10229_ _10202_/X _10203_/X _10226_/X _10228_/Y vssd1 vssd1 vccd1 vccd1 _10246_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_67_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05770_ _05767_/Y _10568_/Q _05769_/Y _08317_/A vssd1 vssd1 vccd1 vccd1 _05770_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07440_ _07573_/A _07574_/A _07726_/B _07732_/B vssd1 vssd1 vccd1 vccd1 _07717_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_35_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07371_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07373_/B sky130_fd_sc_hd__or2_1
X_09110_ _09228_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__and2_1
X_06322_ _06734_/A _06320_/Y _06321_/A _06318_/X vssd1 vssd1 vccd1 vccd1 _06322_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_136_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _10577_/Q _08972_/X _08974_/A _09040_/X vssd1 vssd1 vccd1 vccd1 _09041_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07928__A2_N _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06253_ hold17/A _06253_/B vssd1 vssd1 vccd1 vccd1 _06253_/X sky130_fd_sc_hd__or2_1
XFILLER_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06206__A input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06184_ _10594_/Q vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__inv_2
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09943_ _09943_/A _09943_/B _09943_/C vssd1 vssd1 vccd1 vccd1 _09944_/B sky130_fd_sc_hd__nor3_1
XFILLER_131_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09874_ _09943_/A _09874_/B vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__nor2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08825_ _08825_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08841_/A sky130_fd_sc_hd__and2_1
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08756_ _10809_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08758_/A sky130_fd_sc_hd__nand2_1
X_05968_ input14/X input49/X input1/X vssd1 vssd1 vccd1 vccd1 _08939_/C sky130_fd_sc_hd__nand3b_4
XFILLER_26_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05899_ _05388_/A _05904_/A _05295_/A vssd1 vssd1 vccd1 vccd1 _05900_/B sky130_fd_sc_hd__a21o_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _08808_/A vssd1 vssd1 vccd1 vccd1 _08688_/A sky130_fd_sc_hd__buf_2
XFILLER_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07707_ _09969_/A _09969_/B _07706_/X vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__a21oi_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _07715_/D _07638_/B vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07569_ _10912_/Q vssd1 vssd1 vccd1 vccd1 _09379_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09308_ _09449_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09396_/A sky130_fd_sc_hd__nand2_2
X_10580_ _10839_/CLK _10583_/Q vssd1 vssd1 vccd1 vccd1 _10580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09239_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05955__A _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10017_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10916_ _10980_/CLK _10916_/D vssd1 vssd1 vccd1 vccd1 _10916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ _10847_/CLK _10847_/D vssd1 vssd1 vccd1 vccd1 _10847_/Q sky130_fd_sc_hd__dfxtp_1
X_10778_ _10836_/CLK _10778_/D vssd1 vssd1 vccd1 vccd1 _10778_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08506__A _08514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ _06940_/A _06940_/B vssd1 vssd1 vccd1 vccd1 _07636_/A sky130_fd_sc_hd__xnor2_4
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06871_ _06871_/A _06871_/B vssd1 vssd1 vccd1 vccd1 _07799_/A sky130_fd_sc_hd__xnor2_4
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05822_ _05886_/B vssd1 vssd1 vccd1 vccd1 _05823_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08610_ _10786_/Q _08498_/X _08600_/A _08597_/B _10787_/Q vssd1 vssd1 vccd1 vccd1
+ _08612_/B sky130_fd_sc_hd__a41o_1
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09590_ _09591_/B _09590_/B vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__and2b_1
X_05753_ _08251_/B vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__clkbuf_2
X_08541_ _08541_/A vssd1 vssd1 vccd1 vccd1 _10768_/D sky130_fd_sc_hd__clkbuf_1
X_05684_ _08327_/A _05684_/B vssd1 vssd1 vccd1 vccd1 _05684_/X sky130_fd_sc_hd__or2_1
XANTENNA__08684__A1 _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08472_ _08472_/A vssd1 vssd1 vccd1 vccd1 _10740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09881__B1 _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07423_ _07424_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__and2_1
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07354_ _07461_/B _07471_/A _07461_/A vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__o21a_1
X_06305_ _06305_/A _06374_/B _06305_/C vssd1 vssd1 vccd1 vccd1 _06305_/X sky130_fd_sc_hd__or3_1
X_07285_ _07285_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07286_/B sky130_fd_sc_hd__and2_1
XFILLER_136_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06236_ _10608_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06236_/X sky130_fd_sc_hd__or2_1
X_09024_ _10198_/A _08418_/B _09168_/A _10801_/Q _08999_/X vssd1 vssd1 vccd1 vccd1
+ _09024_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07947__A0 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06167_ input45/X vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__buf_4
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06098_ _10688_/Q _10687_/Q _08132_/B vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__or3_1
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09926_ _10068_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07990__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09857_ _09930_/B _09919_/B _09930_/C _09716_/A vssd1 vssd1 vccd1 vccd1 _09858_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08808_ _08808_/A vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09788_ _09787_/A _09787_/B _09787_/C vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__o21ai_1
X_08739_ _08688_/X _08736_/X _08738_/X vssd1 vssd1 vccd1 vccd1 _10806_/D sky130_fd_sc_hd__o21a_1
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10701_ _10702_/CLK _10701_/D vssd1 vssd1 vccd1 vccd1 _10701_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10632_ _10811_/CLK _10632_/D vssd1 vssd1 vccd1 vccd1 _10632_/Q sky130_fd_sc_hd__dfxtp_1
X_10563_ _10673_/CLK _10563_/D vssd1 vssd1 vccd1 vccd1 _10563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10494_ _06168_/X _10489_/B _10493_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10970_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08061__A _08061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10473__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__A1 _07393_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07070_ _07070_/A _07070_/B vssd1 vssd1 vccd1 vccd1 _07283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06021_ _08201_/A vssd1 vssd1 vccd1 vccd1 _08837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ _07995_/A vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__buf_2
X_09711_ _09711_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06923_ _06913_/A _06923_/B vssd1 vssd1 vccd1 vccd1 _06923_/X sky130_fd_sc_hd__and2b_1
XFILLER_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06854_ _07675_/A _07780_/B vssd1 vssd1 vccd1 vccd1 _06855_/B sky130_fd_sc_hd__or2_1
X_09642_ _09642_/A vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05805_ _05783_/X _05804_/X _05770_/X vssd1 vssd1 vccd1 vccd1 _05805_/X sky130_fd_sc_hd__o21ba_1
X_09573_ _09567_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__and2b_1
X_06785_ _06785_/A vssd1 vssd1 vccd1 vccd1 _10506_/A sky130_fd_sc_hd__buf_2
X_05736_ _05736_/A _10541_/Q vssd1 vssd1 vccd1 vccd1 _05742_/A sky130_fd_sc_hd__nor2_1
X_08524_ _08524_/A vssd1 vssd1 vccd1 vccd1 _10763_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09530__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05667_ _05662_/X _05665_/X _05666_/X vssd1 vssd1 vccd1 vccd1 _05667_/X sky130_fd_sc_hd__a21o_1
X_08455_ _10773_/Q _10736_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08456_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10464__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05598_ _08251_/A vssd1 vssd1 vccd1 vccd1 _05598_/X sky130_fd_sc_hd__clkbuf_2
X_08386_ _08395_/A hold26/X vssd1 vssd1 vccd1 vccd1 _08386_/X sky130_fd_sc_hd__or2_1
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07406_ _07406_/A vssd1 vssd1 vccd1 vccd1 _07543_/A sky130_fd_sc_hd__inv_2
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07337_ _07522_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07525_/B sky130_fd_sc_hd__nand2_1
XFILLER_109_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07330_/A sky130_fd_sc_hd__xnor2_1
XFILLER_136_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06219_ input24/X _06207_/X _06218_/X _06200_/X vssd1 vssd1 vccd1 vccd1 _10601_/D
+ sky130_fd_sc_hd__o211a_1
X_09007_ _09124_/C _09098_/B vssd1 vssd1 vccd1 vccd1 _10432_/C sky130_fd_sc_hd__nor2_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07199_ _07277_/A _07277_/B vssd1 vssd1 vccd1 vccd1 _07301_/A sky130_fd_sc_hd__or2b_1
XFILLER_105_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08345__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09909_ _09910_/A _10049_/C vssd1 vssd1 vccd1 vccd1 _09911_/A sky130_fd_sc_hd__or2_1
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10455__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10615_ _10669_/CLK _10615_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09073__B2 _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__A1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10546_ _10654_/CLK _10546_/D vssd1 vssd1 vccd1 vccd1 _10546_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_4_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_10477_ _10493_/B vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_6_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08033__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06023__B _06023_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10260__S _10291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06570_ _06570_/A _06570_/B vssd1 vssd1 vccd1 vccd1 _06599_/A sky130_fd_sc_hd__xnor2_1
X_05521_ _05326_/X _05517_/X _05471_/X _07919_/A vssd1 vssd1 vccd1 vccd1 _10569_/D
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07847__C1 hold4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _08238_/X _08240_/B vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__and2b_1
X_05452_ _05452_/A vssd1 vssd1 vccd1 vccd1 _09107_/A sky130_fd_sc_hd__buf_2
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08171_ _08158_/X _08150_/A _08148_/B _05692_/A vssd1 vssd1 vccd1 vccd1 _08171_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_118_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05383_ _05383_/A _05383_/B vssd1 vssd1 vccd1 vccd1 _05383_/X sky130_fd_sc_hd__and2_1
X_07122_ _07135_/A _07136_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07123_/B sky130_fd_sc_hd__o21bai_4
XFILLER_133_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07053_ _10985_/Q vssd1 vssd1 vccd1 vccd1 _07151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06004_ input38/X _10578_/Q _06120_/S vssd1 vssd1 vccd1 vccd1 _06005_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07955_ _07955_/A _07955_/B vssd1 vssd1 vccd1 vccd1 _07956_/A sky130_fd_sc_hd__or2_1
XFILLER_102_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06906_ _06921_/A _06921_/B vssd1 vssd1 vccd1 vccd1 _06906_/X sky130_fd_sc_hd__and2_1
X_07886_ _10603_/Q _07870_/X _07874_/X _07885_/Y vssd1 vssd1 vccd1 vccd1 _07887_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_56_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09625_ _09625_/A _09625_/B _09566_/A vssd1 vssd1 vccd1 vccd1 _09682_/B sky130_fd_sc_hd__or3b_1
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06837_ _06828_/A _06828_/B _06836_/Y _06796_/B _06796_/A vssd1 vssd1 vccd1 vccd1
+ _06839_/B sky130_fd_sc_hd__o32a_1
XFILLER_15_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06768_ _06774_/B vssd1 vssd1 vccd1 vccd1 _06842_/A sky130_fd_sc_hd__clkbuf_2
X_09556_ _09554_/C _09600_/A vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__and2b_1
X_05719_ _05719_/A vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08507_ _10789_/Q _08506_/X _08502_/X _10752_/Q vssd1 vssd1 vccd1 vccd1 _10752_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10437__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09487_ _09487_/A vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__clkbuf_2
X_06699_ _06916_/A _06912_/B _06698_/X vssd1 vssd1 vccd1 vccd1 _06903_/B sky130_fd_sc_hd__a21o_1
X_08438_ _10768_/Q _10731_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08439_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09055__A1 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10251_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _10537_/A _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10400_/X sky130_fd_sc_hd__a21bo_1
XFILLER_137_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ _09379_/B _10283_/X _10330_/Y _10293_/X vssd1 vssd1 vccd1 vccd1 _10912_/D
+ sky130_fd_sc_hd__a22o_1
X_10262_ _07083_/A _10115_/X _10261_/X _10043_/X vssd1 vssd1 vccd1 vccd1 _10905_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06124__A _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10193_ _09634_/A _10198_/B _10192_/X _07394_/X vssd1 vssd1 vccd1 vccd1 _10898_/D
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06041__A1 _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10428__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 io_wbs_m2s_addr[7] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
Xinput24 io_wbs_m2s_data[17] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_4
Xinput46 io_wbs_m2s_data[8] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput35 io_wbs_m2s_data[27] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_6
XANTENNA__08514__A _08514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10529_ _10529_/A vssd1 vssd1 vccd1 vccd1 _10529_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07740_ _07740_/A _07740_/B vssd1 vssd1 vccd1 vccd1 _07741_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07673_/B sky130_fd_sc_hd__xor2_1
XFILLER_65_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06622_ _06663_/A _06622_/B _06692_/A _06692_/B vssd1 vssd1 vccd1 vccd1 _06650_/A
+ sky130_fd_sc_hd__nand4_1
X_09410_ _10966_/Q _10965_/Q _09443_/B _09411_/A vssd1 vssd1 vccd1 vccd1 _09494_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10419__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _10893_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__and2b_1
X_06553_ _06346_/A _06346_/B _10497_/A vssd1 vssd1 vccd1 vccd1 _06555_/A sky130_fd_sc_hd__a21o_1
X_05504_ _05363_/X _05503_/X _05495_/X _07871_/A vssd1 vssd1 vccd1 vccd1 _10556_/D
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06209__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ _09289_/A _09272_/B vssd1 vssd1 vccd1 vccd1 _09273_/A sky130_fd_sc_hd__and2_1
X_06484_ _06458_/A _06458_/B _06647_/A _06453_/A vssd1 vssd1 vccd1 vccd1 _06486_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08223_ _08157_/X _08219_/X _08221_/Y _08222_/X vssd1 vssd1 vccd1 vccd1 _10696_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05435_ _10639_/Q _05340_/X _05434_/X vssd1 vssd1 vccd1 vccd1 _05435_/X sky130_fd_sc_hd__o21a_1
X_08154_ input47/X _08123_/X _08109_/X _08150_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08155_/B sky130_fd_sc_hd__o221a_1
XANTENNA__08245__C1 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05366_ _08198_/A _05369_/A vssd1 vssd1 vccd1 vccd1 _05366_/Y sky130_fd_sc_hd__xnor2_1
X_08085_ _05279_/A _08043_/A _08080_/Y _06117_/C _08084_/X vssd1 vssd1 vccd1 vccd1
+ _08090_/A sky130_fd_sc_hd__a221o_1
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07105_ _10985_/Q _07394_/A vssd1 vssd1 vccd1 vccd1 _07137_/C sky130_fd_sc_hd__nand2_1
XFILLER_134_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08260__A2 _08212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05297_ _10658_/Q _06039_/A _05383_/A vssd1 vssd1 vccd1 vccd1 _05373_/B sky130_fd_sc_hd__or3_1
X_07036_ _07555_/B _07037_/B vssd1 vssd1 vccd1 vccd1 _07428_/B sky130_fd_sc_hd__or2_1
XFILLER_134_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09255__A _09255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08987_ _09211_/B vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07938_ _09154_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07939_/A sky130_fd_sc_hd__or2_1
XFILLER_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07869_ _10577_/Q _07910_/A vssd1 vssd1 vccd1 vccd1 _07906_/A sky130_fd_sc_hd__and2b_2
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06326__A2 _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10880_ _10958_/CLK _10880_/D vssd1 vssd1 vccd1 vccd1 _10880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ _09608_/A _09608_/B vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__xnor2_2
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09539_ _09596_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__or2_2
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06119__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05958__A _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10314_ _10944_/Q _10960_/Q vssd1 vssd1 vccd1 vccd1 _10316_/A sky130_fd_sc_hd__and2b_1
XFILLER_121_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09200__B2 _10727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10245_ _10245_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10252_/A sky130_fd_sc_hd__nor2_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10176_ _07061_/A _10174_/X _10170_/X _10888_/Q vssd1 vssd1 vccd1 vccd1 _10888_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_51_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09503__A2 _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08509__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10282__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08910_ _09153_/A _08910_/B vssd1 vssd1 vccd1 vccd1 _10827_/D sky130_fd_sc_hd__nor2_1
X_09890_ _09889_/B _09890_/B vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__and2b_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ _08841_/A _08841_/B _08841_/C vssd1 vssd1 vccd1 vccd1 _08871_/A sky130_fd_sc_hd__and3_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05984_ _05482_/X _05975_/X _05982_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10574_/D
+ sky130_fd_sc_hd__a211o_1
X_08772_ _10811_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08773_/B sky130_fd_sc_hd__or2_1
XFILLER_85_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07723_ _07555_/B _07556_/A _07418_/Y vssd1 vssd1 vccd1 vccd1 _07724_/B sky130_fd_sc_hd__a21oi_1
XFILLER_81_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07654_ _07654_/A _07654_/B vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06605_ _06607_/C _06605_/B vssd1 vssd1 vccd1 vccd1 _06680_/B sky130_fd_sc_hd__or2_1
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07585_ _07585_/A _07721_/A vssd1 vssd1 vccd1 vccd1 _07586_/B sky130_fd_sc_hd__xor2_4
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09324_ _09402_/A _09324_/B vssd1 vssd1 vccd1 vccd1 _09326_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06536_ _06536_/A _06536_/B vssd1 vssd1 vccd1 vccd1 _06663_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09255_ _09255_/A vssd1 vssd1 vccd1 vccd1 _10857_/D sky130_fd_sc_hd__clkbuf_1
X_06467_ _06456_/A _06460_/B _06917_/A vssd1 vssd1 vccd1 vccd1 _06468_/B sky130_fd_sc_hd__a21boi_1
X_08206_ _08206_/A vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__clkbuf_2
X_05418_ _10624_/Q _05383_/X _05385_/Y _05462_/A _05417_/X vssd1 vssd1 vccd1 vccd1
+ _05418_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09186_ _10945_/Q _09143_/Y _09185_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09186_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06398_ _06456_/A vssd1 vssd1 vccd1 vccd1 _06626_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10834__D _10834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ _08150_/B _08136_/Y _08062_/A vssd1 vssd1 vccd1 vccd1 _08137_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05349_ _10635_/Q vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08068_ _08075_/B _08072_/B _08067_/X _06033_/X vssd1 vssd1 vccd1 vccd1 _08068_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07993__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07019_ _07472_/A _07434_/A _07416_/A vssd1 vssd1 vccd1 vccd1 _07035_/A sky130_fd_sc_hd__and3b_1
XFILLER_103_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10030_ _10031_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10030_/X sky130_fd_sc_hd__and2_1
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10932_ _10935_/CLK _10932_/D vssd1 vssd1 vccd1 vccd1 _10932_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10863_ _10865_/CLK _10863_/D vssd1 vssd1 vccd1 vccd1 _10863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10794_ _10797_/CLK _10794_/D vssd1 vssd1 vccd1 vccd1 _10794_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06235__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06015__C input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10228_ _10228_/A vssd1 vssd1 vccd1 vccd1 _10228_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__xnor2_4
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08696__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07370_ _07412_/C _07370_/B vssd1 vssd1 vccd1 vccd1 _07374_/A sky130_fd_sc_hd__nor2_1
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06982__A _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06321_ _06321_/A _06320_/Y vssd1 vssd1 vccd1 vccd1 _06735_/A sky130_fd_sc_hd__or2b_2
X_09040_ _05279_/A _08995_/X _09039_/X _08981_/A vssd1 vssd1 vccd1 vccd1 _09040_/X
+ sky130_fd_sc_hd__a211o_1
X_06252_ input39/X _06145_/B _06251_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10614_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06183_ _06204_/B vssd1 vssd1 vccd1 vccd1 _06183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _09943_/A _09943_/B _09943_/C vssd1 vssd1 vccd1 vccd1 _10012_/A sky130_fd_sc_hd__o21a_1
XFILLER_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09873_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09874_/B sky130_fd_sc_hd__and2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08824_ _10817_/Q _08856_/B vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__or2_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _08688_/X _08753_/Y _08754_/X vssd1 vssd1 vccd1 vccd1 _10808_/D sky130_fd_sc_hd__o21a_1
XFILLER_73_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05967_ input15/X input6/X input5/X vssd1 vssd1 vccd1 vccd1 _08414_/A sky130_fd_sc_hd__or3_4
X_07706_ _07610_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _07706_/X sky130_fd_sc_hd__and2b_1
X_05898_ _06038_/A _05906_/A vssd1 vssd1 vccd1 vccd1 _05904_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_32_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10694_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _08686_/A _08819_/A vssd1 vssd1 vccd1 vccd1 _08808_/A sky130_fd_sc_hd__nand2_2
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07637_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07988__A _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ _07726_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_47_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10851_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06519_ _06519_/A _06519_/B vssd1 vssd1 vccd1 vccd1 _06523_/C sky130_fd_sc_hd__nor2_1
X_09307_ _09387_/A vssd1 vssd1 vccd1 vccd1 _09443_/B sky130_fd_sc_hd__clkbuf_2
X_07499_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07504_/A sky130_fd_sc_hd__xnor2_1
X_09238_ _08268_/A _09237_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09238_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06217__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08612__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ _10081_/B _10013_/B vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__or2_1
XFILLER_48_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input22_A io_wbs_m2s_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08142__A1 _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10915_ _10980_/CLK _10915_/D vssd1 vssd1 vccd1 vccd1 _10915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10846_ _10848_/CLK _10846_/D vssd1 vssd1 vccd1 vccd1 _10846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _10836_/CLK _10777_/D vssd1 vssd1 vccd1 vccd1 _10777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09337__B _09337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06870_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _06871_/B sky130_fd_sc_hd__xnor2_2
X_05821_ _05906_/A vssd1 vssd1 vccd1 vccd1 _05886_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05752_ _10560_/Q vssd1 vssd1 vccd1 vccd1 _05752_/Y sky130_fd_sc_hd__inv_2
X_08540_ _08543_/B _08580_/B _08540_/C vssd1 vssd1 vccd1 vccd1 _08541_/A sky130_fd_sc_hd__and3b_1
XFILLER_94_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05683_ _08317_/A _05583_/Y _05684_/B _08327_/A vssd1 vssd1 vccd1 vccd1 _05683_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08133__B2 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08471_ _08477_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _08472_/A sky130_fd_sc_hd__or2_1
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08684__A2 _08672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07422_ _07421_/Y _07043_/A _07417_/A _07044_/A vssd1 vssd1 vccd1 vccd1 _07424_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08416__B _08989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07353_ _07369_/B _07353_/B vssd1 vssd1 vccd1 vccd1 _07461_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06304_ _06304_/A _06304_/B vssd1 vssd1 vccd1 vccd1 _06374_/B sky130_fd_sc_hd__nand2_2
X_07284_ _07284_/A _07284_/B vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__and2_1
X_06235_ input31/X _06225_/X _06233_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10607_/D
+ sky130_fd_sc_hd__o211a_1
X_09023_ _10578_/Q _08972_/X _08974_/X _09022_/X vssd1 vssd1 vccd1 vccd1 _09023_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07947__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06166_ _06163_/X _06158_/X _06165_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10590_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06097_ _10686_/Q _08117_/B vssd1 vssd1 vccd1 vccd1 _08132_/B sky130_fd_sc_hd__or2_2
XFILLER_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09925_ _09925_/A _09925_/B vssd1 vssd1 vccd1 vccd1 _10141_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09856_ _10484_/A _09930_/C _09856_/C vssd1 vssd1 vccd1 vccd1 _10076_/A sky130_fd_sc_hd__nand3_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09263__A _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08807_ _08801_/X _08802_/Y _08804_/Y _08806_/Y vssd1 vssd1 vccd1 vccd1 _08810_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09787_ _09787_/A _09787_/B _09787_/C vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__or3_1
XFILLER_39_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06999_ _07007_/A _07570_/C vssd1 vssd1 vccd1 vccd1 _07000_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08738_ _10537_/A _08694_/X _08695_/X _10806_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08738_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _10799_/Q _08669_/B _08669_/C vssd1 vssd1 vccd1 vccd1 _08670_/C sky130_fd_sc_hd__nand3_1
XFILLER_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10700_ _10700_/CLK _10700_/D vssd1 vssd1 vccd1 vccd1 _10700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A2 _08672_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10631_ _10811_/CLK _10631_/D vssd1 vssd1 vccd1 vccd1 _10631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10562_ _10673_/CLK _10562_/D vssd1 vssd1 vccd1 vccd1 _10562_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06127__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10493_/X sky130_fd_sc_hd__or2_1
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08342__A _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 _10981_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08517__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09076__C1 _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10829_ _10847_/CLK _10829_/D vssd1 vssd1 vccd1 vccd1 _10829_/Q sky130_fd_sc_hd__dfxtp_1
X_06020_ _08258_/A vssd1 vssd1 vccd1 vccd1 _06020_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07971_ _10517_/A _09263_/A vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__nor2_1
X_09710_ _09710_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09711_/B sky130_fd_sc_hd__and2_1
X_06922_ _06922_/A _06922_/B vssd1 vssd1 vccd1 vccd1 _06926_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08354__A1 _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08354__B2 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09641_ _09641_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__xor2_1
X_06853_ _06853_/A _06853_/B vssd1 vssd1 vccd1 vccd1 _07780_/B sky130_fd_sc_hd__nor2_1
X_05804_ _08321_/A _05769_/A _10566_/Q _05781_/Y vssd1 vssd1 vccd1 vccd1 _05804_/X
+ sky130_fd_sc_hd__a22o_1
X_09572_ _10115_/A vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06784_ _06828_/A _06828_/B vssd1 vssd1 vccd1 vccd1 _06882_/A sky130_fd_sc_hd__or2_1
XFILLER_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05735_ _08093_/A _05547_/A _05536_/B _05733_/X _05734_/X vssd1 vssd1 vccd1 vccd1
+ _05788_/B sky130_fd_sc_hd__o221ai_2
X_08523_ _08935_/A _10762_/Q vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__and2_1
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09811__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05666_ _10693_/Q _05664_/Y _05615_/Y _05877_/A vssd1 vssd1 vccd1 vccd1 _05666_/X
+ sky130_fd_sc_hd__a22o_1
X_08454_ _08454_/A vssd1 vssd1 vccd1 vccd1 _10735_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05597_ _10700_/Q vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08385_ _10198_/A vssd1 vssd1 vccd1 vccd1 _08395_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07405_ _07405_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _07540_/A sky130_fd_sc_hd__or2_1
XFILLER_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07336_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07522_/B sky130_fd_sc_hd__and2_1
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07985__B _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09006_ _10069_/A vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__clkbuf_4
X_07267_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__or2_1
XFILLER_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06218_ _10601_/Q _06223_/B vssd1 vssd1 vccd1 vccd1 _06218_/X sky130_fd_sc_hd__or2_1
X_07198_ _07193_/A _07193_/B _07194_/B _07210_/A _07260_/A vssd1 vssd1 vccd1 vccd1
+ _07277_/B sky130_fd_sc_hd__a32o_1
XFILLER_117_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06149_ _06149_/A vssd1 vssd1 vccd1 vccd1 _06238_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10842__D _10842_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08345__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _09908_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _10049_/C sky130_fd_sc_hd__nand2_1
XFILLER_86_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09839_ _09974_/A _09839_/B _09839_/C vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__and3_1
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10614_ _10851_/CLK _10614_/D vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10545_ _10654_/CLK _10545_/D vssd1 vssd1 vccd1 vccd1 _10545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10476_ _10517_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10493_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10391__A1 _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05520_ _05329_/X _05517_/X _05513_/X _07914_/A vssd1 vssd1 vccd1 vccd1 _10568_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_05451_ _10620_/Q vssd1 vssd1 vccd1 vccd1 _05453_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08170_ _08180_/B vssd1 vssd1 vccd1 vccd1 _08181_/B sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_46_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05382_ _10656_/Q _05382_/B vssd1 vssd1 vccd1 vccd1 _05383_/B sky130_fd_sc_hd__nand2_1
X_07121_ _07145_/A _07145_/B vssd1 vssd1 vccd1 vccd1 _07136_/A sky130_fd_sc_hd__and2b_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07052_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__nand2_1
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06003_ _06003_/A vssd1 vssd1 vccd1 vccd1 _10577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07954_ input43/X _06038_/X _07983_/A vssd1 vssd1 vccd1 vccd1 _07955_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07885_ _07885_/A vssd1 vssd1 vccd1 vccd1 _07885_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_56_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06905_ _06567_/B _06368_/B _06895_/B vssd1 vssd1 vccd1 vccd1 _06922_/B sky130_fd_sc_hd__a21oi_4
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09624_ _09624_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__and2_2
X_06836_ _06836_/A vssd1 vssd1 vccd1 vccd1 _06836_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06767_ _06775_/A vssd1 vssd1 vccd1 vccd1 _06900_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _09555_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08157__A _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05718_ _05718_/A vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__clkbuf_2
X_08506_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08506_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _09486_/A _09486_/B vssd1 vssd1 vccd1 vccd1 _09562_/A sky130_fd_sc_hd__xnor2_1
X_06698_ _06697_/B _06698_/B vssd1 vssd1 vccd1 vccd1 _06698_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10837__D _10837_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05649_ _05719_/A _05641_/Y _05648_/X vssd1 vssd1 vccd1 vccd1 _05649_/X sky130_fd_sc_hd__a21o_1
X_08437_ _08437_/A vssd1 vssd1 vccd1 vccd1 _10730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07996__A _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08368_ _10729_/Q vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__clkbuf_4
X_08299_ _08305_/B _08253_/X _08297_/Y _08298_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08299_/X sky130_fd_sc_hd__a311o_1
X_07319_ _07319_/A _07319_/B vssd1 vssd1 vccd1 vccd1 _07341_/B sky130_fd_sc_hd__or2_1
XFILLER_125_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10330_ _10330_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10330_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10261_ _10261_/A _10261_/B vssd1 vssd1 vccd1 vccd1 _10261_/X sky130_fd_sc_hd__xor2_1
XFILLER_120_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09716__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10192_ _10192_/A vssd1 vssd1 vccd1 vccd1 _10192_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06041__A2 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput25 io_wbs_m2s_data[18] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_8
XFILLER_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 io_wbs_m2s_addr[8] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput36 io_wbs_m2s_data[28] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_6
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput47 io_wbs_m2s_data[9] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_4
X_10528_ _10528_/A _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10528_/X sky130_fd_sc_hd__or3_1
XFILLER_124_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10459_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10116__A1 _10109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07670_ _07670_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07671_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06621_ _06621_/A _06621_/B vssd1 vssd1 vccd1 vccd1 _06692_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06552_ _10971_/Q vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__inv_2
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09340_ _06993_/A _10894_/Q vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__and2b_1
X_05503_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05503_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09271_ _10825_/Q _09243_/X _09244_/X _09269_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09272_/B sky130_fd_sc_hd__a32o_1
XFILLER_61_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08222_ input23/X _08164_/X _08165_/X _08216_/X _08394_/A vssd1 vssd1 vccd1 vccd1
+ _08222_/X sky130_fd_sc_hd__o221a_1
X_06483_ _06646_/A _06646_/B vssd1 vssd1 vccd1 vccd1 _06647_/A sky130_fd_sc_hd__nor2_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05434_ _07896_/A _05343_/Y _05431_/X _05433_/X vssd1 vssd1 vccd1 vccd1 _05434_/X
+ sky130_fd_sc_hd__a22o_1
X_08153_ _07976_/A _08043_/A _08152_/X _08038_/A _08096_/A vssd1 vssd1 vccd1 vccd1
+ _08155_/A sky130_fd_sc_hd__a221o_1
XFILLER_119_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05365_ _10662_/Q vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__buf_2
X_08084_ _08113_/A _08081_/X _08083_/Y _06024_/A vssd1 vssd1 vccd1 vccd1 _08084_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_119_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07104_ _07142_/B vssd1 vssd1 vccd1 vccd1 _07394_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05296_ _10656_/Q _05382_/B vssd1 vssd1 vccd1 vccd1 _05383_/A sky130_fd_sc_hd__or2_1
XANTENNA__06225__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07035_ _07035_/A _07415_/C vssd1 vssd1 vccd1 vccd1 _07037_/B sky130_fd_sc_hd__xor2_1
XFILLER_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08986_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__and2_1
X_07937_ input16/X _05475_/X _07964_/A vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__mux2_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07868_ _07848_/X _05460_/B _07865_/X hold15/X vssd1 vssd1 vccd1 vccd1 _10630_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06819_ _10502_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _07779_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _09607_/A _09676_/D vssd1 vssd1 vccd1 vccd1 _09608_/B sky130_fd_sc_hd__xor2_2
X_07799_ _07799_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _07799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09538_ _09538_/A _09638_/C vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__and2_1
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09469_ _09534_/C _09469_/B vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__nand2_1
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08787__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06135__A _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10313_ _09920_/B _10283_/X _10312_/X _10293_/X vssd1 vssd1 vccd1 vccd1 _10910_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10244_ _10953_/Q _10937_/Q vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__and2b_1
XFILLER_78_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10175_ _07066_/A _10174_/X _10170_/X _10887_/Q vssd1 vssd1 vccd1 vccd1 _10887_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08711__A1 _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08244__B _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08840_ _10819_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08844_/A sky130_fd_sc_hd__xnor2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05983_ _08445_/A vssd1 vssd1 vccd1 vccd1 _05983_/X sky130_fd_sc_hd__buf_4
X_08771_ _08771_/A _08796_/B vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__nand2_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07722_ _07585_/A _07721_/Y _07584_/A vssd1 vssd1 vccd1 vccd1 _07741_/A sky130_fd_sc_hd__a21oi_1
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07653_ _07653_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07654_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06604_ _06593_/A _06593_/B _06593_/C vssd1 vssd1 vccd1 vccd1 _06605_/B sky130_fd_sc_hd__a21oi_1
XFILLER_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09323_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09324_/B sky130_fd_sc_hd__or2_1
X_07584_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__or2_2
X_06535_ _06534_/B _06535_/B vssd1 vssd1 vccd1 vccd1 _06536_/B sky130_fd_sc_hd__and2b_1
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09254_ _09259_/A _09254_/B vssd1 vssd1 vccd1 vccd1 _09255_/A sky130_fd_sc_hd__and2_4
X_06466_ _06480_/C _06466_/B vssd1 vssd1 vccd1 vccd1 _06688_/A sky130_fd_sc_hd__or2_1
XFILLER_138_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08205_ _08206_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08224_/C sky130_fd_sc_hd__and2_1
X_05417_ _05462_/B _05389_/Y _05385_/Y _10623_/Q _05416_/X vssd1 vssd1 vccd1 vccd1
+ _05417_/X sky130_fd_sc_hd__a221o_1
X_09185_ _10961_/Q _09194_/B vssd1 vssd1 vccd1 vccd1 _09185_/Y sky130_fd_sc_hd__nor2_1
X_08136_ _08132_/A _08132_/B _06035_/A vssd1 vssd1 vccd1 vccd1 _08136_/Y sky130_fd_sc_hd__o21ai_1
X_06397_ _10977_/Q vssd1 vssd1 vccd1 vccd1 _06456_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_134_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05348_ _05854_/A _05348_/B vssd1 vssd1 vccd1 vccd1 _05348_/X sky130_fd_sc_hd__and2_1
X_08067_ _08092_/A vssd1 vssd1 vccd1 vccd1 _08067_/X sky130_fd_sc_hd__buf_2
X_05279_ _05279_/A vssd1 vssd1 vccd1 vccd1 _05818_/A sky130_fd_sc_hd__clkinv_2
XFILLER_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07018_ _07229_/A vssd1 vssd1 vccd1 vccd1 _07416_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08969_ _09142_/B _09142_/C _08965_/B _08968_/X vssd1 vssd1 vccd1 vccd1 _08969_/Y
+ sky130_fd_sc_hd__o31ai_4
XFILLER_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09205__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10931_ _10935_/CLK _10931_/D vssd1 vssd1 vccd1 vccd1 _10931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10862_ _10862_/CLK _10862_/D vssd1 vssd1 vccd1 vccd1 _10862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _10797_/CLK _10793_/D vssd1 vssd1 vccd1 vccd1 _10793_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05969__A _08414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10227_ _10226_/B _10217_/X _10214_/A vssd1 vssd1 vccd1 vccd1 _10228_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10115__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06312__B _10909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10158_ _10158_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__xnor2_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10089_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10090_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06171__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06320_ _10924_/Q _10907_/Q vssd1 vssd1 vccd1 vccd1 _06320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06251_ hold25/A _06253_/B vssd1 vssd1 vccd1 vccd1 _06251_/X sky130_fd_sc_hd__or2_1
XFILLER_90_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06182_ input17/X vssd1 vssd1 vccd1 vccd1 _06182_/X sky130_fd_sc_hd__buf_4
XANTENNA__09948__B1 _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _10009_/B _09941_/B vssd1 vssd1 vccd1 vccd1 _09943_/C sky130_fd_sc_hd__and2_1
XANTENNA__10025__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09872_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__nor2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _10817_/Q _08865_/B vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__nand2_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08754_ _06178_/X _08694_/X _08695_/X _10808_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08754_/X sky130_fd_sc_hd__o221a_1
X_05966_ _09016_/A _09126_/A vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__or2_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07705_ _07616_/X _09899_/B _07704_/Y vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__a21bo_1
X_05897_ _10656_/Q _05900_/A vssd1 vssd1 vccd1 vccd1 _05897_/X sky130_fd_sc_hd__xor2_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08685_ _08683_/X _08684_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10801_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07636_ _07636_/A _07636_/B vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__xor2_4
XFILLER_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07567_ _07567_/A vssd1 vssd1 vccd1 vccd1 _07726_/A sky130_fd_sc_hd__clkbuf_4
X_06518_ _06521_/A _06521_/B _06612_/A _06503_/Y vssd1 vssd1 vccd1 vccd1 _06519_/B
+ sky130_fd_sc_hd__a211oi_1
X_09306_ _09306_/A _09316_/A vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__or2_1
XANTENNA__10845__D _10845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08165__A _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09237_ _08267_/A _07893_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09237_/X sky130_fd_sc_hd__mux2_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07498_ _07534_/B _07534_/C _07534_/A vssd1 vssd1 vccd1 vccd1 _07535_/A sky130_fd_sc_hd__o21a_1
X_06449_ _06472_/A _06470_/A _06426_/A _06568_/B vssd1 vssd1 vccd1 vccd1 _06450_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09168_ _09168_/A vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ _08119_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _10493_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__nor2_2
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10580__D _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10012_ _10012_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__nor2_1
XFILLER_130_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input15_A io_wbs_m2s_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08059__B _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ _10955_/CLK _10914_/D vssd1 vssd1 vccd1 vccd1 _10914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10845_ _10845_/CLK _10845_/D vssd1 vssd1 vccd1 vccd1 _10845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10776_ _10836_/CLK _10776_/D vssd1 vssd1 vccd1 vccd1 _10776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06307__B _10906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09634__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05820_ _05905_/A _05905_/B vssd1 vssd1 vccd1 vccd1 _05906_/A sky130_fd_sc_hd__or2_1
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05751_ _10700_/Q vssd1 vssd1 vccd1 vccd1 _05751_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05682_ _10707_/Q vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__clkbuf_2
X_08470_ _10777_/Q _10740_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__mux2_1
XFILLER_63_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06993__A _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07421_ _07421_/A vssd1 vssd1 vccd1 vccd1 _07421_/Y sky130_fd_sc_hd__inv_2
XFILLER_23_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07352_ _07366_/B _07291_/B _07291_/C vssd1 vssd1 vccd1 vccd1 _07353_/B sky130_fd_sc_hd__a21oi_1
X_06303_ _06303_/A _06305_/C vssd1 vssd1 vccd1 vccd1 _06730_/B sky130_fd_sc_hd__or2_1
X_07283_ _07357_/C _07283_/B vssd1 vssd1 vccd1 vccd1 _07284_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09022_ _06065_/X _08976_/X _09020_/X _09021_/Y _09078_/B vssd1 vssd1 vccd1 vccd1
+ _09022_/X sky130_fd_sc_hd__a221o_1
X_06234_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06234_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06165_ _06165_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06096_ _10685_/Q _10684_/Q _08098_/B vssd1 vssd1 vccd1 vccd1 _08117_/B sky130_fd_sc_hd__or3_2
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06080__B1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09924_ _10131_/A _09924_/B vssd1 vssd1 vccd1 vccd1 _09925_/B sky130_fd_sc_hd__nand2_1
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09855_ _09855_/A _09855_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__xor2_2
XANTENNA_input7_A io_wbs_m2s_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08806_ _08806_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _08806_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09786_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09787_/C sky130_fd_sc_hd__xnor2_1
X_06998_ _07028_/A _07008_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07570_/C sky130_fd_sc_hd__or3_1
X_05949_ _08350_/A _05829_/X _05826_/X _05528_/X _05948_/X vssd1 vssd1 vccd1 vccd1
+ _05949_/X sky130_fd_sc_hd__o221a_1
X_08737_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08737_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _08669_/B _08669_/C _10799_/Q vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__a21o_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07619_ _07625_/A _07624_/B _07624_/A vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__a21oi_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10811_/CLK _10630_/D vssd1 vssd1 vccd1 vccd1 _10630_/Q sky130_fd_sc_hd__dfxtp_1
X_08599_ _09403_/B _08624_/B vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__or2_2
XANTENNA__05312__A _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ _10673_/CLK _10561_/D vssd1 vssd1 vccd1 vccd1 _10561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ _06163_/X _10489_/B _10491_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10969_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05949__B2 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06143__A _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05982__A _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10828_ _10830_/CLK _10828_/D vssd1 vssd1 vccd1 vccd1 _10828_/Q sky130_fd_sc_hd__dfxtp_1
X_10759_ _10798_/CLK _10759_/D vssd1 vssd1 vccd1 vccd1 _10759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08533__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10695_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09348__B _10907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06062__B1 _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07970_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06921_ _06921_/A _06921_/B vssd1 vssd1 vccd1 vccd1 _06922_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_42_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10830_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_95_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06852_ _06852_/A _06852_/B vssd1 vssd1 vccd1 vccd1 _06855_/A sky130_fd_sc_hd__xor2_2
X_09640_ _09640_/A _09640_/B vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__xnor2_1
X_05803_ _05803_/A vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__inv_2
X_09571_ hold12/A _09408_/X _09570_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10872_/D
+ sky130_fd_sc_hd__a22o_1
X_06783_ _06902_/A _06892_/B _06782_/A vssd1 vssd1 vccd1 vccd1 _06828_/B sky130_fd_sc_hd__a21oi_1
X_05734_ _05726_/A _05549_/A _05729_/Y _05728_/X vssd1 vssd1 vccd1 vccd1 _05734_/X
+ sky130_fd_sc_hd__o22a_1
X_08522_ _08522_/A vssd1 vssd1 vccd1 vccd1 _10762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08453_ _08460_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__or2_1
XFILLER_24_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05665_ _05885_/A _05619_/X _05664_/Y _10693_/Q vssd1 vssd1 vccd1 vccd1 _05665_/X
+ sky130_fd_sc_hd__o22a_1
X_07404_ _07404_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _07405_/B sky130_fd_sc_hd__and2_1
XFILLER_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05596_ _05596_/A _05596_/B vssd1 vssd1 vccd1 vccd1 _05596_/X sky130_fd_sc_hd__and2_1
X_08384_ _10251_/S vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__buf_4
XFILLER_51_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07335_ _07335_/A _07335_/B vssd1 vssd1 vccd1 vccd1 _07511_/B sky130_fd_sc_hd__and2_1
XFILLER_109_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07266_ _07266_/A _07270_/A vssd1 vssd1 vccd1 vccd1 _07268_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08443__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06217_ input23/X _06207_/X _06216_/X _06200_/X vssd1 vssd1 vccd1 vccd1 _10600_/D
+ sky130_fd_sc_hd__o211a_1
X_09005_ _09931_/A vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__buf_2
X_07197_ _07197_/A _07197_/B _07197_/C vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__and3_1
X_06148_ _10587_/Q vssd1 vssd1 vccd1 vccd1 _06151_/A sky130_fd_sc_hd__inv_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06079_ _06113_/A _08342_/A _06038_/X _08105_/A _06078_/X vssd1 vssd1 vccd1 vccd1
+ _06082_/C sky130_fd_sc_hd__a221o_1
XFILLER_78_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09274__A _09274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09907_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08345__A2 _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09838_ _09906_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09839_/C sky130_fd_sc_hd__and2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09769_ _09769_/A _09769_/B _09769_/C vssd1 vssd1 vccd1 vccd1 _09771_/C sky130_fd_sc_hd__and3_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10613_ _10851_/CLK _10613_/D vssd1 vssd1 vccd1 vccd1 _10613_/Q sky130_fd_sc_hd__dfxtp_1
X_10544_ _10651_/CLK _10544_/D vssd1 vssd1 vccd1 vccd1 _10544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08281__B2 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ _10489_/B vssd1 vssd1 vccd1 vccd1 _10475_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08033__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06044__B1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10123__A _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06320__B _10907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09297__A0 _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05450_ _05490_/A vssd1 vssd1 vccd1 vccd1 _05470_/A sky130_fd_sc_hd__inv_2
XFILLER_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05381_ _10625_/Q vssd1 vssd1 vccd1 vccd1 _05461_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07120_ _07135_/A _07511_/A _07149_/C _07235_/B vssd1 vssd1 vccd1 vccd1 _07145_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08263__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07051_ _07051_/A _07414_/A vssd1 vssd1 vccd1 vccd1 _07371_/B sky130_fd_sc_hd__xnor2_1
XFILLER_126_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08024__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A0 _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06002_ _08483_/A _06002_/B vssd1 vssd1 vccd1 vccd1 _06003_/A sky130_fd_sc_hd__and2_1
XFILLER_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07953_ _07953_/A vssd1 vssd1 vccd1 vccd1 _10652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07884_ _07898_/A _07884_/B vssd1 vssd1 vccd1 vccd1 _10634_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06904_ _06921_/A _06921_/B vssd1 vssd1 vccd1 vccd1 _06904_/X sky130_fd_sc_hd__or2_1
XFILLER_110_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06835_ _06835_/A _06835_/B vssd1 vssd1 vccd1 vccd1 _06839_/A sky130_fd_sc_hd__xnor2_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ _09623_/A _09623_/B _09623_/C vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__or3_1
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06766_ _06766_/A _06766_/B vssd1 vssd1 vccd1 vccd1 _06828_/A sky130_fd_sc_hd__or2_1
X_09554_ _09805_/A _09692_/A _09554_/C vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__and3_1
X_05717_ _05798_/A _05717_/B _05717_/C _05717_/D vssd1 vssd1 vccd1 vccd1 _05717_/X
+ sky130_fd_sc_hd__or4_1
X_08505_ _10788_/Q _08496_/X _08502_/X hold26/A vssd1 vssd1 vccd1 vccd1 _10751_/D
+ sky130_fd_sc_hd__a22o_1
X_09485_ _09904_/A _09744_/A vssd1 vssd1 vccd1 vccd1 _09486_/B sky130_fd_sc_hd__nand2_1
X_06697_ _06698_/B _06697_/B vssd1 vssd1 vccd1 vccd1 _06912_/B sky130_fd_sc_hd__xnor2_2
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05648_ _05719_/A _05641_/Y _05644_/Y _08082_/C _05647_/X vssd1 vssd1 vccd1 vccd1
+ _05648_/X sky130_fd_sc_hd__o221a_1
X_08436_ _08443_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__or2_1
X_08367_ _08419_/A vssd1 vssd1 vccd1 vccd1 _08367_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05579_ _10566_/Q _05588_/A vssd1 vssd1 vccd1 vccd1 _05580_/B sky130_fd_sc_hd__nand2_1
X_07318_ _07318_/A _07318_/B _07324_/A vssd1 vssd1 vccd1 vccd1 _07319_/B sky130_fd_sc_hd__and3_1
XFILLER_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08298_ _08298_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08298_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07926__A2_N _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ _07517_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _07250_/B sky130_fd_sc_hd__and2b_1
XFILLER_124_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10260_ _10258_/Y _10259_/X _10291_/S vssd1 vssd1 vccd1 vccd1 _10261_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08901__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10191_ _10197_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10198_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07951__S _07983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06140__B _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08348__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput37 io_wbs_m2s_data[29] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_6
Xinput26 io_wbs_m2s_data[19] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_6
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput15 io_wbs_m2s_addr[9] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_4
Xinput48 io_wbs_m2s_sel[0] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
X_10527_ _07726_/A _10522_/X _10526_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10981_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10458_ _06178_/X _10446_/X _10456_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10956_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06315__B _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10389_ _10408_/A vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10521__C1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ _06620_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _06621_/B sky130_fd_sc_hd__and2_1
XFILLER_65_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06551_ _06561_/B _06561_/C _06587_/B vssd1 vssd1 vccd1 vccd1 _06564_/A sky130_fd_sc_hd__and3_1
X_05502_ _05366_/Y _05497_/X _05490_/A _05460_/B vssd1 vssd1 vccd1 vccd1 _10555_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09270_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09270_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06482_ _06658_/A _06657_/B _06657_/A vssd1 vssd1 vccd1 vccd1 _06646_/B sky130_fd_sc_hd__o21ba_1
X_08221_ _08216_/X _08224_/C _08220_/Y vssd1 vssd1 vccd1 vccd1 _08221_/Y sky130_fd_sc_hd__a21oi_1
X_05433_ _10638_/Q _05343_/Y _05348_/X _07893_/A vssd1 vssd1 vccd1 vccd1 _05433_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08065_/B _08147_/X _08149_/Y _08151_/Y _08074_/A vssd1 vssd1 vccd1 vccd1
+ _08152_/X sky130_fd_sc_hd__a32o_1
XFILLER_119_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05364_ _10630_/Q vssd1 vssd1 vccd1 vccd1 _05460_/B sky130_fd_sc_hd__clkbuf_2
X_08083_ _08095_/B vssd1 vssd1 vccd1 vccd1 _08083_/Y sky130_fd_sc_hd__inv_2
X_05295_ _05295_/A _05389_/A vssd1 vssd1 vccd1 vccd1 _05382_/B sky130_fd_sc_hd__nand2_1
X_07103_ _07382_/A vssd1 vssd1 vccd1 vccd1 _07142_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_134_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07034_ _07043_/A _07034_/B vssd1 vssd1 vccd1 vccd1 _07415_/C sky130_fd_sc_hd__xnor2_1
XFILLER_115_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08985_ _09168_/A vssd1 vssd1 vccd1 vccd1 _08985_/X sky130_fd_sc_hd__clkbuf_2
X_07936_ _07950_/A vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__buf_2
XFILLER_102_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07867_ _06204_/A _07849_/X _07850_/X _07866_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ hold15/A sky130_fd_sc_hd__o221ai_4
XFILLER_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06818_ _06818_/A _06818_/B vssd1 vssd1 vccd1 vccd1 _07767_/B sky130_fd_sc_hd__xnor2_4
X_09606_ _09369_/X _09606_/B vssd1 vssd1 vccd1 vccd1 _09676_/D sky130_fd_sc_hd__and2b_1
X_07798_ _07798_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _07802_/A sky130_fd_sc_hd__xnor2_1
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09537_ _09538_/A _09638_/C vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__nor2_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06749_ _06769_/A _06758_/C vssd1 vssd1 vccd1 vccd1 _06772_/A sky130_fd_sc_hd__and2_1
XANTENNA__10848__D _10848_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _09534_/C _09469_/B vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__or2_1
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08419_ _08419_/A _08419_/B vssd1 vssd1 vccd1 vccd1 _08419_/Y sky130_fd_sc_hd__nand2_1
X_09399_ _09400_/B _09399_/B vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__and2b_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ _10312_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10312_/X sky130_fd_sc_hd__xor2_1
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10243_ _10243_/A vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__inv_2
XANTENNA_input45_A io_wbs_m2s_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10174_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10174_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_120_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05289__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10282__A1 _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08525__B _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06061__A _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05982_ _05982_/A _05993_/S vssd1 vssd1 vccd1 vccd1 _05982_/Y sky130_fd_sc_hd__nor2_1
X_08770_ _10811_/Q vssd1 vssd1 vccd1 vccd1 _08771_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06996__A _10907_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07721_ _07721_/A vssd1 vssd1 vccd1 vccd1 _07721_/Y sky130_fd_sc_hd__inv_2
XFILLER_65_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07652_ _07653_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07654_/A sky130_fd_sc_hd__or2_1
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05405__A _05405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06603_ _06616_/A _06616_/B vssd1 vssd1 vccd1 vccd1 _06672_/A sky130_fd_sc_hd__xor2_1
X_07583_ _07582_/B _07583_/B vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__and2b_1
X_09322_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__nand2_1
X_06534_ _06535_/B _06534_/B vssd1 vssd1 vccd1 vccd1 _06536_/A sky130_fd_sc_hd__and2b_1
XFILLER_61_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ _10822_/Q _09243_/X _09244_/X _09252_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09254_/B sky130_fd_sc_hd__a32o_1
XFILLER_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10273__A1 _06997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06465_ _06465_/A _06465_/B vssd1 vssd1 vccd1 vccd1 _06466_/B sky130_fd_sc_hd__nor2_1
X_08204_ _08204_/A vssd1 vssd1 vccd1 vccd1 _10694_/D sky130_fd_sc_hd__clkbuf_1
X_05416_ _10622_/Q _05389_/Y _05393_/X _05415_/X vssd1 vssd1 vccd1 vccd1 _05416_/X
+ sky130_fd_sc_hd__o22a_1
X_09184_ _09202_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _10847_/D sky130_fd_sc_hd__nor2_2
X_06396_ _06396_/A vssd1 vssd1 vccd1 vccd1 _06871_/A sky130_fd_sc_hd__clkinv_2
X_08135_ _08131_/X _08133_/X _08134_/X vssd1 vssd1 vccd1 vccd1 _10687_/D sky130_fd_sc_hd__o21a_1
X_05347_ _10669_/Q _05347_/B vssd1 vssd1 vccd1 vccd1 _05348_/B sky130_fd_sc_hd__nand2_1
XFILLER_107_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08066_ _08113_/A vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__clkbuf_2
X_05278_ _10651_/Q vssd1 vssd1 vccd1 vccd1 _05279_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__05988__C1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ _07186_/A vssd1 vssd1 vccd1 vccd1 _07229_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08968_ _08968_/A vssd1 vssd1 vccd1 vccd1 _08968_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07919_ _07919_/A vssd1 vssd1 vccd1 vccd1 _07919_/Y sky130_fd_sc_hd__clkinv_2
X_08899_ input35/X _08785_/X _08786_/X _10826_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08899_/X sky130_fd_sc_hd__o221a_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10930_ _10930_/CLK _10930_/D vssd1 vssd1 vccd1 vccd1 _10930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05315__A _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10861_ _10865_/CLK _10861_/D vssd1 vssd1 vccd1 vccd1 _10861_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09221__S _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10792_ _10797_/CLK _10792_/D vssd1 vssd1 vccd1 vccd1 _10792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05969__B _08939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05985__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10226_ _10226_/A _10226_/B _10226_/C vssd1 vssd1 vccd1 vccd1 _10226_/X sky130_fd_sc_hd__and3_1
XFILLER_121_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10157_ _10157_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__xnor2_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_67_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10088_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__or2_1
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08696__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08536__A _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06250_ input37/X _06238_/X _06249_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10613_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_90_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06056__A _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06181_ _06178_/X _06158_/X _06180_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10593_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09940_ _09940_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09871_ _09933_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__nand2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08822_ _08814_/X _08817_/X _08818_/Y _08821_/X vssd1 vssd1 vccd1 vccd1 _10816_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_58_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08753_ _08759_/B _08753_/B vssd1 vssd1 vccd1 vccd1 _08753_/Y sky130_fd_sc_hd__xnor2_1
X_05965_ input8/X _09142_/C vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__or2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08136__B1 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07704_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _07704_/Y sky130_fd_sc_hd__nand2_1
X_05896_ _05896_/A vssd1 vssd1 vccd1 vccd1 _06035_/A sky130_fd_sc_hd__buf_2
X_08684_ _10526_/A _08672_/X _08674_/X _10801_/Q vssd1 vssd1 vccd1 vccd1 _08684_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10494__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07635_ _07635_/A _07635_/B vssd1 vssd1 vccd1 vccd1 _07636_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__xnor2_1
X_06517_ _06517_/A _06517_/B _06517_/C vssd1 vssd1 vccd1 vccd1 _06612_/A sky130_fd_sc_hd__and3_1
X_09305_ _10898_/Q _10882_/Q vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__and2b_4
X_09236_ _09236_/A vssd1 vssd1 vccd1 vccd1 _10854_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_37_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07497_ _07497_/A _07497_/B vssd1 vssd1 vccd1 vccd1 _07534_/A sky130_fd_sc_hd__xor2_1
X_06448_ _06469_/B _06448_/B vssd1 vssd1 vccd1 vccd1 _06470_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _09113_/X _09166_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09167_/Y sky130_fd_sc_hd__o21ai_1
X_06379_ _06408_/B _06409_/C _06393_/A vssd1 vssd1 vccd1 vccd1 _06381_/C sky130_fd_sc_hd__a21oi_1
XFILLER_135_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08118_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__buf_2
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09098_ _09098_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__or2_2
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08049_ input8/X _09124_/C vssd1 vssd1 vccd1 vccd1 _08416_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08375__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _10012_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10081_/B sky130_fd_sc_hd__and2_1
XFILLER_0_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06015__D_N input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _10920_/CLK _10913_/D vssd1 vssd1 vccd1 vccd1 _10913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10844_ _10848_/CLK _10844_/D vssd1 vssd1 vccd1 vccd1 _10844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10775_ _10781_/CLK _10775_/D vssd1 vssd1 vccd1 vccd1 _10775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06323__B _10909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10209_ _10202_/X _10203_/X _10208_/X vssd1 vssd1 vccd1 vccd1 _10209_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07435__A _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05750_ _05744_/Y _10557_/Q _05747_/X _05749_/X vssd1 vssd1 vccd1 vccd1 _05750_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_82_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05681_ _10568_/Q _05681_/B vssd1 vssd1 vccd1 vccd1 _05684_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07420_ _07555_/B _07418_/Y _07419_/X vssd1 vssd1 vccd1 vccd1 _07426_/A sky130_fd_sc_hd__o21ai_1
XFILLER_35_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07351_ _07470_/B _07482_/A _07470_/A vssd1 vssd1 vccd1 vccd1 _07471_/A sky130_fd_sc_hd__o21a_1
X_06302_ _06386_/A _06302_/B _06416_/A vssd1 vssd1 vccd1 vccd1 _06305_/C sky130_fd_sc_hd__or3b_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07282_ _07282_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _07291_/B sky130_fd_sc_hd__or2_1
XFILLER_129_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09021_ _06066_/Y _06212_/B _08995_/X vssd1 vssd1 vccd1 vccd1 _09021_/Y sky130_fd_sc_hd__a21oi_1
X_06233_ _10607_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06233_/X sky130_fd_sc_hd__or2_1
XFILLER_117_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06164_ _10590_/Q vssd1 vssd1 vccd1 vccd1 _06165_/A sky130_fd_sc_hd__inv_2
XANTENNA__10400__A1 _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06095_ _10683_/Q _10682_/Q _08075_/B vssd1 vssd1 vccd1 vccd1 _08098_/B sky130_fd_sc_hd__or3_2
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09923_ _09923_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09924_/B sky130_fd_sc_hd__or2_1
XFILLER_112_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09854_ _09795_/A _09795_/B _09853_/Y vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__a21bo_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08805_ _10814_/Q _10813_/Q _10812_/Q _08771_/A _08801_/B vssd1 vssd1 vccd1 vccd1
+ _08806_/B sky130_fd_sc_hd__o41a_1
XFILLER_58_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09661_/X _09724_/A _09723_/Y vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__o21ai_1
XFILLER_39_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06997_ _07013_/A _06997_/B _06997_/C vssd1 vssd1 vccd1 vccd1 _07007_/B sky130_fd_sc_hd__or3_1
X_05948_ _08350_/A _05829_/X _05946_/X _05947_/X vssd1 vssd1 vccd1 vccd1 _05948_/X
+ sky130_fd_sc_hd__a22o_1
X_08736_ _08740_/C _08736_/B vssd1 vssd1 vccd1 vccd1 _08736_/X sky130_fd_sc_hd__xor2_1
X_05879_ _10661_/Q vssd1 vssd1 vccd1 vccd1 _07988_/A sky130_fd_sc_hd__buf_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _10800_/Q _08678_/A vssd1 vssd1 vccd1 vccd1 _08669_/C sky130_fd_sc_hd__or2_1
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07618_ _07618_/A _07618_/B vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__xor2_2
XANTENNA__05894__A1 _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08598_ _10283_/A vssd1 vssd1 vccd1 vccd1 _08649_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10856__D _10856_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07549_ _07549_/A _07549_/B vssd1 vssd1 vccd1 vccd1 _07550_/B sky130_fd_sc_hd__and2_1
XFILLER_14_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ _10702_/CLK _10560_/D vssd1 vssd1 vccd1 vccd1 _10560_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08832__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09245_/S sky130_fd_sc_hd__clkbuf_2
X_10491_ _10491_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__or2_1
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__S _07983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08899__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10458__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08520__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07702__B _07702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05503__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10827_ _10847_/CLK _10827_/D vssd1 vssd1 vccd1 vccd1 _10827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10758_ _10798_/CLK _10758_/D vssd1 vssd1 vccd1 vccd1 _10758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10689_ _10841_/CLK _10689_/D vssd1 vssd1 vccd1 vccd1 _10689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06920_ _06939_/A _06939_/B vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__nor2_2
XFILLER_95_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06851_ _06851_/A _06851_/B vssd1 vssd1 vccd1 vccd1 _06852_/B sky130_fd_sc_hd__nand2_1
X_05802_ _05802_/A _05802_/B vssd1 vssd1 vccd1 vccd1 _05802_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09570_ _09570_/A _09574_/B vssd1 vssd1 vccd1 vccd1 _09570_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06782_ _06782_/A _06782_/B vssd1 vssd1 vccd1 vccd1 _06892_/B sky130_fd_sc_hd__nor2_2
X_05733_ _08082_/A vssd1 vssd1 vccd1 vccd1 _05733_/X sky130_fd_sc_hd__clkbuf_2
X_08521_ _08935_/A input3/X vssd1 vssd1 vccd1 vccd1 _08522_/A sky130_fd_sc_hd__and2_1
XFILLER_82_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10449__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08452_ _10772_/Q _10735_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08453_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05664_ _05664_/A _05664_/B vssd1 vssd1 vccd1 vccd1 _05664_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07403_ _07404_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__nor2_1
X_05595_ _10561_/Q _05602_/A _10562_/Q vssd1 vssd1 vccd1 vccd1 _05596_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09067__A1 _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _08419_/A vssd1 vssd1 vccd1 vccd1 _08383_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07334_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07335_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07265_ _07269_/A _07514_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__a21oi_1
X_06216_ _10600_/Q _06223_/B vssd1 vssd1 vccd1 vccd1 _06216_/X sky130_fd_sc_hd__or2_1
X_09004_ _09867_/A vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_0_clock_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07196_ _07196_/A _07196_/B vssd1 vssd1 vccd1 vccd1 _07197_/C sky130_fd_sc_hd__xor2_1
XFILLER_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06147_ _10528_/A vssd1 vssd1 vccd1 vccd1 _06147_/X sky130_fd_sc_hd__clkbuf_4
X_06078_ _08251_/B _08244_/A vssd1 vssd1 vccd1 vccd1 _06078_/X sky130_fd_sc_hd__xor2_1
X_09906_ _09906_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__xor2_1
XFILLER_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09837_ _09837_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09838_/B sky130_fd_sc_hd__or2_1
XANTENNA__10213__B _10934_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08750__B1 _08676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09768_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__nor2_1
XFILLER_46_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09290__A _09290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08865_/B vssd1 vssd1 vccd1 vccd1 _08840_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09769_/A _09764_/A _09810_/B _09769_/B vssd1 vssd1 vccd1 vccd1 _09844_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10612_ _10851_/CLK _10612_/D vssd1 vssd1 vccd1 vccd1 _10612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10543_ _10651_/CLK _10543_/D vssd1 vssd1 vccd1 vccd1 _10543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10474_ _10495_/A _10474_/B vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__nand2_2
XFILLER_6_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08033__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06044__B2 _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_6_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07713__A _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09049__A1 _10934_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05380_ _05380_/A _05380_/B vssd1 vssd1 vccd1 vccd1 _05380_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07050_ _07048_/A _07048_/B _07464_/A vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__a21oi_1
X_06001_ _10528_/A _07849_/A _06120_/S vssd1 vssd1 vccd1 vccd1 _06002_/B sky130_fd_sc_hd__mux2_1
XFILLER_114_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07952_ _07955_/A _07952_/B vssd1 vssd1 vccd1 vccd1 _07953_/A sky130_fd_sc_hd__or2_1
XFILLER_102_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07883_ _10602_/Q _07870_/X _07874_/X _07882_/Y vssd1 vssd1 vccd1 vccd1 _07884_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_06903_ _06903_/A _06903_/B vssd1 vssd1 vccd1 vccd1 _06921_/B sky130_fd_sc_hd__xor2_2
XFILLER_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06834_ _06834_/A _06834_/B vssd1 vssd1 vccd1 vccd1 _06835_/B sky130_fd_sc_hd__nor2_1
X_09622_ _09623_/A _09623_/B _09623_/C vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__o21ai_1
XFILLER_55_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09553_ _09553_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09554_/C sky130_fd_sc_hd__xnor2_1
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08504_ _10787_/Q _08496_/X _08502_/X hold23/A vssd1 vssd1 vccd1 vccd1 _10750_/D
+ sky130_fd_sc_hd__a22o_1
X_06765_ _06834_/A _06765_/B vssd1 vssd1 vccd1 vccd1 _06766_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05716_ _08196_/A _10555_/Q _05663_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _05717_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06239__A _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09484_ _10967_/Q _09579_/A vssd1 vssd1 vccd1 vccd1 _09486_/A sky130_fd_sc_hd__and2_1
X_06696_ _06693_/A _06693_/B _06691_/A vssd1 vssd1 vccd1 vccd1 _06697_/B sky130_fd_sc_hd__o21a_1
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05647_ _05912_/B _05539_/Y _05540_/X _05646_/X vssd1 vssd1 vccd1 vccd1 _05647_/X
+ sky130_fd_sc_hd__a31o_1
X_08435_ _10767_/Q _10730_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08366_ _08531_/A vssd1 vssd1 vccd1 vccd1 _08419_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05578_ _08315_/B vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__clkbuf_2
X_07317_ _07317_/A _07317_/B vssd1 vssd1 vccd1 vccd1 _07341_/A sky130_fd_sc_hd__or2_1
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08297_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07248_ _07248_/A _07382_/A vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__and2_1
XFILLER_133_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07179_ _07188_/B vssd1 vssd1 vccd1 vccd1 _07587_/B sky130_fd_sc_hd__buf_2
XFILLER_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10190_ _10947_/Q _10931_/Q vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__or2b_1
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08420__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10666_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10669_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput27 io_wbs_m2s_data[1] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_6
Xinput16 io_wbs_m2s_data[0] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_4
XFILLER_128_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10526_ _10526_/A _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10526_/X sky130_fd_sc_hd__or3_1
Xinput49 io_wbs_m2s_stb vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_2
Xinput38 io_wbs_m2s_data[2] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_4
X_10457_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10457_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07708__A _07708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10388_ _10365_/X _10716_/Q _10386_/X _10387_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10935_/D sky130_fd_sc_hd__o221a_1
XANTENNA__07765__A1 _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06550_ _10971_/Q _06550_/B _06550_/C vssd1 vssd1 vccd1 vccd1 _06587_/B sky130_fd_sc_hd__and3_1
X_05501_ _05369_/Y _05497_/X _05495_/X _05460_/C vssd1 vssd1 vccd1 vccd1 _10554_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_06481_ _06480_/B _06480_/C _06480_/A vssd1 vssd1 vccd1 vccd1 _06657_/A sky130_fd_sc_hd__o21a_1
X_08220_ _08216_/X _08224_/C _08067_/X vssd1 vssd1 vccd1 vccd1 _08220_/Y sky130_fd_sc_hd__o21ai_1
X_05432_ _10637_/Q vssd1 vssd1 vccd1 vccd1 _07893_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08274__A input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08151_ _08160_/B _08151_/B vssd1 vssd1 vccd1 vccd1 _08151_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08245__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05363_ _05363_/A _05363_/B vssd1 vssd1 vccd1 vccd1 _05363_/X sky130_fd_sc_hd__and2_1
X_08082_ _08082_/A _08082_/B _08082_/C _08082_/D vssd1 vssd1 vccd1 vccd1 _08095_/B
+ sky130_fd_sc_hd__and4_1
X_05294_ _05388_/A _05392_/A vssd1 vssd1 vccd1 vccd1 _05389_/A sky130_fd_sc_hd__and2_1
X_07102_ _07102_/A vssd1 vssd1 vccd1 vccd1 _07382_/A sky130_fd_sc_hd__clkbuf_2
X_07033_ _07044_/A _07421_/A _07417_/A vssd1 vssd1 vccd1 vccd1 _07034_/B sky130_fd_sc_hd__and3_1
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08984_ _09035_/B vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07935_ _10432_/B _07935_/B vssd1 vssd1 vccd1 vccd1 _07950_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05519__B1 _05474_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ _10880_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09605_ _09549_/A _09549_/B _09678_/A vssd1 vssd1 vccd1 vccd1 _09608_/A sky130_fd_sc_hd__o21ai_1
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06817_ _07670_/A _06817_/B vssd1 vssd1 vccd1 vccd1 _06818_/B sky130_fd_sc_hd__nand2_1
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07797_ _07797_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__xnor2_1
X_09536_ _10969_/Q _09536_/B vssd1 vssd1 vccd1 vccd1 _09638_/C sky130_fd_sc_hd__nand2_1
XFILLER_43_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06748_ _06758_/B _06774_/B vssd1 vssd1 vccd1 vccd1 _06748_/X sky130_fd_sc_hd__and2_2
X_09467_ _09516_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__or2_1
X_08418_ _10394_/B _08418_/B vssd1 vssd1 vccd1 vccd1 _08419_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06679_ _06678_/A _06678_/C _06678_/B vssd1 vssd1 vccd1 vccd1 _06945_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09398_ _09433_/A _09398_/B vssd1 vssd1 vccd1 vccd1 _09399_/B sky130_fd_sc_hd__xnor2_2
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08349_ _08351_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08349_/X sky130_fd_sc_hd__and2_1
XFILLER_7_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _10310_/X _10309_/A _10329_/S vssd1 vssd1 vccd1 vccd1 _10312_/B sky130_fd_sc_hd__mux2_1
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10242_ _10937_/Q _10953_/Q vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__or2b_1
XFILLER_120_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10173_ _07056_/A _10167_/X _10170_/X _10886_/Q vssd1 vssd1 vccd1 vccd1 _10886_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input38_A io_wbs_m2s_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10282__A2 _10253_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07986__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10509_ _05958_/X _10496_/X _10508_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10975_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07438__A _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06061__B _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05981_ _10533_/A vssd1 vssd1 vccd1 vccd1 _05982_/A sky130_fd_sc_hd__buf_4
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _07720_/A _07720_/B vssd1 vssd1 vccd1 vccd1 _07745_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07651_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07653_/B sky130_fd_sc_hd__xnor2_2
XFILLER_92_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06602_ _06602_/A _06602_/B vssd1 vssd1 vccd1 vccd1 _06616_/B sky130_fd_sc_hd__or2_2
X_07582_ _07583_/B _07582_/B vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__and2b_1
XFILLER_80_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09321_ _09396_/B _09396_/C vssd1 vssd1 vccd1 vccd1 _09323_/B sky130_fd_sc_hd__xor2_4
X_06533_ _06533_/A _06538_/B vssd1 vssd1 vccd1 vccd1 _06534_/B sky130_fd_sc_hd__xnor2_1
X_09252_ _08289_/A _09251_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10273__A2 _10115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06464_ _06465_/A _06465_/B vssd1 vssd1 vccd1 vccd1 _06480_/C sky130_fd_sc_hd__and2_1
XFILLER_21_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08203_ _08200_/X _08203_/B vssd1 vssd1 vccd1 vccd1 _08204_/A sky130_fd_sc_hd__and2b_1
X_05415_ _05462_/C _05393_/B _05414_/X vssd1 vssd1 vccd1 vccd1 _05415_/X sky130_fd_sc_hd__o21a_1
X_09183_ _09112_/A _09178_/Y _09182_/X vssd1 vssd1 vccd1 vccd1 _09184_/B sky130_fd_sc_hd__a21oi_1
X_06395_ _06874_/A _06395_/B vssd1 vssd1 vccd1 vccd1 _06396_/A sky130_fd_sc_hd__xnor2_1
X_08134_ _06168_/X _08047_/X _08052_/X _08132_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08134_/X sky130_fd_sc_hd__o221a_1
X_05346_ _05347_/B _05346_/B vssd1 vssd1 vccd1 vccd1 _05346_/X sky130_fd_sc_hd__and2_1
XFILLER_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08065_ _10580_/Q _08065_/B vssd1 vssd1 vccd1 vccd1 _08113_/A sky130_fd_sc_hd__and2_2
X_05277_ _05291_/A _05818_/B vssd1 vssd1 vccd1 vccd1 _05277_/Y sky130_fd_sc_hd__nand2_1
XFILLER_122_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07016_ _07235_/C vssd1 vssd1 vccd1 vccd1 _07186_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08967_ _08962_/Y _10495_/B _08966_/Y vssd1 vssd1 vccd1 vccd1 _08967_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08154__A1 input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07918_ _09154_/A vssd1 vssd1 vccd1 vccd1 _08284_/A sky130_fd_sc_hd__clkbuf_4
X_08898_ _08889_/A _08892_/Y _08896_/X _08688_/A vssd1 vssd1 vccd1 vccd1 _08898_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10502__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08154__B2 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07849_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07849_/X sky130_fd_sc_hd__buf_4
XFILLER_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10859__D _10859_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10860_ _10865_/CLK _10860_/D vssd1 vssd1 vccd1 vccd1 _10860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07811__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09519_ _09562_/B _09562_/C _09562_/A vssd1 vssd1 vccd1 vccd1 _09520_/C sky130_fd_sc_hd__a21oi_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _10791_/CLK _10791_/D vssd1 vssd1 vccd1 vccd1 _10791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05985__B input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06162__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10225_ _10225_/A _10225_/B vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10156_ _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _10157_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10412__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _10087_/A _10087_/B vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__xnor2_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__05506__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06180_ hold3/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__or3_1
XANTENNA__10204__B_N _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08821_ input24/X _08819_/X _08820_/X _10816_/Q _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08821_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09377__B_N _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08748_/X _08815_/B _08759_/A vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__a21oi_1
X_05964_ input7/X input4/X input9/X vssd1 vssd1 vccd1 vccd1 _09142_/C sky130_fd_sc_hd__or3_4
XFILLER_57_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08683_ _08778_/A _08683_/B _08692_/B vssd1 vssd1 vccd1 vccd1 _08683_/X sky130_fd_sc_hd__and3_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07703_ _09824_/A _09824_/B _07702_/X vssd1 vssd1 vccd1 vccd1 _09899_/B sky130_fd_sc_hd__a21o_1
X_05895_ _05895_/A _05895_/B vssd1 vssd1 vccd1 vccd1 _05895_/X sky130_fd_sc_hd__and2_1
X_07634_ _07670_/A vssd1 vssd1 vccd1 vccd1 _07635_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07565_ _07563_/X _07565_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__and2b_1
XANTENNA__06247__A _07977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07534_/C sky130_fd_sc_hd__nor2_1
X_06516_ _06517_/A _06517_/B _06680_/A vssd1 vssd1 vccd1 vccd1 _06521_/B sky130_fd_sc_hd__and3_1
X_09304_ _09304_/A _10882_/Q vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ _09259_/A _09235_/B vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__and2_1
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06447_ _06472_/A _06472_/B _06675_/A _06675_/B vssd1 vssd1 vccd1 vccd1 _06448_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_09166_ _09114_/X _09165_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__o21a_1
X_06378_ _06872_/A _06409_/C vssd1 vssd1 vccd1 vccd1 _06393_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05329_ _05329_/A _05329_/B vssd1 vssd1 vccd1 vccd1 _05329_/X sky130_fd_sc_hd__and2_1
X_08117_ _08117_/A _08117_/B vssd1 vssd1 vccd1 vccd1 _08117_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09097_ _10129_/A vssd1 vssd1 vccd1 vccd1 _10493_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08048_ _08048_/A vssd1 vssd1 vccd1 vccd1 _09124_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10010_ _10081_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09999_ _09999_/A vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__inv_2
XFILLER_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05326__A _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10912_ _10960_/CLK _10912_/D vssd1 vssd1 vccd1 vccd1 _10912_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10843_ _10848_/CLK _10843_/D vssd1 vssd1 vccd1 vccd1 _10843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10774_ _10833_/CLK _10774_/D vssd1 vssd1 vccd1 vccd1 _10774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05996__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08063__B1 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10208_ _10226_/A _10206_/Y _10279_/S vssd1 vssd1 vccd1 vccd1 _10208_/X sky130_fd_sc_hd__mux2_1
X_10139_ _10138_/B _10138_/Y _10139_/S vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__mux2_1
XANTENNA__07435__B _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09866__B2 _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05680_ _05803_/A vssd1 vssd1 vccd1 vccd1 _08317_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07350_ _07461_/B _07350_/B vssd1 vssd1 vccd1 vccd1 _07470_/A sky130_fd_sc_hd__nor2_1
X_06301_ _10921_/Q _10904_/Q vssd1 vssd1 vccd1 vccd1 _06386_/A sky130_fd_sc_hd__xnor2_2
X_09020_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _09020_/X sky130_fd_sc_hd__or2_1
X_07281_ _07282_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _07366_/B sky130_fd_sc_hd__nand2_1
X_06232_ input30/X _06225_/X _06231_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10606_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06163_ _10535_/A vssd1 vssd1 vccd1 vccd1 _06163_/X sky130_fd_sc_hd__buf_4
XFILLER_132_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06094_ _10681_/Q _10680_/Q vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__or2_2
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06080__A2 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09922_ _10065_/D _09922_/B vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__xnor2_2
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09853_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09853_/Y sky130_fd_sc_hd__nand2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08804_ _08804_/A _08804_/B _08804_/C _08804_/D vssd1 vssd1 vccd1 vccd1 _08804_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09784_ _09784_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__or2_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08735_ _10805_/Q _08815_/B _08726_/Y vssd1 vssd1 vccd1 vccd1 _08736_/B sky130_fd_sc_hd__a21bo_1
X_06996_ _10907_/Q vssd1 vssd1 vccd1 vccd1 _07013_/A sky130_fd_sc_hd__buf_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05947_ _08339_/A _05947_/B vssd1 vssd1 vccd1 vccd1 _05947_/X sky130_fd_sc_hd__or2_1
XFILLER_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09857__A1 _09930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__B2 _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05878_ _07991_/A _05878_/B vssd1 vssd1 vccd1 vccd1 _05878_/Y sky130_fd_sc_hd__xnor2_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _10800_/Q _08678_/A vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__nand2_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _08661_/A _08597_/B vssd1 vssd1 vccd1 vccd1 _08617_/B sky130_fd_sc_hd__and2_1
XFILLER_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07617_ _07622_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07618_/A sky130_fd_sc_hd__nand2_1
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07548_ _07549_/A _07549_/B vssd1 vssd1 vccd1 vccd1 _07743_/B sky130_fd_sc_hd__nor2_1
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07479_ _07497_/A _07497_/B vssd1 vssd1 vccd1 vccd1 _07504_/B sky130_fd_sc_hd__and2_1
XFILLER_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09218_ _09218_/A vssd1 vssd1 vccd1 vccd1 _10851_/D sky130_fd_sc_hd__clkbuf_1
X_10490_ _05982_/A _10489_/B _10489_/Y _10485_/X vssd1 vssd1 vccd1 vccd1 _10968_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08045__B1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09149_ _05461_/B _09136_/X _09148_/X _08160_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09149_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_2_2_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input20_A io_wbs_m2s_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10826_ _10826_/CLK _10826_/D vssd1 vssd1 vccd1 vccd1 _10826_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_2_clock_A _10981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10757_ _10798_/CLK _10757_/D vssd1 vssd1 vccd1 vccd1 _10757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10688_ _10841_/CLK _10688_/D vssd1 vssd1 vccd1 vccd1 _10688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06062__A2 _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06850_ _06850_/A _06288_/X vssd1 vssd1 vccd1 vccd1 _06852_/A sky130_fd_sc_hd__or2b_1
X_05801_ _05717_/X _05742_/C _05796_/X _05800_/X _05702_/X vssd1 vssd1 vccd1 vccd1
+ _05802_/B sky130_fd_sc_hd__o32a_1
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06781_ _06781_/A _06781_/B vssd1 vssd1 vccd1 vccd1 _06782_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05732_ _05794_/A _05732_/B _05732_/C _05732_/D vssd1 vssd1 vccd1 vccd1 _05788_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08520_ _10798_/Q _08514_/X _08517_/X _10761_/Q vssd1 vssd1 vccd1 vccd1 _10761_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05663_ _05663_/A _05663_/B vssd1 vssd1 vccd1 vccd1 _05664_/B sky130_fd_sc_hd__and2_1
X_08451_ _08451_/A vssd1 vssd1 vccd1 vccd1 _10734_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07181__A _07229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07402_ _07402_/A _07402_/B vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__xnor2_1
X_05594_ _10701_/Q vssd1 vssd1 vccd1 vccd1 _08277_/B sky130_fd_sc_hd__clkbuf_2
X_08382_ _08367_/X _10734_/Q _08380_/X _08381_/X vssd1 vssd1 vccd1 vccd1 _10716_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07333_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07522_/A sky130_fd_sc_hd__xnor2_1
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07264_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07266_/A sky130_fd_sc_hd__xor2_1
X_06215_ _06206_/X _06207_/X _06214_/X _06200_/X vssd1 vssd1 vccd1 vccd1 _10599_/D
+ sky130_fd_sc_hd__o211a_1
X_09003_ _09610_/A vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07195_ _07195_/A _07334_/A vssd1 vssd1 vccd1 vccd1 _07196_/B sky130_fd_sc_hd__or2b_1
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06146_ _06143_/X _06131_/X _06145_/Y _06137_/X vssd1 vssd1 vccd1 vccd1 _10586_/D
+ sky130_fd_sc_hd__o211a_1
X_06077_ _08355_/A _08352_/A _08029_/A _10709_/Q _06076_/X vssd1 vssd1 vccd1 vccd1
+ _06082_/B sky130_fd_sc_hd__a221o_1
XFILLER_132_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09905_ _09971_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09836_ _09837_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__nand2_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _09767_/A _09767_/B vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__and2_1
X_06979_ _10900_/Q vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08856_/B vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10510__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09698_ _09767_/A _09767_/B vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__xnor2_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _08649_/A _08649_/B _08649_/C vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__and3_1
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _10851_/CLK _10611_/D vssd1 vssd1 vccd1 vccd1 _10611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10542_ _10682_/CLK _10542_/D vssd1 vssd1 vccd1 vccd1 _10542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10473_ _06206_/X _10459_/A _10472_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10962_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06044__A2 _10671_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10809_ _10813_/CLK _10809_/D vssd1 vssd1 vccd1 vccd1 _10809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06000_ _10577_/Q vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__buf_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09375__B _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08980__A1 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ input42/X _05905_/A _07983_/A vssd1 vssd1 vccd1 vccd1 _07952_/B sky130_fd_sc_hd__mux2_1
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06902_ _06902_/A _06902_/B vssd1 vssd1 vccd1 vccd1 _06921_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08193__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07882_ _07882_/A vssd1 vssd1 vccd1 vccd1 _07882_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06833_ _06833_/A _06833_/B vssd1 vssd1 vccd1 vccd1 _06835_/A sky130_fd_sc_hd__nand2_1
X_09621_ _09621_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09623_/C sky130_fd_sc_hd__xor2_1
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06764_ _06834_/A _06765_/B vssd1 vssd1 vccd1 vccd1 _06766_/A sky130_fd_sc_hd__and2_1
X_09552_ _09610_/A _09552_/B _09599_/B vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__and3_1
X_05715_ _08139_/A _10549_/Q _05702_/X _05708_/Y _05714_/X vssd1 vssd1 vccd1 vccd1
+ _05717_/C sky130_fd_sc_hd__a2111o_1
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08503_ _10786_/Q _08496_/X _08502_/X hold27/A vssd1 vssd1 vccd1 vccd1 _10749_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_91_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06695_ _06695_/A _06695_/B vssd1 vssd1 vccd1 vccd1 _06698_/B sky130_fd_sc_hd__xor2_2
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09483_ _09483_/A _09483_/B vssd1 vssd1 vccd1 vccd1 _09527_/A sky130_fd_sc_hd__xor2_2
X_05646_ _10681_/Q _05644_/Y _05541_/X vssd1 vssd1 vccd1 vccd1 _05646_/X sky130_fd_sc_hd__a21bo_1
X_08434_ _08476_/S vssd1 vssd1 vccd1 vccd1 _08486_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05577_ _10705_/Q vssd1 vssd1 vccd1 vccd1 _08315_/B sky130_fd_sc_hd__clkbuf_2
X_08365_ _10729_/Q vssd1 vssd1 vccd1 vccd1 _08531_/A sky130_fd_sc_hd__inv_2
XANTENNA__08799__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _07309_/A _07152_/B _07322_/A vssd1 vssd1 vccd1 vccd1 _07317_/B sky130_fd_sc_hd__a21oi_1
XFILLER_20_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08296_ _08297_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08296_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07247_ _07269_/A _07247_/B vssd1 vssd1 vccd1 vccd1 _07513_/A sky130_fd_sc_hd__nand2_1
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07178_ _07178_/A vssd1 vssd1 vccd1 vccd1 _07398_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06129_ _10432_/B _06129_/B vssd1 vssd1 vccd1 vccd1 _06149_/A sky130_fd_sc_hd__nand2_2
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09819_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09820_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10530__A1 _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput17 io_wbs_m2s_data[10] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput28 io_wbs_m2s_data[20] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_28_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_1_0_clock _10985_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clock/X sky130_fd_sc_hd__clkbuf_16
Xinput39 io_wbs_m2s_data[30] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_4
X_10525_ _07442_/X _10522_/X _10524_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10980_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08380__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ _10956_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10456_/X sky130_fd_sc_hd__or2_1
XANTENNA__10349__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _10935_/Q _10379_/B _10376_/X vssd1 vssd1 vccd1 vccd1 _10387_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__05776__B2 _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10521__A1 _06124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05500_ _05371_/Y _05497_/X _05495_/X _05460_/D vssd1 vssd1 vccd1 vccd1 _10553_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06480_ _06480_/A _06480_/B _06480_/C vssd1 vssd1 vccd1 vccd1 _06657_/B sky130_fd_sc_hd__nor3_1
X_05431_ _07889_/A _05346_/X _05348_/X _10637_/Q _05430_/X vssd1 vssd1 vccd1 vccd1
+ _05431_/X sky130_fd_sc_hd__a221o_1
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__nand2_1
XFILLER_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06075__A _10677_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05362_ _10663_/Q _05362_/B vssd1 vssd1 vccd1 vccd1 _05363_/B sky130_fd_sc_hd__nand2_1
X_07101_ _10986_/Q _07327_/A vssd1 vssd1 vccd1 vccd1 _07384_/A sky130_fd_sc_hd__nand2_1
X_08081_ _08075_/A _08059_/A _08082_/D _05733_/X vssd1 vssd1 vccd1 vccd1 _08081_/X
+ sky130_fd_sc_hd__a31o_1
X_05293_ _10653_/Q _05391_/B vssd1 vssd1 vccd1 vccd1 _05392_/A sky130_fd_sc_hd__nor2_1
X_07032_ _07042_/A _07042_/B vssd1 vssd1 vccd1 vccd1 _07043_/A sky130_fd_sc_hd__and2_1
XFILLER_115_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10970__D _10970_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06803__A _07682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08953__A1 _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08983_ _06019_/A _08972_/X _08974_/X _08982_/X vssd1 vssd1 vccd1 vccd1 _08983_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07934_ _08995_/A vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07865_ _08557_/A vssd1 vssd1 vccd1 vccd1 _07865_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07634__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08159__B1_N _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _09655_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09613_/B sky130_fd_sc_hd__and2_1
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10060__A _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06816_ _06856_/A vssd1 vssd1 vccd1 vccd1 _10502_/A sky130_fd_sc_hd__buf_2
X_07796_ _07796_/A _07796_/B _07795_/X vssd1 vssd1 vccd1 vccd1 _07797_/B sky130_fd_sc_hd__or3b_1
X_09535_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__xnor2_1
X_06747_ _06785_/A _06747_/B _06776_/A vssd1 vssd1 vccd1 vccd1 _06763_/A sky130_fd_sc_hd__and3_1
X_06678_ _06678_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__and3_1
XFILLER_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09552_/B _09466_/B vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__and2_1
X_05629_ _10548_/Q _05629_/B vssd1 vssd1 vccd1 vccd1 _05630_/B sky130_fd_sc_hd__nand2_1
X_08417_ _09037_/A vssd1 vssd1 vccd1 vccd1 _08418_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ _10131_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09398_/B sky130_fd_sc_hd__nand2_1
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08348_ input39/X vssd1 vssd1 vccd1 vccd1 _08348_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08279_ _08278_/A _08278_/B _08255_/A vssd1 vssd1 vccd1 vccd1 _08279_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08912__B _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07809__A hold16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _10292_/A _10289_/A _10298_/B _10309_/Y vssd1 vssd1 vccd1 vccd1 _10310_/X
+ sky130_fd_sc_hd__a31o_1
X_10241_ _07066_/A _10192_/X _10240_/Y vssd1 vssd1 vccd1 vccd1 _10903_/D sky130_fd_sc_hd__a21o_1
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _07113_/A _10167_/X _10170_/X _10885_/Q vssd1 vssd1 vccd1 vccd1 _10885_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10503__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05999__A input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10508_ _10508_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10508_/X sky130_fd_sc_hd__or2_1
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10439_ _10949_/Q _10431_/X _10438_/X vssd1 vssd1 vccd1 vccd1 _10949_/D sky130_fd_sc_hd__a21o_1
XFILLER_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05980_ input43/X vssd1 vssd1 vccd1 vccd1 _10533_/A sky130_fd_sc_hd__buf_4
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07650_ _07659_/A _07658_/B _07635_/A vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__o21a_1
XFILLER_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06601_ _06775_/A _06409_/B _06522_/C vssd1 vssd1 vccd1 vccd1 _06602_/B sky130_fd_sc_hd__a21oi_1
X_07581_ _07581_/A _07581_/B vssd1 vssd1 vccd1 vccd1 _07582_/B sky130_fd_sc_hd__xor2_1
X_09320_ _10069_/A _09744_/A vssd1 vssd1 vccd1 vccd1 _09396_/C sky130_fd_sc_hd__nand2_2
XFILLER_18_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06532_ _06532_/A _06532_/B vssd1 vssd1 vccd1 vccd1 _06538_/B sky130_fd_sc_hd__xor2_1
X_09251_ _08287_/A _07900_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09251_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08202_ input21/X _08123_/X _08124_/X _05877_/X _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08203_/B sky130_fd_sc_hd__o221a_1
XANTENNA__10965__D _10965_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06463_ _06479_/A _06479_/B vssd1 vssd1 vccd1 vccd1 _06465_/B sky130_fd_sc_hd__xor2_1
XFILLER_119_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05414_ _10620_/Q _05487_/A _05413_/X vssd1 vssd1 vccd1 vccd1 _05414_/X sky130_fd_sc_hd__a21o_1
X_09182_ _10812_/Q _09168_/X _09079_/X _10725_/Q _09181_/X vssd1 vssd1 vccd1 vccd1
+ _09182_/X sky130_fd_sc_hd__a221o_1
X_06394_ _06394_/A _06394_/B vssd1 vssd1 vccd1 vccd1 _06395_/B sky130_fd_sc_hd__xnor2_1
X_08133_ _08038_/X _08074_/X _08132_/Y _08044_/X _06050_/X vssd1 vssd1 vccd1 vccd1
+ _08133_/X sky130_fd_sc_hd__a32o_1
X_05345_ _10667_/Q _05350_/B _10668_/Q vssd1 vssd1 vccd1 vccd1 _05346_/B sky130_fd_sc_hd__o21ai_1
X_08064_ _05813_/A _08058_/X _08063_/X vssd1 vssd1 vccd1 vccd1 _08064_/X sky130_fd_sc_hd__o21ba_1
XFILLER_119_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05276_ _10576_/Q vssd1 vssd1 vccd1 vccd1 _05818_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07015_ _10982_/Q vssd1 vssd1 vccd1 vccd1 _07235_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08966_ _07780_/C _08964_/A _08965_/Y vssd1 vssd1 vccd1 vccd1 _08966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_44_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10673_/CLK sky130_fd_sc_hd__clkbuf_16
X_07917_ _08462_/A vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__buf_4
X_08897_ _08889_/A _08892_/Y _08896_/X vssd1 vssd1 vccd1 vccd1 _08897_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07848_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07848_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07779_ _07779_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__nor2_1
X_09518_ _09562_/A _09562_/B _09562_/C vssd1 vssd1 vccd1 vccd1 _09520_/B sky130_fd_sc_hd__and3_1
XFILLER_25_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08311__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _10790_/CLK _10790_/D vssd1 vssd1 vccd1 vccd1 _10790_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_59_clock clkbuf_opt_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _10862_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ _09449_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__nand2_1
XFILLER_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07539__A _07539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05979__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input50_A io_wbs_m2s_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10224_ _10224_/A _10935_/Q vssd1 vssd1 vccd1 vccd1 _10225_/B sky130_fd_sc_hd__and2_1
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10156_/B sky130_fd_sc_hd__xnor2_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_10086_ _09998_/A _10138_/B _09997_/B _10017_/A vssd1 vssd1 vccd1 vccd1 _10087_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08908__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08820_ _08820_/A vssd1 vssd1 vccd1 vccd1 _08820_/X sky130_fd_sc_hd__clkbuf_2
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08751_ _10808_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08759_/B sky130_fd_sc_hd__xor2_1
X_05963_ _07967_/A vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05894_ _07974_/A _05900_/A _06039_/A vssd1 vssd1 vccd1 vccd1 _05895_/B sky130_fd_sc_hd__o21ai_1
X_08682_ _08669_/B _08670_/C _08679_/X _08680_/Y vssd1 vssd1 vccd1 vccd1 _08692_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_66_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07702_ _07621_/A _07702_/B vssd1 vssd1 vccd1 vccd1 _07702_/X sky130_fd_sc_hd__and2b_1
XFILLER_93_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07633_ _07633_/A _07633_/B vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__xor2_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07564_ _07563_/A _07727_/B _07563_/C vssd1 vssd1 vccd1 vccd1 _07565_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07631__B _07698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07495_ _07495_/A _07495_/B vssd1 vssd1 vccd1 vccd1 _07506_/B sky130_fd_sc_hd__xnor2_1
X_06515_ _06758_/B _06515_/B vssd1 vssd1 vccd1 vccd1 _06680_/A sky130_fd_sc_hd__nand2_1
X_09303_ _09303_/A _09303_/B vssd1 vssd1 vccd1 vccd1 _09310_/C sky130_fd_sc_hd__nor2_1
X_09234_ _08847_/X _09210_/X _09212_/X _09233_/X _09203_/X vssd1 vssd1 vccd1 vccd1
+ _09235_/B sky130_fd_sc_hd__a32o_1
X_06446_ _06461_/B _06459_/B vssd1 vssd1 vccd1 vccd1 _06675_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ _10943_/Q _09008_/X _09164_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09165_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_08116_ _08117_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _08116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06377_ _06436_/A _06513_/D vssd1 vssd1 vccd1 vccd1 _06409_/C sky130_fd_sc_hd__and2_1
X_05328_ _10675_/Q _05834_/A vssd1 vssd1 vccd1 vccd1 _05329_/B sky130_fd_sc_hd__nand2_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09096_ _09977_/A vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__06083__B1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08047_ _08248_/A vssd1 vssd1 vccd1 vccd1 _08047_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_107_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09998_ _09998_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10513__A _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08949_ input10/X vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__inv_2
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06138__A1 _06124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10911_ _10960_/CLK _10911_/D vssd1 vssd1 vccd1 vccd1 _10911_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09088__A0 _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _10842_/CLK _10842_/D vssd1 vssd1 vccd1 vccd1 _10842_/Q sky130_fd_sc_hd__dfxtp_1
X_10773_ _10833_/CLK _10773_/D vssd1 vssd1 vccd1 vccd1 _10773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06074__B1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09012__A0 _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10207_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10279_/S sky130_fd_sc_hd__buf_2
XANTENNA__05517__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10138_ _10487_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10138_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10069_ _10069_/A _10069_/B _10140_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__and3_1
XFILLER_48_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07732__A _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09659__A _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06300_ _06262_/A _06304_/A _06304_/B vssd1 vssd1 vccd1 vccd1 _06303_/A sky130_fd_sc_hd__a21bo_1
X_07280_ _07280_/A _07280_/B _07280_/C _07289_/A vssd1 vssd1 vccd1 vccd1 _07282_/B
+ sky130_fd_sc_hd__or4_1
X_06231_ _10606_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06231_/X sky130_fd_sc_hd__or2_1
XANTENNA__08563__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08282__B _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_76_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06162_ input44/X vssd1 vssd1 vccd1 vccd1 _10535_/A sky130_fd_sc_hd__buf_4
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06093_ _08236_/A vssd1 vssd1 vccd1 vccd1 _08062_/A sky130_fd_sc_hd__buf_2
XFILLER_117_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _09921_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _10065_/D sky130_fd_sc_hd__nor2_1
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09852_ _09852_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__nor2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07626__B _07700_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08803_ _08777_/A _08803_/B _08803_/C _08803_/D vssd1 vssd1 vccd1 vccd1 _08804_/D
+ sky130_fd_sc_hd__and4b_1
XANTENNA__08762__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ _09713_/B _09718_/Y _09781_/Y _09780_/X vssd1 vssd1 vccd1 vccd1 _09784_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08734_ _08928_/B vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__buf_2
XFILLER_65_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06995_ _09344_/B vssd1 vssd1 vccd1 vccd1 _07008_/A sky130_fd_sc_hd__buf_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05946_ _08339_/A _05947_/B _05836_/X _08332_/A _05945_/X vssd1 vssd1 vccd1 vccd1
+ _05946_/X sky130_fd_sc_hd__a221o_1
XFILLER_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05877_ _05877_/A vssd1 vssd1 vccd1 vccd1 _05877_/X sky130_fd_sc_hd__buf_2
X_08665_ _10832_/Q _10764_/Q vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__xnor2_2
XFILLER_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06258__A _07849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ _08623_/C vssd1 vssd1 vccd1 vccd1 _08597_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07616_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _07616_/X sky130_fd_sc_hd__or2_1
XFILLER_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07547_ _07743_/A _07547_/B vssd1 vssd1 vccd1 vccd1 _07549_/B sky130_fd_sc_hd__or2_1
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09349__A_N _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07478_ _07477_/A _07477_/B _07480_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07497_/B
+ sky130_fd_sc_hd__o2bb2ai_1
X_09217_ _09228_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09218_/A sky130_fd_sc_hd__and2_1
XANTENNA__10508__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06429_ _06630_/A _06407_/B _06425_/Y _06656_/A vssd1 vssd1 vccd1 vccd1 _06430_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__08045__A1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09148_ _09148_/A vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09079_ _09079_/A vssd1 vssd1 vccd1 vccd1 _09079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input13_A io_wbs_m2s_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06168__A _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10825_ _10826_/CLK _10825_/D vssd1 vssd1 vccd1 vccd1 _10825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10756_ _10791_/CLK _10756_/D vssd1 vssd1 vccd1 vccd1 _10756_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09481__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10687_ _10841_/CLK _10687_/D vssd1 vssd1 vccd1 vccd1 _10687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07727__A _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05800_ _05717_/D _05799_/X _05708_/B vssd1 vssd1 vccd1 vccd1 _05800_/X sky130_fd_sc_hd__o21a_1
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06780_ _06781_/A _06781_/B vssd1 vssd1 vccd1 vccd1 _06782_/A sky130_fd_sc_hd__and2_1
X_05731_ _05728_/X _05729_/Y _05547_/A _08093_/A vssd1 vssd1 vccd1 vccd1 _05732_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05662_ _08169_/A _05617_/X _05619_/X _05885_/A _05661_/X vssd1 vssd1 vccd1 vccd1
+ _05662_/X sky130_fd_sc_hd__a221o_1
X_08450_ _08460_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08451_/A sky130_fd_sc_hd__or2_1
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08381_ _08381_/A hold23/X vssd1 vssd1 vccd1 vccd1 _08381_/X sky130_fd_sc_hd__or2_1
XFILLER_51_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07401_ _07070_/A _07359_/A _07398_/B _07562_/A vssd1 vssd1 vccd1 vccd1 _07402_/B
+ sky130_fd_sc_hd__o211a_1
X_05593_ _05593_/A _05593_/B vssd1 vssd1 vccd1 vccd1 _05593_/X sky130_fd_sc_hd__and2_1
X_07332_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07525_/A sky130_fd_sc_hd__or2b_1
X_07263_ _07334_/A _07195_/A _07262_/X vssd1 vssd1 vccd1 vccd1 _07268_/A sky130_fd_sc_hd__o21ai_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06214_ _10599_/Q _06223_/B vssd1 vssd1 vccd1 vccd1 _06214_/X sky130_fd_sc_hd__or2_1
X_09002_ _10964_/Q vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07194_ _07194_/A _07194_/B vssd1 vssd1 vccd1 vccd1 _07210_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06145_ _06145_/A _06145_/B vssd1 vssd1 vccd1 vccd1 _06145_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06076_ _05781_/Y _05844_/A _08256_/A _05751_/Y vssd1 vssd1 vccd1 vccd1 _06076_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09904_ _09904_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _09905_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09835_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__nor2_1
XANTENNA_input5_A io_wbs_m2s_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09766_ _09842_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__or2_1
X_06978_ _10902_/Q vssd1 vssd1 vccd1 vccd1 _07056_/A sky130_fd_sc_hd__buf_2
XFILLER_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05929_ _05877_/X _05878_/Y _05876_/X _08206_/A _05928_/X vssd1 vssd1 vccd1 vccd1
+ _05929_/X sky130_fd_sc_hd__a221o_1
XFILLER_92_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08717_ _08801_/B vssd1 vssd1 vccd1 vccd1 _08856_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_73_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09697_ _09588_/A _09640_/A _09639_/B _09769_/B vssd1 vssd1 vccd1 vccd1 _09767_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _10797_/Q _08648_/B vssd1 vssd1 vccd1 vccd1 _08649_/C sky130_fd_sc_hd__nand2_1
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07710__B1 _07539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08579_ _10778_/Q _08578_/C _08578_/D _10779_/Q vssd1 vssd1 vccd1 vccd1 _08580_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _10851_/CLK _10610_/D vssd1 vssd1 vccd1 vccd1 _10610_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09299__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10541_ _10682_/CLK _10541_/D vssd1 vssd1 vccd1 vccd1 _10541_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08634__C _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09215__A0 _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06029__B1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ _10962_/Q _10472_/B vssd1 vssd1 vccd1 vccd1 _10472_/X sky130_fd_sc_hd__or2_1
XFILLER_123_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10808_ _10808_/CLK _10808_/D vssd1 vssd1 vccd1 vccd1 _10808_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10739_ _10836_/CLK _10739_/D vssd1 vssd1 vccd1 vccd1 _10739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07950_ _07950_/A vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__buf_2
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06901_ _10504_/A _07776_/B _06773_/C vssd1 vssd1 vccd1 vccd1 _06902_/B sky130_fd_sc_hd__a21oi_1
X_07881_ _07899_/A vssd1 vssd1 vccd1 vccd1 _07898_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06832_ _06832_/A _06794_/B vssd1 vssd1 vccd1 vccd1 _06833_/B sky130_fd_sc_hd__or2b_1
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10968__D _10968_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06763_ _06763_/A _06763_/B vssd1 vssd1 vccd1 vccd1 _06765_/B sky130_fd_sc_hd__xor2_1
X_09551_ _09867_/B _09760_/B vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05951__C1 _05950_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05714_ _05709_/Y _10551_/Q _10550_/Q _05711_/Y _05713_/X vssd1 vssd1 vccd1 vccd1
+ _05714_/X sky130_fd_sc_hd__a221o_1
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08502_ _10177_/A vssd1 vssd1 vccd1 vccd1 _08502_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09482_ _09479_/Y _09481_/X hold18/A _09406_/X vssd1 vssd1 vccd1 vccd1 _10870_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_06694_ _06915_/B _06942_/A _06915_/A vssd1 vssd1 vccd1 vccd1 _06916_/A sky130_fd_sc_hd__o21a_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05645_ _10681_/Q vssd1 vssd1 vccd1 vccd1 _08082_/C sky130_fd_sc_hd__clkbuf_2
X_08433_ _10218_/A _08661_/A _08432_/Y vssd1 vssd1 vccd1 vccd1 _08476_/S sky130_fd_sc_hd__a21oi_2
XFILLER_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08364_ _08364_/A vssd1 vssd1 vccd1 vccd1 _10711_/D sky130_fd_sc_hd__clkbuf_1
X_05576_ _05576_/A _05576_/B vssd1 vssd1 vccd1 vccd1 _05576_/X sky130_fd_sc_hd__and2_1
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09996__A1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09996__B2 _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _07347_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07470_/B sky130_fd_sc_hd__and2b_1
XFILLER_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08295_ _10704_/Q _10703_/Q _08295_/C vssd1 vssd1 vccd1 vccd1 _08315_/C sky130_fd_sc_hd__and3_1
XFILLER_109_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07246_ _07246_/A _07246_/B vssd1 vssd1 vccd1 vccd1 _07247_/B sky130_fd_sc_hd__or2_1
XFILLER_133_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07177_ _07200_/A _07200_/B _07176_/A vssd1 vssd1 vccd1 vccd1 _07183_/A sky130_fd_sc_hd__o21ai_2
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06128_ _09250_/A vssd1 vssd1 vccd1 vccd1 _06129_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__08420__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06059_ _08232_/A _08235_/A _07991_/A _05877_/X vssd1 vssd1 vccd1 vccd1 _06059_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_105_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09818_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__and2_1
XFILLER_74_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09749_ _09749_/A _09749_/B vssd1 vssd1 vccd1 vccd1 _09750_/B sky130_fd_sc_hd__and2_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07830__A _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08239__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 io_wbs_m2s_data[11] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_4
Xinput29 io_wbs_m2s_data[21] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08661__A _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10524_ input27/X _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__or3_1
XANTENNA__09757__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10455_ _06172_/X _10446_/X _10454_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10955_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _10531_/A _10394_/B _10394_/C vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__and3_1
XFILLER_2_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05430_ _07885_/A _05350_/X _05346_/X _10636_/Q _05429_/X vssd1 vssd1 vccd1 vccd1
+ _05430_/X sky130_fd_sc_hd__o221a_1
XFILLER_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05361_ _10631_/Q vssd1 vssd1 vccd1 vccd1 _07871_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06356__A _10978_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07100_ _07235_/B vssd1 vssd1 vccd1 vccd1 _07327_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08080_ _08098_/B _08079_/Y _06117_/D vssd1 vssd1 vccd1 vccd1 _08080_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05292_ _05277_/Y _05398_/A _05397_/B vssd1 vssd1 vccd1 vccd1 _05391_/B sky130_fd_sc_hd__a21o_1
XFILLER_9_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07031_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07042_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08982_ _05475_/X _08976_/X _08979_/X _08980_/Y _09078_/B vssd1 vssd1 vccd1 vccd1
+ _08982_/X sky130_fd_sc_hd__a221o_1
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07933_ _09124_/B _09092_/A vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__nor2_2
X_07864_ _07848_/X _05460_/C _07844_/X _07863_/Y vssd1 vssd1 vccd1 vccd1 _10629_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10341__A _10341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05519__A2 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06815_ _07780_/C _07766_/B vssd1 vssd1 vccd1 vccd1 _07779_/A sky130_fd_sc_hd__nand2_1
X_09603_ _09610_/B _09610_/C vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__and2_1
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07795_ _06719_/B _06718_/A _06718_/B _07791_/A vssd1 vssd1 vccd1 vccd1 _07795_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_71_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09534_ _10968_/Q _09579_/A _09534_/C vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__and3_1
X_06746_ _06746_/A _06746_/B vssd1 vssd1 vccd1 vccd1 _06776_/A sky130_fd_sc_hd__xnor2_2
XFILLER_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06677_ _06678_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06943_/B sky130_fd_sc_hd__nand3_1
X_09465_ _09552_/B _09466_/B vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__nor2_2
X_05628_ _10549_/Q _05630_/A vssd1 vssd1 vccd1 vccd1 _05628_/X sky130_fd_sc_hd__xor2_1
X_08416_ _08416_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__and2_1
XFILLER_52_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09396_ _09396_/A _09396_/B _09396_/C vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__nand3_1
X_08347_ _08347_/A vssd1 vssd1 vccd1 vccd1 _10709_/D sky130_fd_sc_hd__clkbuf_1
X_05559_ _10563_/Q _05596_/A vssd1 vssd1 vccd1 vccd1 _05593_/A sky130_fd_sc_hd__or2_1
XFILLER_138_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _08278_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08278_/Y sky130_fd_sc_hd__nand2_1
X_07229_ _07229_/A _07229_/B _07244_/A vssd1 vssd1 vccd1 vccd1 _07231_/B sky130_fd_sc_hd__and3_1
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ _10246_/C _10238_/X _10239_/Y vssd1 vssd1 vccd1 vccd1 _10240_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10171_ _07747_/A _10167_/X _10170_/X _10884_/Q vssd1 vssd1 vccd1 vccd1 _10884_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08656__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06176__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07840__C1 _07839_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10507_ _06147_/X _10496_/X _10506_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10974_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10438_ _06143_/X _10440_/B _05977_/X vssd1 vssd1 vccd1 vccd1 _10438_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10369_ _10369_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__and2_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06600_ _06600_/A vssd1 vssd1 vccd1 vccd1 _06775_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ _07580_/A _07580_/B vssd1 vssd1 vccd1 vccd1 _07581_/B sky130_fd_sc_hd__nand2_1
X_06531_ _06521_/A _06519_/A _06507_/A vssd1 vssd1 vccd1 vccd1 _06532_/B sky130_fd_sc_hd__o21bai_1
X_09250_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09276_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_61_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08201_ _08201_/A vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__clkbuf_2
X_06462_ _06470_/A _06462_/B vssd1 vssd1 vccd1 vccd1 _06479_/B sky130_fd_sc_hd__xor2_1
XFILLER_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05413_ _10620_/Q _05487_/A _05485_/A _10619_/Q _05412_/X vssd1 vssd1 vccd1 vccd1
+ _05413_/X sky130_fd_sc_hd__o221a_1
X_09181_ _07988_/A _09226_/S _09203_/A _09180_/X vssd1 vssd1 vccd1 vccd1 _09181_/X
+ sky130_fd_sc_hd__o211a_1
X_06393_ _06393_/A _06393_/B vssd1 vssd1 vccd1 vccd1 _06394_/B sky130_fd_sc_hd__xor2_1
X_08132_ _08132_/A _08132_/B vssd1 vssd1 vccd1 vccd1 _08132_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05344_ _10636_/Q vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__clkbuf_2
X_08063_ _08075_/B _08072_/B _08306_/B _08062_/X vssd1 vssd1 vccd1 vccd1 _08063_/X
+ sky130_fd_sc_hd__a31o_1
X_05275_ _10652_/Q vssd1 vssd1 vccd1 vccd1 _05291_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__10981__D _10981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07014_ _07039_/C vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08965_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08965_/Y sky130_fd_sc_hd__nor2_4
X_07916_ _07916_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _10643_/D sky130_fd_sc_hd__nor2_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08896_ _10826_/Q _08902_/B vssd1 vssd1 vccd1 vccd1 _08896_/X sky130_fd_sc_hd__xor2_2
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10071__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07847_ _07827_/X _05461_/C _07844_/X hold4/X vssd1 vssd1 vccd1 vccd1 _10625_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07778_ _07778_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07787_/A sky130_fd_sc_hd__xnor2_1
XFILLER_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06729_ _06729_/A _06729_/B vssd1 vssd1 vccd1 vccd1 _06752_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09517_ _09516_/B _09516_/C _09516_/A vssd1 vssd1 vccd1 vccd1 _09562_/C sky130_fd_sc_hd__a21o_1
XANTENNA__08311__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08862__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09448_ _09448_/A _09448_/B vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__xnor2_2
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09379_ _10896_/Q _09379_/B vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__and2b_1
XFILLER_40_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07822__C1 _07821_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ _10224_/A _10935_/Q vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10185__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _10154_/A _10154_/B vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input43_A io_wbs_m2s_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07555__A _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10488__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10987_ _10987_/CLK _10987_/D vssd1 vssd1 vccd1 vccd1 _10987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08853__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08747_/X _08749_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10807_/D sky130_fd_sc_hd__o21a_1
X_05962_ input10/X _09142_/B vssd1 vssd1 vccd1 vccd1 _07967_/A sky130_fd_sc_hd__or2_2
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05893_ _10656_/Q vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__buf_2
X_08681_ _08679_/X _08680_/Y _08669_/B _08670_/C vssd1 vssd1 vccd1 vccd1 _08683_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__10479__A1 _06124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07701_ _09759_/A _09759_/B _07700_/Y vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__a21o_1
XFILLER_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07632_ _07715_/D _07632_/B vssd1 vssd1 vccd1 vccd1 _07633_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06809__A _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__D _10976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07563_ _07563_/A _07727_/B _07563_/C vssd1 vssd1 vccd1 vccd1 _07563_/X sky130_fd_sc_hd__and3_1
X_09302_ _10497_/A _09302_/B vssd1 vssd1 vccd1 vccd1 _09303_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07494_ _07508_/B _07508_/A vssd1 vssd1 vccd1 vccd1 _07506_/A sky130_fd_sc_hd__or2b_1
X_06514_ _06527_/A _06522_/B _06517_/B _06567_/A vssd1 vssd1 vccd1 vccd1 _06523_/B
+ sky130_fd_sc_hd__a22o_1
X_09233_ _08256_/A _09231_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09233_/X sky130_fd_sc_hd__mux2_1
X_06445_ _10975_/Q _06576_/B vssd1 vssd1 vccd1 vccd1 _06675_/A sky130_fd_sc_hd__nand2_1
X_09164_ _10959_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09164_/Y sky130_fd_sc_hd__nor2_1
X_08115_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08130_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10403__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06376_ _06517_/B vssd1 vssd1 vccd1 vccd1 _06513_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05327_ _10643_/Q vssd1 vssd1 vccd1 vccd1 _07914_/A sky130_fd_sc_hd__clkbuf_2
X_09095_ _09769_/A vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08046_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08248_/A sky130_fd_sc_hd__buf_2
XFILLER_123_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09021__A1 _06066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09997_ _10138_/B _09997_/B vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08948_ _08968_/A vssd1 vssd1 vccd1 vccd1 _08948_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08879_ input32/X _08830_/X _08831_/X _08876_/A vssd1 vssd1 vccd1 vccd1 _08879_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08918__B _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10910_ _10924_/CLK _10910_/D vssd1 vssd1 vccd1 vccd1 _10910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10841_ _10841_/CLK _10841_/D vssd1 vssd1 vccd1 vccd1 _10841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10772_ _10833_/CLK _10772_/D vssd1 vssd1 vccd1 vccd1 _10772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ _10197_/A _10196_/B _10204_/X vssd1 vssd1 vccd1 vccd1 _10206_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_79_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _10137_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__xnor2_1
XFILLER_94_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _10068_/A _10068_/B vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06230_ input29/X _06225_/X _06229_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10605_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_19_clock_A _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10646_/CLK sky130_fd_sc_hd__clkbuf_16
X_06161_ _05982_/A _06158_/X _06160_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10589_/D
+ sky130_fd_sc_hd__o211a_1
X_06092_ _08037_/A vssd1 vssd1 vccd1 vccd1 _06117_/C sky130_fd_sc_hd__buf_2
XFILLER_105_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09920_ _10894_/Q _09920_/B vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__and2b_1
XFILLER_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08211__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09851_ _09851_/A _09851_/B _09851_/C vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__nor3_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08802_ _10815_/Q _08856_/B vssd1 vssd1 vccd1 vccd1 _08802_/Y sky130_fd_sc_hd__nor2_1
X_06994_ _10909_/Q vssd1 vssd1 vccd1 vccd1 _07028_/A sky130_fd_sc_hd__clkbuf_2
X_09782_ _09780_/X _09781_/Y _09718_/Y _09713_/B vssd1 vssd1 vccd1 vccd1 _09784_/A
+ sky130_fd_sc_hd__a211oi_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05945_ _08324_/A _05839_/X _05836_/X _08339_/B _05944_/X vssd1 vssd1 vccd1 vccd1
+ _05945_/X sky130_fd_sc_hd__o221a_1
X_08733_ _08918_/B vssd1 vssd1 vccd1 vccd1 _08928_/B sky130_fd_sc_hd__clkbuf_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10840__CLK _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05876_ _05848_/B _05823_/A _05875_/Y vssd1 vssd1 vccd1 vccd1 _05876_/X sky130_fd_sc_hd__o21a_1
X_08664_ _08778_/A vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__buf_2
XFILLER_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08595_ _10784_/Q _10783_/Q vssd1 vssd1 vccd1 vccd1 _08623_/C sky130_fd_sc_hd__and2_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07615_ _07615_/A _07615_/B vssd1 vssd1 vccd1 vccd1 _09898_/B sky130_fd_sc_hd__xnor2_4
XFILLER_41_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07546_ _07545_/B _07546_/B vssd1 vssd1 vccd1 vccd1 _07547_/B sky130_fd_sc_hd__and2b_1
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ _10816_/Q _09210_/X _09212_/X _09203_/X _09215_/X vssd1 vssd1 vccd1 vccd1
+ _09217_/B sky130_fd_sc_hd__a32o_1
X_07477_ _07477_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07480_/B sky130_fd_sc_hd__xnor2_1
XFILLER_22_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06428_ _06800_/A _06428_/B _06690_/A vssd1 vssd1 vccd1 vccd1 _06656_/A sky130_fd_sc_hd__and3_1
X_09147_ _09113_/X _09146_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09147_/Y sky130_fd_sc_hd__o21ai_1
X_06359_ _09302_/B _06736_/A vssd1 vssd1 vccd1 vccd1 _06359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09078_ _09078_/A _09078_/B vssd1 vssd1 vccd1 vccd1 _09078_/Y sky130_fd_sc_hd__nand2_1
X_08029_ _08029_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10524__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10824_ _10847_/CLK _10824_/D vssd1 vssd1 vccd1 vccd1 _10824_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10755_ _10791_/CLK _10755_/D vssd1 vssd1 vccd1 vccd1 _10755_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_20_clock_A _10857_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ _10841_/CLK _10686_/D vssd1 vssd1 vccd1 vccd1 _10686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06047__B2 _08018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05730_ _08095_/A vssd1 vssd1 vccd1 vccd1 _08093_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_36_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05661_ _08169_/B _05623_/X _05617_/X _08169_/A _05660_/X vssd1 vssd1 vccd1 vccd1
+ _05661_/X sky130_fd_sc_hd__o221a_1
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08380_ _08394_/A vssd1 vssd1 vccd1 vccd1 _08380_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07400_ _07406_/A _07753_/A _07399_/X vssd1 vssd1 vccd1 vccd1 _07404_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05592_ _10563_/Q _05596_/A vssd1 vssd1 vccd1 vccd1 _05593_/B sky130_fd_sc_hd__nand2_1
X_07331_ _07331_/A _07331_/B vssd1 vssd1 vccd1 vccd1 _07333_/B sky130_fd_sc_hd__and2_1
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09389__B _09396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ _07169_/A _07197_/B _07186_/B _07166_/A vssd1 vssd1 vccd1 vccd1 _07262_/X
+ sky130_fd_sc_hd__a22o_1
X_06213_ _06253_/B vssd1 vssd1 vccd1 vccd1 _06223_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09001_ _10713_/Q _08990_/C _09000_/X vssd1 vssd1 vccd1 vccd1 _09001_/X sky130_fd_sc_hd__o21a_1
X_07193_ _07193_/A _07193_/B vssd1 vssd1 vccd1 vccd1 _07194_/A sky130_fd_sc_hd__nand2_1
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07918__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06144_ _10586_/Q vssd1 vssd1 vccd1 vccd1 _06145_/A sky130_fd_sc_hd__inv_2
X_06075_ _10677_/Q vssd1 vssd1 vccd1 vccd1 _08029_/A sky130_fd_sc_hd__inv_2
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _09903_/A vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_113_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09834_ _09834_/A _09834_/B _09977_/B _09903_/A vssd1 vssd1 vccd1 vccd1 _09835_/B
+ sky130_fd_sc_hd__and4_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09765_ _09763_/C _09829_/A vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__and2b_1
X_06977_ _10903_/Q vssd1 vssd1 vccd1 vccd1 _07066_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05928_ _08188_/A _05884_/Y _05878_/Y _05877_/A _05927_/X vssd1 vssd1 vccd1 vccd1
+ _05928_/X sky130_fd_sc_hd__o221a_1
X_08716_ _08789_/B vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__clkbuf_2
X_09696_ _09696_/A vssd1 vssd1 vccd1 vccd1 _09769_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05859_ _10668_/Q _05863_/B vssd1 vssd1 vccd1 vccd1 _05859_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09160__B1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _10796_/Q _08600_/A _08643_/C _10797_/Q vssd1 vssd1 vccd1 vccd1 _08649_/B
+ sky130_fd_sc_hd__a31o_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _10779_/Q _10778_/Q _08578_/C _08578_/D vssd1 vssd1 vccd1 vccd1 _08585_/C
+ sky130_fd_sc_hd__and4_1
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07529_ _07529_/A _07529_/B vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__or2_1
X_10540_ _10839_/CLK _10540_/D vssd1 vssd1 vccd1 vccd1 _10540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ _06202_/X _10459_/X _10469_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10961_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06029__A1 _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07828__A _07849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06201__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05811__A _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08394__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10807_ _10811_/CLK _10807_/D vssd1 vssd1 vccd1 vccd1 _10807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10738_ _10791_/CLK _10738_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10669_ _10669_/CLK _10669_/D vssd1 vssd1 vccd1 vccd1 _10669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06900_ _06900_/A vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__buf_2
XANTENNA__08193__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07880_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _10633_/D sky130_fd_sc_hd__nor2_1
XFILLER_95_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06831_ _06875_/A _06875_/B vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__and2b_1
XFILLER_55_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06762_ _06762_/A _06762_/B vssd1 vssd1 vccd1 vccd1 _06763_/B sky130_fd_sc_hd__xor2_2
X_09550_ _09610_/C vssd1 vssd1 vccd1 vccd1 _09760_/B sky130_fd_sc_hd__clkbuf_2
X_05713_ _10549_/Q _08139_/A _08146_/A _05712_/Y vssd1 vssd1 vccd1 vccd1 _05713_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_08501_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__clkbuf_4
X_09481_ _09479_/A _09479_/B _09480_/X vssd1 vssd1 vccd1 vccd1 _09481_/X sky130_fd_sc_hd__a21o_1
X_08432_ _08432_/A _08432_/B _08578_/C vssd1 vssd1 vccd1 vccd1 _08432_/Y sky130_fd_sc_hd__nor3b_1
X_06693_ _06693_/A _06693_/B vssd1 vssd1 vccd1 vccd1 _06915_/A sky130_fd_sc_hd__xor2_1
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05644_ _05913_/A _05644_/B vssd1 vssd1 vccd1 vccd1 _05644_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06817__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ _08363_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__and2_1
X_05575_ _10568_/Q _05769_/A _05582_/B _10569_/Q vssd1 vssd1 vccd1 vccd1 _05576_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_51_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10984__D _10984_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _08294_/A vssd1 vssd1 vccd1 vccd1 _10703_/D sky130_fd_sc_hd__clkbuf_1
X_07314_ _07344_/A _07344_/B _07345_/B _07313_/A vssd1 vssd1 vccd1 vccd1 _07347_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07245_ _07264_/A _07264_/B _07269_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07254_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07759__A1 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _07176_/A _07176_/B vssd1 vssd1 vccd1 vccd1 _07200_/B sky130_fd_sc_hd__nand2_1
XFILLER_117_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06127_ input9/X _10432_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__and3_4
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06058_ _10666_/Q vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__buf_2
XFILLER_120_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08184__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08184__B2 _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__xnor2_1
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08198__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _09749_/A _09749_/B vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__nor2_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09679_ _09679_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__xor2_1
XFILLER_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08239__A2 _08212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 io_wbs_m2s_data[12] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_2
X_10523_ _10523_/A vssd1 vssd1 vccd1 vccd1 _10533_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_10_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10454_ _10955_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10454_/X sky130_fd_sc_hd__or2_1
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10385_ _10365_/X _10715_/Q _10383_/X _10384_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10934_/D sky130_fd_sc_hd__o221a_1
XFILLER_104_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05360_ _06052_/A _05848_/B vssd1 vssd1 vccd1 vccd1 _05360_/X sky130_fd_sc_hd__xor2_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07989__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05291_ _05291_/A _10576_/Q vssd1 vssd1 vccd1 vccd1 _05397_/B sky130_fd_sc_hd__nor2_1
X_07030_ _07169_/A _07166_/A _07030_/C _07417_/A vssd1 vssd1 vccd1 vccd1 _07031_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_127_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08981_ _08981_/A vssd1 vssd1 vccd1 vccd1 _09078_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_87_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07932_ _09016_/A _09013_/A vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__or2_1
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07863_ _06197_/A _07849_/X _07850_/X _07862_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ _07863_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_56_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10979__D _10979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06814_ _06814_/A _06853_/B vssd1 vssd1 vccd1 vccd1 _07766_/B sky130_fd_sc_hd__xnor2_2
X_09602_ _09780_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09533_ _10967_/Q _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__and3_1
X_07794_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07796_/B sky130_fd_sc_hd__nor2_1
X_06745_ _07675_/A _06745_/B vssd1 vssd1 vccd1 vccd1 _06746_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06676_ _06674_/A _06674_/C _06681_/A vssd1 vssd1 vccd1 vccd1 _06678_/C sky130_fd_sc_hd__a21o_1
X_09464_ _09501_/A _09464_/B vssd1 vssd1 vccd1 vccd1 _09466_/B sky130_fd_sc_hd__or2_1
X_05627_ _10688_/Q vssd1 vssd1 vccd1 vccd1 _05896_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09395_ _09678_/A vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08415_ input1/X input49/X input14/X _08415_/D vssd1 vssd1 vccd1 vccd1 _08989_/B
+ sky130_fd_sc_hd__and4_4
X_08346_ _08344_/X _08346_/B vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__and2b_1
XANTENNA__10069__A _10069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05558_ _10562_/Q _10561_/Q _05602_/A vssd1 vssd1 vccd1 vccd1 _05596_/A sky130_fd_sc_hd__or3_1
X_08277_ _08277_/A _08277_/B _08277_/C vssd1 vssd1 vccd1 vccd1 _08295_/C sky130_fd_sc_hd__and3_1
X_05489_ _05489_/A vssd1 vssd1 vccd1 vccd1 _05489_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_67_clock_A _10981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07228_ _07232_/A _07232_/B _07225_/X vssd1 vssd1 vccd1 vccd1 _07231_/A sky130_fd_sc_hd__a21o_1
XFILLER_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07159_ _07229_/A _07164_/B _07178_/A _07188_/A vssd1 vssd1 vccd1 vccd1 _07159_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10170_ _10177_/A vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_105_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08002__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10506_ _10506_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__or2_1
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10437_ _06008_/X _10431_/X _10436_/X _08563_/X vssd1 vssd1 vccd1 vccd1 _10948_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10368_ _10931_/Q _10379_/B vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__and2_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10442__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ _10301_/A _10289_/X _10300_/A vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__o21ba_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06530_ _06541_/C _06528_/Y _06529_/X vssd1 vssd1 vccd1 vccd1 _06533_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08320__A1 _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__B2 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06461_ _06472_/A _06461_/B _06547_/C vssd1 vssd1 vccd1 vccd1 _06462_/B sky130_fd_sc_hd__and3b_1
X_08200_ _08114_/X _08207_/B _08196_/X _08199_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08200_/X sky130_fd_sc_hd__o311a_1
X_05412_ _10619_/Q _05485_/A _05402_/X _05411_/X vssd1 vssd1 vccd1 vccd1 _05412_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09180_ _05460_/C _09136_/X _09148_/X _08191_/A _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09180_/X sky130_fd_sc_hd__a221o_1
X_06392_ _10515_/A _06627_/B vssd1 vssd1 vccd1 vccd1 _06393_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08084__B1 _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _08092_/X _08129_/X _08139_/B _08096_/X vssd1 vssd1 vccd1 vccd1 _08131_/X
+ sky130_fd_sc_hd__a31o_1
X_05343_ _08013_/A _05854_/A vssd1 vssd1 vccd1 vccd1 _05343_/Y sky130_fd_sc_hd__xnor2_1
X_08062_ _08062_/A vssd1 vssd1 vccd1 vccd1 _08062_/X sky130_fd_sc_hd__buf_4
X_05274_ _10654_/Q vssd1 vssd1 vccd1 vccd1 _05388_/A sky130_fd_sc_hd__clkinv_2
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07013_ _07013_/A _07013_/B vssd1 vssd1 vccd1 vccd1 _07039_/C sky130_fd_sc_hd__xnor2_2
XFILLER_127_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08964_ _08964_/A vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_130_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07915_ _10611_/Q _07906_/X _07910_/X _07914_/Y vssd1 vssd1 vccd1 vccd1 _07916_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08895_ _08893_/X _08894_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10825_/D sky130_fd_sc_hd__o21a_1
XFILLER_96_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07846_ hold3/X _07828_/X _07829_/X _07845_/Y _07832_/X vssd1 vssd1 vccd1 vccd1 hold4/A
+ sky130_fd_sc_hd__o221ai_4
XFILLER_56_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07777_ _07777_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07778_/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06728_ _06734_/A _06734_/B _06320_/Y _06321_/A vssd1 vssd1 vccd1 vccd1 _06729_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09516_ _09516_/A _09516_/B _09516_/C vssd1 vssd1 vccd1 vccd1 _09562_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08311__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09447_ _09678_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09448_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06659_ _06660_/A _06660_/B vssd1 vssd1 vccd1 vccd1 _06661_/A sky130_fd_sc_hd__and2_1
XANTENNA__08492__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09378_ _09921_/B _09922_/B _10065_/B _09377_/X vssd1 vssd1 vccd1 vccd1 _10063_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08329_ _08339_/C _08329_/B vssd1 vssd1 vccd1 vccd1 _08329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10222_ _10951_/Q vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__inv_2
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10153_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10154_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10084_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__or2_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input36_A io_wbs_m2s_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07571__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06187__A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ _10986_/CLK _10986_/D vssd1 vssd1 vccd1 vccd1 _10986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08081__A3 _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05961_ input11/X input13/X input12/X vssd1 vssd1 vccd1 vccd1 _09142_/B sky130_fd_sc_hd__or3_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07700_ _07700_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _07700_/Y sky130_fd_sc_hd__nor2_1
X_05892_ _08169_/B _05892_/B vssd1 vssd1 vccd1 vccd1 _05892_/X sky130_fd_sc_hd__and2_1
X_08680_ _10801_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07631_ _07698_/A _07698_/B vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__xnor2_2
XFILLER_80_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07562_ _07562_/A _07729_/B _07562_/C vssd1 vssd1 vccd1 vccd1 _07563_/C sky130_fd_sc_hd__and3_1
XANTENNA__08829__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__buf_2
X_06513_ _06527_/A _06600_/A _06522_/B _06513_/D vssd1 vssd1 vccd1 vccd1 _06532_/A
+ sky130_fd_sc_hd__nand4_2
X_07493_ _07493_/A _07493_/B vssd1 vssd1 vccd1 vccd1 _07508_/A sky130_fd_sc_hd__xor2_2
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09232_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09257_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__06825__A _06845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06444_ _10976_/Q _06587_/A _06947_/A vssd1 vssd1 vccd1 vccd1 _06472_/B sky130_fd_sc_hd__and3_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09163_ _09202_/A _09163_/B vssd1 vssd1 vccd1 vccd1 _10845_/D sky130_fd_sc_hd__nor2_4
X_06375_ _06375_/A _06387_/B vssd1 vssd1 vccd1 vccd1 _06517_/B sky130_fd_sc_hd__xnor2_4
XFILLER_135_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08114_/X sky130_fd_sc_hd__buf_2
X_05326_ _05830_/A _05831_/B vssd1 vssd1 vccd1 vccd1 _05326_/X sky130_fd_sc_hd__xor2_1
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09094_ _10970_/Q vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08045_ _05475_/X _08044_/X _06033_/X vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__a21o_1
XFILLER_116_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09996_ _10123_/A _09919_/B _10122_/B _10487_/A vssd1 vssd1 vccd1 vccd1 _09997_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09309__B1 _09396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08947_ _08947_/A vssd1 vssd1 vccd1 vccd1 _10430_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08487__A _08935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _08883_/A _08876_/Y _08871_/Y _08873_/Y vssd1 vssd1 vccd1 vccd1 _08878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07829_ _07850_/A vssd1 vssd1 vccd1 vccd1 _07829_/X sky130_fd_sc_hd__buf_4
XFILLER_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10840_ _10840_/CLK _10840_/D vssd1 vssd1 vccd1 vccd1 _10840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10771_ _10855_/CLK _10771_/D vssd1 vssd1 vccd1 vccd1 _10771_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06846__A1 _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09111__A _09111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08063__A3 _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06074__A2 _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08220__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10205_ _10191_/B _10204_/X _10196_/B vssd1 vssd1 vccd1 vccd1 _10226_/A sky130_fd_sc_hd__a21o_1
XFILLER_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _10491_/A _10129_/B _10061_/A _10059_/A vssd1 vssd1 vccd1 vccd1 _10137_/B
+ sky130_fd_sc_hd__a31o_1
X_10067_ _10131_/B _10067_/B vssd1 vssd1 vccd1 vccd1 _10068_/B sky130_fd_sc_hd__xnor2_2
XFILLER_48_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10969_ _10970_/CLK _10969_/D vssd1 vssd1 vccd1 vccd1 _10969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08039__B1 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10167__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06160_ _06160_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06160_/Y sky130_fd_sc_hd__nand2_1
X_06091_ _10580_/Q vssd1 vssd1 vccd1 vccd1 _08037_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08333__C_N _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09850_ _09851_/A _09851_/B _09851_/C vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__o21a_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08801_ _10815_/Q _08801_/B vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__and2_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06993_ _06993_/A vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__clkbuf_2
X_09781_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__nand2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05944_ _05939_/X _05940_/X _05942_/X _05943_/X vssd1 vssd1 vccd1 vccd1 _05944_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_112_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08732_ _10806_/Q _08732_/B vssd1 vssd1 vccd1 vccd1 _08740_/C sky130_fd_sc_hd__xor2_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10987__D _10987_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _10799_/Q _08658_/X _08662_/X vssd1 vssd1 vccd1 vccd1 _10799_/D sky130_fd_sc_hd__a21boi_1
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05875_ _08198_/A _05878_/B _10663_/Q vssd1 vssd1 vccd1 vccd1 _05875_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_94_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10321__A1 _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _10783_/Q _08550_/X _08593_/Y vssd1 vssd1 vccd1 vccd1 _10783_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ _07620_/A _06962_/B _07624_/A vssd1 vssd1 vccd1 vccd1 _07615_/B sky130_fd_sc_hd__a21oi_2
XFILLER_81_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07545_ _07546_/B _07545_/B vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__and2b_1
XFILLER_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07476_ _07589_/A vssd1 vssd1 vccd1 vccd1 _07480_/A sky130_fd_sc_hd__inv_2
X_09215_ _08000_/A _09214_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__mux2_1
X_06427_ _06690_/A _06630_/A _06425_/Y _06428_/B _06800_/A vssd1 vssd1 vccd1 vccd1
+ _06631_/A sky130_fd_sc_hd__o2111a_1
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09146_ _09114_/X _09145_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__o21a_1
X_06358_ _06558_/B _06558_/C vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05309_ _10672_/Q _05340_/A vssd1 vssd1 vccd1 vccd1 _05336_/A sky130_fd_sc_hd__or2_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09077_ _08119_/A _08976_/X _09076_/X _09078_/B vssd1 vssd1 vccd1 vccd1 _09077_/X
+ sky130_fd_sc_hd__a211o_1
X_06289_ _10928_/Q _10911_/Q vssd1 vssd1 vccd1 vccd1 _06851_/A sky130_fd_sc_hd__or2_1
XFILLER_123_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08028_ input36/X _07985_/B _08027_/X _08019_/X vssd1 vssd1 vccd1 vccd1 _10676_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _10049_/C _09976_/Y _09978_/X vssd1 vssd1 vccd1 vccd1 _09980_/B sky130_fd_sc_hd__o21a_1
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10823_ _10823_/CLK _10823_/D vssd1 vssd1 vccd1 vccd1 _10823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10754_ _10798_/CLK _10754_/D vssd1 vssd1 vccd1 vccd1 _10754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10685_ _10839_/CLK _10685_/D vssd1 vssd1 vccd1 vccd1 _10685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10119_ _10107_/A _10107_/B _10118_/X vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__a21oi_2
XFILLER_76_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05660_ _08148_/A _05626_/X _05623_/X _10690_/Q _05659_/X vssd1 vssd1 vccd1 vccd1
+ _05660_/X sky130_fd_sc_hd__a221o_1
XFILLER_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05591_ _10702_/Q vssd1 vssd1 vccd1 vccd1 _08277_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07330_ _07330_/A _07335_/A vssd1 vssd1 vccd1 vccd1 _07331_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09000_ _10766_/Q _08418_/B _09168_/A _10800_/Q _08999_/X vssd1 vssd1 vccd1 vccd1
+ _09000_/X sky130_fd_sc_hd__a221o_1
X_07261_ _07273_/A _07273_/B vssd1 vssd1 vccd1 vccd1 _07318_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07483__A1 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07483__B2 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06212_ _10517_/A _06212_/B vssd1 vssd1 vccd1 vccd1 _06253_/B sky130_fd_sc_hd__nor2_4
XANTENNA__08590__A _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ _07192_/A _07192_/B vssd1 vssd1 vccd1 vccd1 _07194_/B sky130_fd_sc_hd__xnor2_1
XFILLER_117_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06143_ _10526_/A vssd1 vssd1 vccd1 vccd1 _06143_/X sky130_fd_sc_hd__buf_4
XANTENNA__08983__A1 _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06074_ _10711_/Q _08034_/A _07979_/A _05709_/Y _06073_/X vssd1 vssd1 vccd1 vccd1
+ _06082_/A sky130_fd_sc_hd__a221o_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _10023_/A _09829_/A vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__or2b_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09833_ _09834_/A _09977_/B _09903_/A _10057_/A vssd1 vssd1 vccd1 vccd1 _09835_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09764_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__nand2_1
X_06976_ _10906_/Q vssd1 vssd1 vccd1 vccd1 _06997_/B sky130_fd_sc_hd__buf_2
XFILLER_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05927_ _10693_/Q _05884_/Y _05888_/X _05926_/X vssd1 vssd1 vccd1 vccd1 _05927_/X
+ sky130_fd_sc_hd__a22o_1
X_08715_ _08744_/B vssd1 vssd1 vccd1 vccd1 _08789_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__08499__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ _09646_/B _09695_/B vssd1 vssd1 vccd1 vccd1 _09707_/A sky130_fd_sc_hd__and2b_1
XFILLER_26_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05858_ _05858_/A _05858_/B vssd1 vssd1 vccd1 vccd1 _05858_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09160__A1 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08646_ _08648_/B _08646_/B vssd1 vssd1 vccd1 vccd1 _10796_/D sky130_fd_sc_hd__nor2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05789_ _05789_/A _05764_/A vssd1 vssd1 vccd1 vccd1 _05789_/X sky130_fd_sc_hd__or2b_1
X_08577_ _08583_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _10778_/D sky130_fd_sc_hd__nor2_1
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07528_ _07528_/A _07528_/B _07528_/C vssd1 vssd1 vccd1 vccd1 _07529_/B sky130_fd_sc_hd__and3_1
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07459_ _09304_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07460_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10470_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06029__A2 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ _08748_/X _08985_/X _08988_/X _10720_/Q _09128_/X vssd1 vssd1 vccd1 vccd1
+ _09129_/X sky130_fd_sc_hd__a221o_1
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10535__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07844__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06737__B1 _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__A4 _08701_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_42_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10676_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09151__B2 _10722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ _10806_/CLK _10806_/D vssd1 vssd1 vccd1 vccd1 _10806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06195__A input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10970_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__08662__B1 _08820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ _10737_/CLK _10737_/D vssd1 vssd1 vccd1 vccd1 _10737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05476__B1 _05474_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10668_ _10702_/CLK _10668_/D vssd1 vssd1 vccd1 vccd1 _10668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _10811_/CLK _10599_/D vssd1 vssd1 vccd1 vccd1 _10599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05779__B2 _05778_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06830_ _06844_/C _06856_/C _06884_/A vssd1 vssd1 vccd1 vccd1 _06875_/B sky130_fd_sc_hd__o21bai_2
XFILLER_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06761_ _06772_/A _06786_/A _06856_/A vssd1 vssd1 vccd1 vccd1 _06762_/B sky130_fd_sc_hd__and3b_1
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05712_ _10550_/Q vssd1 vssd1 vccd1 vccd1 _05712_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08500_ _08633_/A vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__buf_2
X_09480_ _09757_/A vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__clkbuf_4
X_06692_ _06692_/A _06692_/B vssd1 vssd1 vccd1 vccd1 _06693_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05643_ _05643_/A _10541_/Q vssd1 vssd1 vccd1 vccd1 _05644_/B sky130_fd_sc_hd__xor2_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08431_ _10729_/Q _08565_/C vssd1 vssd1 vccd1 vccd1 _08578_/C sky130_fd_sc_hd__and2_1
XFILLER_64_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08362_ input40/X _08123_/X _08109_/X _05528_/X _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08363_/B sky130_fd_sc_hd__o221a_1
X_05574_ _08332_/A vssd1 vssd1 vccd1 vccd1 _05574_/X sky130_fd_sc_hd__clkbuf_2
X_08293_ _08291_/X _08293_/B vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__and2b_1
X_07313_ _07313_/A _07313_/B vssd1 vssd1 vccd1 vccd1 _07345_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ _07244_/A _07244_/B vssd1 vssd1 vccd1 vccd1 _07269_/B sky130_fd_sc_hd__xor2_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10355__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07175_ _07193_/A _07175_/B vssd1 vssd1 vccd1 vccd1 _07176_/B sky130_fd_sc_hd__nand2_1
X_06126_ input7/X input4/X _07967_/A _06126_/D vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__nor4_4
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06057_ _10668_/Q vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__buf_2
XFILLER_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09816_ _09961_/A _09753_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__o21a_1
XFILLER_100_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09747_ _10478_/A _09672_/B _10129_/B _09670_/Y vssd1 vssd1 vccd1 vccd1 _09749_/B
+ sky130_fd_sc_hd__a31oi_1
XANTENNA_clkbuf_leaf_63_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ _07636_/A _07635_/B vssd1 vssd1 vccd1 vccd1 _07629_/B sky130_fd_sc_hd__nor2_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09678_ _09678_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09679_/B sky130_fd_sc_hd__nand2_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _10792_/Q _08631_/C _08642_/D _08550_/X vssd1 vssd1 vccd1 vccd1 _08630_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _10522_/A vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10453_ _06168_/X _10446_/X _10452_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10954_/D
+ sky130_fd_sc_hd__o211a_1
X_10384_ _10528_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__a21bo_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06186__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05822__A _05886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06918__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05290_ _05818_/A _05910_/B _05289_/Y vssd1 vssd1 vccd1 vccd1 _05398_/A sky130_fd_sc_hd__a21oi_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05269__A _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08980_ _05736_/A _06212_/B _08976_/X vssd1 vssd1 vccd1 vccd1 _08980_/Y sky130_fd_sc_hd__a21oi_1
X_07931_ _08944_/A _09142_/C vssd1 vssd1 vccd1 vccd1 _09013_/A sky130_fd_sc_hd__or2_1
XFILLER_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07862_ hold14/X _07866_/B vssd1 vssd1 vccd1 vccd1 _07862_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06177__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06813_ _06813_/A _06813_/B vssd1 vssd1 vccd1 vccd1 _06853_/B sky130_fd_sc_hd__xor2_4
X_09601_ _09599_/A _09692_/A _09761_/C _09805_/A vssd1 vssd1 vccd1 vccd1 _09602_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07793_ _06869_/A _06869_/B _06868_/A vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__a21oi_1
X_09532_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__xor2_2
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06744_ _06775_/A _06774_/B vssd1 vssd1 vccd1 vccd1 _06747_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06675_ _06675_/A _06675_/B vssd1 vssd1 vccd1 vccd1 _06678_/B sky130_fd_sc_hd__xor2_2
XFILLER_24_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09463_ _09462_/A _09462_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _09464_/B sky130_fd_sc_hd__a21oi_1
X_05626_ _05626_/A _05626_/B vssd1 vssd1 vccd1 vccd1 _05626_/X sky130_fd_sc_hd__and2_1
XFILLER_52_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09394_ _09424_/A vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08414_ _08414_/A vssd1 vssd1 vccd1 vccd1 _08415_/D sky130_fd_sc_hd__inv_2
X_08345_ input37/X _08248_/A _08052_/A _05570_/X _08175_/A vssd1 vssd1 vccd1 vccd1
+ _08346_/B sky130_fd_sc_hd__o221a_1
X_05557_ _10560_/Q _05604_/A vssd1 vssd1 vccd1 vccd1 _05602_/A sky130_fd_sc_hd__or2_1
XFILLER_51_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08276_ _08278_/A _08276_/B vssd1 vssd1 vccd1 vccd1 _08276_/Y sky130_fd_sc_hd__nor2_1
X_05488_ _05818_/B _05470_/B _05495_/A _05453_/A _05487_/Y vssd1 vssd1 vccd1 vccd1
+ _10545_/D sky130_fd_sc_hd__a221o_1
X_07227_ _07225_/X _07227_/B vssd1 vssd1 vccd1 vccd1 _07232_/B sky130_fd_sc_hd__and2b_1
XFILLER_105_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09051__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _07186_/A _07188_/A _07164_/B _07178_/A vssd1 vssd1 vccd1 vccd1 _07280_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06109_ _10705_/Q _08305_/B vssd1 vssd1 vccd1 vccd1 _08317_/B sky130_fd_sc_hd__or2_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07089_ _07089_/A _07089_/B vssd1 vssd1 vccd1 vccd1 _07090_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05915__A1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__A1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__B _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07569__A _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10505_ _06143_/X _10496_/X _10504_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10973_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10436_ _10948_/Q _10440_/B vssd1 vssd1 vccd1 vccd1 _10436_/X sky130_fd_sc_hd__or2_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10367_ _10427_/B vssd1 vssd1 vccd1 vccd1 _10379_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10298_ _10298_/A _10298_/B vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__nand2_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06460_ _10978_/Q _06460_/B _06670_/A vssd1 vssd1 vccd1 vccd1 _06479_/A sky130_fd_sc_hd__and3_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05411_ _10618_/Q _05483_/A _05407_/X _05410_/X vssd1 vssd1 vccd1 vccd1 _05411_/X
+ sky130_fd_sc_hd__a22o_1
X_08130_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08139_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06391_ _06489_/B vssd1 vssd1 vccd1 vccd1 _06627_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09281__A0 _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05342_ _10670_/Q vssd1 vssd1 vccd1 vccd1 _08013_/A sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_11_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08061_ _08061_/A vssd1 vssd1 vccd1 vccd1 _08306_/B sky130_fd_sc_hd__buf_2
X_05273_ _10655_/Q vssd1 vssd1 vccd1 vccd1 _05295_/A sky130_fd_sc_hd__inv_2
XANTENNA__09033__A0 _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07012_ _06997_/B _06997_/C _07007_/A vssd1 vssd1 vccd1 vccd1 _07013_/B sky130_fd_sc_hd__o21ai_1
XFILLER_88_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ _09092_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07914_ _07914_/A vssd1 vssd1 vccd1 vccd1 _07914_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08894_ input34/X _08830_/X _08831_/X _10825_/Q vssd1 vssd1 vccd1 vccd1 _08894_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07845_ _10875_/Q _07845_/B vssd1 vssd1 vccd1 vccd1 _07845_/Y sky130_fd_sc_hd__nand2_1
X_07776_ _10515_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07777_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09515_ _09514_/A _09514_/B _09514_/C vssd1 vssd1 vccd1 vccd1 _09516_/C sky130_fd_sc_hd__a21o_1
X_06727_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07761_/A sky130_fd_sc_hd__xnor2_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09446_ _09811_/B _09677_/B vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__or2_2
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06658_ _06658_/A _06658_/B vssd1 vssd1 vccd1 vccd1 _06660_/B sky130_fd_sc_hd__xnor2_1
X_05609_ _10557_/Q _05612_/A vssd1 vssd1 vccd1 vccd1 _05610_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08492__B _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ _10894_/Q _06993_/A vssd1 vssd1 vccd1 vccd1 _09377_/X sky130_fd_sc_hd__or2b_1
X_06589_ _06589_/A _06589_/B vssd1 vssd1 vccd1 vccd1 _06951_/B sky130_fd_sc_hd__or2_1
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08328_ _08324_/A _08327_/B _08067_/X vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__o21ai_1
XFILLER_138_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06086__B1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _08114_/X _08277_/C _08252_/Y _08257_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08259_/X sky130_fd_sc_hd__o311a_1
XFILLER_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10221_ _07113_/A _10115_/X _10220_/Y _10043_/X vssd1 vssd1 vccd1 vccd1 _10901_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10152_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10153_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10083_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input29_A io_wbs_m2s_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10985_ _10985_/CLK _10985_/D vssd1 vssd1 vccd1 vccd1 _10985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09015__A0 _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10419_ _06191_/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__a21bo_1
XFILLER_124_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05960_ _10369_/A vssd1 vssd1 vccd1 vccd1 _10432_/B sky130_fd_sc_hd__buf_2
XFILLER_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05891_ _05891_/A _05891_/B vssd1 vssd1 vccd1 vccd1 _05892_/B sky130_fd_sc_hd__and2_1
XFILLER_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06001__A0 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07630_ _07630_/A _07630_/B vssd1 vssd1 vccd1 vccd1 _07698_/B sky130_fd_sc_hd__xnor2_4
XFILLER_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07561_ _07729_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__nand2_1
X_09300_ _09300_/A vssd1 vssd1 vccd1 vccd1 _10865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06512_ _06541_/C _06512_/B vssd1 vssd1 vccd1 vccd1 _06620_/A sky130_fd_sc_hd__xnor2_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07492_ _07490_/A _07490_/B _07510_/A vssd1 vssd1 vccd1 vccd1 _07508_/B sky130_fd_sc_hd__o21ba_1
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09231_ _05598_/X _07889_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09231_/X sky130_fd_sc_hd__mux2_1
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06443_ _10975_/Q _06575_/B vssd1 vssd1 vccd1 vccd1 _06947_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09162_ _09112_/X _09158_/Y _09161_/X vssd1 vssd1 vccd1 vccd1 _09163_/B sky130_fd_sc_hd__a21oi_1
X_06374_ _06374_/A _06374_/B vssd1 vssd1 vccd1 vccd1 _06387_/B sky130_fd_sc_hd__xnor2_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08113_ _08113_/A vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__06068__B1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05325_ _10644_/Q vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09093_ _10515_/A _09118_/A vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__nor2_1
X_08044_ _08044_/A vssd1 vssd1 vccd1 vccd1 _08044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09995_ _10489_/A _10056_/C _10122_/B vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08946_ _09124_/A _08968_/A vssd1 vssd1 vccd1 vccd1 _08947_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08877_ _08871_/Y _08873_/Y _08883_/A _08876_/Y vssd1 vssd1 vccd1 vccd1 _08891_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_84_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07828_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07828_/X sky130_fd_sc_hd__buf_4
XFILLER_57_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07759_ _07635_/A _06966_/A _06966_/B vssd1 vssd1 vccd1 vccd1 _07764_/A sky130_fd_sc_hd__a21oi_2
X_10770_ _10855_/CLK _10770_/D vssd1 vssd1 vccd1 vccd1 _10770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09429_ _09429_/A _09460_/B vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__xnor2_2
XFILLER_138_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08950__B _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ _10948_/Q _10932_/Q vssd1 vssd1 vccd1 vccd1 _10204_/X sky130_fd_sc_hd__or2b_1
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10135_ _10049_/B _09880_/A _09976_/Y _09879_/B vssd1 vssd1 vccd1 vccd1 _10137_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10066_ _10066_/A _10131_/C vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__nor2_1
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06198__A _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10968_ _10968_/CLK _10968_/D vssd1 vssd1 vccd1 vccd1 _10968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05830__A _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ _10920_/CLK _10899_/D vssd1 vssd1 vccd1 vccd1 _10899_/Q sky130_fd_sc_hd__dfxtp_2
X_06090_ _06036_/X _06071_/X _06082_/X _06089_/X _10579_/Q vssd1 vssd1 vccd1 vccd1
+ _08065_/B sky130_fd_sc_hd__o41a_2
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08211__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05277__A _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08688_/X _08798_/X _08799_/X vssd1 vssd1 vccd1 vccd1 _10814_/D sky130_fd_sc_hd__o21a_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09780_ _09780_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__or2b_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _07021_/A vssd1 vssd1 vccd1 vccd1 _07574_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05943_ _08315_/A _05838_/B _05941_/Y _05839_/X _08327_/A vssd1 vssd1 vccd1 vccd1
+ _05943_/X sky130_fd_sc_hd__a32o_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08731_ _08727_/X _08730_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10805_/D sky130_fd_sc_hd__o21a_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08662_ _06124_/A _08819_/A _08820_/A _10799_/Q _09090_/A vssd1 vssd1 vccd1 vccd1
+ _08662_/X sky130_fd_sc_hd__o221a_1
X_05874_ _10661_/Q _05883_/A _05886_/A _05886_/B vssd1 vssd1 vccd1 vccd1 _05878_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ _07613_/A vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__inv_2
XFILLER_38_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08593_ _10783_/Q _08550_/X _08630_/A vssd1 vssd1 vccd1 vccd1 _08593_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07544_ _07544_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07545_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09212__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07475_ _07728_/A _07475_/B _07475_/C vssd1 vssd1 vccd1 vccd1 _07589_/A sky130_fd_sc_hd__and3_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09214_ _06061_/A _07878_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09214_/X sky130_fd_sc_hd__mux2_1
X_06426_ _06426_/A vssd1 vssd1 vccd1 vccd1 _06800_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09145_ _10941_/Q _09143_/Y _09144_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09145_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06357_ _06436_/A vssd1 vssd1 vccd1 vccd1 _06719_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05308_ _10671_/Q _10670_/Q _05854_/A vssd1 vssd1 vccd1 vccd1 _05340_/A sky130_fd_sc_hd__or3_1
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09076_ _05462_/B _09020_/B _06129_/B _08117_/A _09297_/S vssd1 vssd1 vccd1 vccd1
+ _09076_/X sky130_fd_sc_hd__o221a_1
X_06288_ _10929_/Q _10912_/Q vssd1 vssd1 vccd1 vccd1 _06288_/X sky130_fd_sc_hd__or2_1
XANTENNA__07667__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08027_/X sky130_fd_sc_hd__or2_1
XFILLER_104_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08202__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_opt_1_0_clock_A _10985_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__A0 _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ _09908_/A _10049_/B _10095_/A vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__a21bo_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08929_ _08920_/A _08927_/X _08928_/X vssd1 vssd1 vccd1 vccd1 _08929_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_92_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10822_ _10823_/CLK _10822_/D vssd1 vssd1 vccd1 vccd1 _10822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _10791_/CLK _10753_/D vssd1 vssd1 vccd1 vccd1 _10753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10684_ _10839_/CLK _10684_/D vssd1 vssd1 vccd1 vccd1 _10684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07401__C1 _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ _10104_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10118_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08201__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10049_ _10129_/A _10049_/B _10049_/C vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__and3_1
XFILLER_63_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05590_ _10564_/Q _05593_/A vssd1 vssd1 vccd1 vccd1 _05590_/X sky130_fd_sc_hd__xor2_1
XFILLER_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07260_ _07260_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _07273_/B sky130_fd_sc_hd__nor2_1
X_06211_ _09148_/A vssd1 vssd1 vccd1 vccd1 _06212_/B sky130_fd_sc_hd__buf_2
X_07191_ _07229_/A _07197_/B _07186_/B _07188_/A vssd1 vssd1 vccd1 vccd1 _07193_/B
+ sky130_fd_sc_hd__a22o_1
X_06142_ input38/X vssd1 vssd1 vccd1 vccd1 _10526_/A sky130_fd_sc_hd__buf_4
X_06073_ _05702_/A _08209_/A _05818_/A _08082_/A vssd1 vssd1 vccd1 vccd1 _06073_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ _09901_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08217__B1_N _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09832_ _09647_/A _09971_/A _09834_/A _09761_/C vssd1 vssd1 vccd1 vccd1 _09837_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09207__A _09228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09763_ _09908_/A _09947_/B _09763_/C vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__and3_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08714_ _10805_/Q _08744_/B vssd1 vssd1 vccd1 vccd1 _08740_/A sky130_fd_sc_hd__xor2_1
XFILLER_39_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06975_ _07086_/B vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05926_ _05885_/A _05888_/B _05889_/X _05692_/A _05925_/X vssd1 vssd1 vccd1 vccd1
+ _05926_/X sky130_fd_sc_hd__a221o_1
XFILLER_94_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09694_ _09904_/A _09828_/B _09647_/A _09693_/Y vssd1 vssd1 vccd1 vccd1 _09710_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05857_ _08268_/A _05857_/B vssd1 vssd1 vccd1 vccd1 _05858_/A sky130_fd_sc_hd__and2_1
XFILLER_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08645_ _10796_/Q _08638_/X _10192_/A vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__o21ai_1
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08576_ _10778_/Q _08576_/B vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__xor2_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05788_ _05788_/A _05788_/B _05788_/C _05802_/A vssd1 vssd1 vccd1 vccd1 _05788_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__10058__A1 _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07527_ _07648_/B _07527_/B _07643_/A vssd1 vssd1 vccd1 vccd1 _07638_/B sky130_fd_sc_hd__or3b_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07458_ _07493_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__xor2_1
XFILLER_22_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07389_ _07728_/A vssd1 vssd1 vccd1 vccd1 _07592_/A sky130_fd_sc_hd__buf_4
X_06409_ _06626_/A _06409_/B _06409_/C vssd1 vssd1 vccd1 vccd1 _06717_/A sky130_fd_sc_hd__and3_1
X_09128_ _07974_/A _09123_/X _09125_/X _09127_/X vssd1 vssd1 vccd1 vccd1 _09128_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ _10057_/A vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08021__A _08021_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input11_A io_wbs_m2s_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09439__B1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10805_ _10808_/CLK _10805_/D vssd1 vssd1 vccd1 vccd1 _10805_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10736_ _10737_/CLK _10736_/D vssd1 vssd1 vccd1 vccd1 _10736_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08662__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05476__A1 _10616_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05476__B2 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10667_ _10814_/CLK _10667_/D vssd1 vssd1 vccd1 vccd1 _10667_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10598_ _10819_/CLK _10598_/D vssd1 vssd1 vccd1 vccd1 _10598_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10221__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06760_ _06779_/A _06779_/B vssd1 vssd1 vccd1 vccd1 _06762_/A sky130_fd_sc_hd__and2b_1
X_05711_ _08146_/A vssd1 vssd1 vccd1 vccd1 _05711_/Y sky130_fd_sc_hd__inv_2
X_06691_ _06691_/A _06691_/B vssd1 vssd1 vccd1 vccd1 _06693_/A sky130_fd_sc_hd__nand2_1
X_05642_ _10680_/Q vssd1 vssd1 vccd1 vccd1 _05913_/A sky130_fd_sc_hd__inv_2
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08430_ _10774_/Q _10773_/Q _08559_/B vssd1 vssd1 vccd1 vccd1 _08565_/C sky130_fd_sc_hd__and3_1
XFILLER_64_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08361_ _10679_/Q _08044_/A _08359_/Y _08360_/X vssd1 vssd1 vccd1 vccd1 _08363_/A
+ sky130_fd_sc_hd__a211o_1
X_05573_ _08339_/B vssd1 vssd1 vccd1 vccd1 _08332_/A sky130_fd_sc_hd__buf_2
XFILLER_16_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08292_ input31/X _08212_/X _08052_/A _08287_/A _08175_/A vssd1 vssd1 vccd1 vccd1
+ _08293_/B sky130_fd_sc_hd__o221a_1
X_07312_ _07312_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07313_/B sky130_fd_sc_hd__and2_1
X_07243_ _07246_/A _07246_/B vssd1 vssd1 vccd1 vccd1 _07269_/A sky130_fd_sc_hd__nand2_1
XFILLER_118_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07174_ _07193_/A _07175_/B vssd1 vssd1 vccd1 vccd1 _07176_/A sky130_fd_sc_hd__or2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06125_ input8/X vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__buf_2
XFILLER_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06056_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__inv_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09815_ _09815_/A _09815_/B vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__xor2_2
XANTENNA_input3_A io_qei_ch_b vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09746_ _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__xnor2_1
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06958_ _07641_/A _07645_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07635_/B sky130_fd_sc_hd__nand3_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05909_ _05909_/A _05909_/B vssd1 vssd1 vccd1 vccd1 _05909_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09811_/B _09677_/B _09676_/X vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__or3b_1
XFILLER_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05912__B _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08628_ _10792_/Q _10791_/Q _08628_/C vssd1 vssd1 vccd1 vccd1 _08642_/D sky130_fd_sc_hd__and3_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06889_ _06886_/A _06886_/B _06891_/A _06891_/B vssd1 vssd1 vccd1 vccd1 _06890_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08559_ _10773_/Q _08559_/B vssd1 vssd1 vccd1 vccd1 _08559_/X sky130_fd_sc_hd__and2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10451__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10521_ _06124_/X _10522_/A _10520_/X _05983_/X vssd1 vssd1 vccd1 vccd1 _10979_/D
+ sky130_fd_sc_hd__a211o_2
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08016__A _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10452_ _10954_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__or2_1
XFILLER_124_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10383_ _10934_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__and2_1
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08686__A _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09281__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06918__B _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10719_ _10737_/CLK _10719_/D vssd1 vssd1 vccd1 vccd1 _10719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07843__C1 _07842_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07930_ input8/X vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__inv_2
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07861_ _07848_/X _05460_/D _07844_/X hold10/X vssd1 vssd1 vccd1 vccd1 _10628_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06812_ _06805_/A _06805_/B _06293_/A vssd1 vssd1 vccd1 vccd1 _06813_/B sky130_fd_sc_hd__a21oi_2
X_07792_ _07792_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__xnor2_1
X_09600_ _09600_/A _09653_/A vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__or2_1
XFILLER_95_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09531_ hold11/A _09408_/X _09529_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10871_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06743_ _06752_/B _06743_/B vssd1 vssd1 vccd1 vccd1 _06774_/B sky130_fd_sc_hd__xnor2_2
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06674_ _06674_/A _06681_/A _06674_/C vssd1 vssd1 vccd1 vccd1 _06678_/A sky130_fd_sc_hd__nand3_1
XFILLER_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09462_ _09462_/A _09462_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__and3_1
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05625_ _10549_/Q _05630_/A _10550_/Q vssd1 vssd1 vccd1 vccd1 _05626_/B sky130_fd_sc_hd__o21ai_1
X_08413_ _10495_/A vssd1 vssd1 vccd1 vccd1 _10394_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09393_ _09430_/A _09393_/B vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__nor2_2
X_08344_ _08263_/X _08350_/B _08340_/Y _08343_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08344_/X sky130_fd_sc_hd__o311a_1
X_05556_ _10559_/Q _10558_/Q _05610_/A vssd1 vssd1 vccd1 vccd1 _05604_/A sky130_fd_sc_hd__or3_1
XANTENNA__06844__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08275_ _08277_/A vssd1 vssd1 vccd1 vccd1 _08278_/A sky130_fd_sc_hd__clkbuf_2
X_05487_ _05487_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05487_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07834__C1 _07833_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07226_ _07235_/C _07142_/B _07224_/X _07223_/X _07217_/Y vssd1 vssd1 vccd1 vccd1
+ _07227_/B sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_41_clock _10704_/CLK vssd1 vssd1 vccd1 vccd1 _10865_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_118_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07157_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07282_/A sky130_fd_sc_hd__xor2_1
X_06108_ _10704_/Q _08297_/B vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__or2_1
XANTENNA__07675__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07088_ _07089_/A _07089_/B vssd1 vssd1 vccd1 vccd1 _07359_/A sky130_fd_sc_hd__and2_1
X_06039_ _06039_/A vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_56_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10968_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__09400__A_N _09399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05915__A2 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ _09647_/A _09647_/B _09728_/X vssd1 vssd1 vccd1 vccd1 _09730_/B sky130_fd_sc_hd__a21oi_1
XFILLER_47_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ _10504_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10504_/X sky130_fd_sc_hd__or2_1
XFILLER_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09042__A1 _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ _06124_/X _10431_/X _10434_/X _08563_/X vssd1 vssd1 vccd1 vccd1 _10947_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10188__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_7_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 _10704_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10495_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10427_/B sky130_fd_sc_hd__nand2_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10297_ _10297_/A vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__inv_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05833__A _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05410_ _05408_/Y _10616_/Q _05480_/A _08994_/A vssd1 vssd1 vccd1 vccd1 _05410_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06390_ _06502_/C vssd1 vssd1 vccd1 vccd1 _06489_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__07816__C1 _07815_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05341_ _10638_/Q vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08060_ _08352_/B vssd1 vssd1 vccd1 vccd1 _08061_/A sky130_fd_sc_hd__buf_2
XFILLER_119_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05272_ _10657_/Q vssd1 vssd1 vccd1 vccd1 _06039_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07011_ _07567_/A _07433_/A vssd1 vssd1 vccd1 vccd1 _07472_/A sky130_fd_sc_hd__and2_1
XFILLER_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08962_ _10947_/Q _10430_/B _08961_/X vssd1 vssd1 vccd1 vccd1 _08962_/Y sky130_fd_sc_hd__a21oi_1
X_07913_ _07916_/A _07913_/B vssd1 vssd1 vccd1 vccd1 _10642_/D sky130_fd_sc_hd__nor2_1
X_08893_ _08889_/X _08890_/X _08891_/X _08892_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08893_/X sky130_fd_sc_hd__o311a_1
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07844_ _08557_/A vssd1 vssd1 vccd1 vccd1 _07844_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07775_ _07773_/Y _07773_/B _07775_/S vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09514_ _09514_/A _09514_/B _09514_/C vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__nand3_1
X_06726_ _07796_/A _06726_/B vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__or2_1
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06657_ _06657_/A _06657_/B vssd1 vssd1 vccd1 vccd1 _06658_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09445_ _09676_/B _09445_/B vssd1 vssd1 vccd1 vccd1 _09448_/A sky130_fd_sc_hd__xor2_4
X_05608_ _10696_/Q vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10406__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09376_ _09376_/A vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__inv_2
X_06588_ _06576_/B _06587_/C _06587_/B vssd1 vssd1 vccd1 vccd1 _06589_/B sky130_fd_sc_hd__a21oi_1
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08327_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08339_/C sky130_fd_sc_hd__and2_1
X_05539_ _10541_/Q vssd1 vssd1 vccd1 vccd1 _05539_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10096__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ _08258_/A vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__buf_2
XANTENNA__06086__B2 _06066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09024__A1 _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07209_ _07280_/C _07209_/B vssd1 vssd1 vccd1 vccd1 _07279_/B sky130_fd_sc_hd__or2_1
X_08189_ _08191_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08189_/X sky130_fd_sc_hd__or2_1
XFILLER_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10220_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10220_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10151_ _10151_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__xnor2_1
XFILLER_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08013__B _08021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _10126_/A _10082_/B vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__and2_1
XFILLER_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10342__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08838__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10984_ _10984_/CLK _10984_/D vssd1 vssd1 vccd1 vccd1 _10984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05521__B1 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07813__A2 _10616_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10418_ _10943_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__and2_1
XFILLER_97_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _09312_/X _06371_/C _10346_/X _10918_/Q vssd1 vssd1 vccd1 vccd1 _10918_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07329__A1 _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05890_ _10658_/Q _05895_/A vssd1 vssd1 vccd1 vccd1 _05891_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06001__A1 _07849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07560_ _07560_/A vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06511_ _06511_/A _06511_/B vssd1 vssd1 vccd1 vccd1 _06512_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ _10441_/A vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07491_ _07509_/A _07509_/B vssd1 vssd1 vccd1 vccd1 _07510_/A sky130_fd_sc_hd__nor2_1
X_06442_ _06442_/A _06442_/B vssd1 vssd1 vccd1 vccd1 _06469_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _10810_/Q _08985_/X _08988_/X _10723_/Q _09160_/X vssd1 vssd1 vccd1 vccd1
+ _09161_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06373_ _06305_/A _06274_/B _06262_/A vssd1 vssd1 vccd1 vccd1 _06374_/A sky130_fd_sc_hd__o21ai_2
X_08112_ _08112_/A vssd1 vssd1 vccd1 vccd1 _10685_/D sky130_fd_sc_hd__clkbuf_1
X_05324_ _05827_/A _05324_/B vssd1 vssd1 vccd1 vccd1 _05324_/X sky130_fd_sc_hd__and2_1
XANTENNA__06068__B2 _06066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09092_ _09092_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09118_/A sky130_fd_sc_hd__or2_1
XFILLER_30_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08043_ _08043_/A vssd1 vssd1 vccd1 vccd1 _08044_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__05815__A1 _05405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08114__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09994_ _10123_/A vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__inv_2
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08945_ _09124_/C _09142_/D vssd1 vssd1 vccd1 vccd1 _08968_/A sky130_fd_sc_hd__or2_1
XFILLER_130_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08876_ _08876_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _08876_/Y sky130_fd_sc_hd__nor2_1
X_07827_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07827_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06288__B _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07758_ _07758_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _10117_/A sky130_fd_sc_hd__xnor2_4
XFILLER_72_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06709_ _06717_/A _06717_/B vssd1 vssd1 vccd1 vccd1 _06711_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07689_ _07689_/A _09441_/A vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__or2b_1
X_09428_ _09454_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09460_/B sky130_fd_sc_hd__xor2_2
XFILLER_100_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09359_ _09359_/A vssd1 vssd1 vccd1 vccd1 _09361_/A sky130_fd_sc_hd__inv_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10203_ _10949_/Q _10933_/Q vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__or2b_1
XANTENNA_input41_A io_wbs_m2s_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10134_ _10134_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08959__A _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10065_ _09924_/B _10065_/B _10065_/C _10065_/D vssd1 vssd1 vccd1 vccd1 _10131_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_54_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08694__A _08819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10967_ _10968_/CLK _10967_/D vssd1 vssd1 vccd1 vccd1 _10967_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _10982_/CLK _10898_/D vssd1 vssd1 vccd1 vccd1 _10898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06222__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _07166_/A vssd1 vssd1 vccd1 vccd1 _07021_/A sky130_fd_sc_hd__clkbuf_2
X_05942_ _05838_/B _05941_/Y _05803_/A vssd1 vssd1 vccd1 vccd1 _05942_/X sky130_fd_sc_hd__a21o_1
X_08730_ _06163_/X _08728_/X _08729_/X _10805_/Q vssd1 vssd1 vccd1 vccd1 _08730_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05873_ _10660_/Q vssd1 vssd1 vccd1 vccd1 _05883_/A sky130_fd_sc_hd__buf_2
X_08661_ _08661_/A _08671_/A vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__or2_2
XFILLER_78_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07612_ _07539_/A _07505_/A _07505_/B _07536_/X _07611_/Y vssd1 vssd1 vccd1 vccd1
+ _07613_/A sky130_fd_sc_hd__a41o_1
X_08592_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07543_ _07543_/A _07753_/A vssd1 vssd1 vccd1 vccd1 _07544_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07474_ _07747_/B _07474_/B vssd1 vssd1 vccd1 vccd1 _07475_/C sky130_fd_sc_hd__nand2_1
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08109__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09213_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09296_/S sky130_fd_sc_hd__buf_2
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06425_ _06425_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06425_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07013__A _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _10957_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09144_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06356_ _10978_/Q _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06451_/C sky130_fd_sc_hd__and3_1
XFILLER_108_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05307_ _10669_/Q _05347_/B vssd1 vssd1 vccd1 vccd1 _05854_/A sky130_fd_sc_hd__or2_2
X_09075_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09297_/S sky130_fd_sc_hd__buf_4
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06287_ _06287_/A _06287_/B vssd1 vssd1 vccd1 vccd1 _06371_/C sky130_fd_sc_hd__nor2_2
XFILLER_135_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08026_ input35/X _08015_/X _08025_/X _08019_/X vssd1 vssd1 vccd1 vccd1 _10675_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07961__A1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09977_ _09977_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _10095_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08928_ _10830_/Q _08928_/B vssd1 vssd1 vccd1 vccd1 _08928_/X sky130_fd_sc_hd__xor2_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08859_ _08845_/Y _08870_/B _08858_/X vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__a21o_1
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10821_ _10823_/CLK _10821_/D vssd1 vssd1 vccd1 vccd1 _10821_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09403__A _09403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _10791_/CLK _10752_/D vssd1 vssd1 vccd1 vccd1 _10752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08019__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10683_ _10839_/CLK _10683_/D vssd1 vssd1 vccd1 vccd1 _10683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10117_ _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__xor2_1
X_10048_ _09980_/A _09980_/B _09975_/A vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06002__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06210_ _09104_/B vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07190_ _07190_/A _07190_/B vssd1 vssd1 vccd1 vccd1 _07277_/A sky130_fd_sc_hd__or2_1
XFILLER_117_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06141_ _06008_/X _06131_/X _06140_/Y _06137_/X vssd1 vssd1 vccd1 vccd1 _10585_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06072_ _10658_/Q vssd1 vssd1 vccd1 vccd1 _07979_/A sky130_fd_sc_hd__buf_2
XFILLER_132_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09900_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09915_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08599__A _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09831_ _09908_/A _09828_/B _09830_/X vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__a21o_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09762_ _09971_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09763_/C sky130_fd_sc_hd__xor2_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _10983_/Q vssd1 vssd1 vccd1 vccd1 _07086_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05925_ _05892_/X _05924_/X _05889_/X _08169_/A vssd1 vssd1 vccd1 vccd1 _05925_/X
+ sky130_fd_sc_hd__o22a_1
X_08713_ _08732_/B vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09693_ _09904_/A _09947_/B _09828_/B _10057_/A vssd1 vssd1 vccd1 vccd1 _09693_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05856_ _10669_/Q vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_81_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08644_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__buf_4
XFILLER_54_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05787_ _05787_/A _05787_/B vssd1 vssd1 vccd1 vccd1 _05802_/A sky130_fd_sc_hd__nand2_2
XANTENNA__09223__A _09228_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08575_ _08575_/A vssd1 vssd1 vccd1 vccd1 _10777_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10369__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _07526_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__xor2_1
XFILLER_23_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07457_ _07394_/X _07327_/X _07378_/Y vssd1 vssd1 vccd1 vccd1 _07493_/A sky130_fd_sc_hd__a21o_1
XFILLER_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06408_ _06626_/A _06408_/B _06408_/C vssd1 vssd1 vccd1 vccd1 _06645_/A sky130_fd_sc_hd__and3_1
X_07388_ _07456_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07454_/C sky130_fd_sc_hd__nor2_1
XANTENNA__07678__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__buf_2
X_06339_ _06575_/B vssd1 vssd1 vccd1 vccd1 _06459_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ _09834_/B vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__clkbuf_2
X_08009_ _08009_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08009_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08021__B _08021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10804_ _10806_/CLK _10804_/D vssd1 vssd1 vccd1 vccd1 _10804_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10735_ _10768_/CLK _10735_/D vssd1 vssd1 vccd1 vccd1 _10735_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08662__A2 _08819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05476__A2 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ _10666_/CLK _10666_/D vssd1 vssd1 vccd1 vccd1 _10666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10597_ _10878_/CLK _10597_/D vssd1 vssd1 vccd1 vccd1 _10597_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10221__A2 _10115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput80 _10865_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[31] sky130_fd_sc_hd__buf_2
XFILLER_110_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05710_ _08148_/A vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06690_ _06690_/A _06690_/B vssd1 vssd1 vccd1 vccd1 _06691_/B sky130_fd_sc_hd__or2_1
X_05641_ _05641_/A _05641_/B vssd1 vssd1 vccd1 vccd1 _05641_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08360_ _05528_/A _06011_/A _08037_/A _06115_/B _06024_/A vssd1 vssd1 vccd1 vccd1
+ _08360_/X sky130_fd_sc_hd__a41o_1
XFILLER_64_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05572_ _10708_/Q vssd1 vssd1 vccd1 vccd1 _08339_/B sky130_fd_sc_hd__clkbuf_2
X_07311_ _07312_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07313_/A sky130_fd_sc_hd__nor2_1
X_08291_ _08263_/X _08296_/B _08287_/Y _08290_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08291_/X sky130_fd_sc_hd__o311a_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07242_ _07242_/A _07242_/B vssd1 vssd1 vccd1 vccd1 _07246_/B sky130_fd_sc_hd__xnor2_1
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07173_ _07184_/A _07185_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07175_/B sky130_fd_sc_hd__o21bai_1
X_06124_ _06124_/A vssd1 vssd1 vccd1 vccd1 _06124_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06055_ _08173_/A _07981_/A _06050_/X _09104_/A _06054_/X vssd1 vssd1 vccd1 vccd1
+ _06071_/C sky130_fd_sc_hd__a221o_1
XFILLER_113_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_09814_ _09825_/B _09814_/B vssd1 vssd1 vccd1 vccd1 _09815_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09745_ _10493_/A _09810_/A _09745_/C vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__and3_1
X_06957_ _07651_/A _07659_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__nor3_1
X_05908_ _05908_/A _05908_/B vssd1 vssd1 vccd1 vccd1 _05909_/B sky130_fd_sc_hd__nor2_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09676_/A _09676_/B _09676_/C _09676_/D vssd1 vssd1 vccd1 vccd1 _09676_/X
+ sky130_fd_sc_hd__and4_1
X_06888_ _06872_/A _07801_/A _06873_/B vssd1 vssd1 vccd1 vccd1 _06891_/B sky130_fd_sc_hd__o21a_2
XANTENNA__08341__A1 _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05839_ _05831_/B _05831_/C _05838_/Y vssd1 vssd1 vccd1 vccd1 _05839_/X sky130_fd_sc_hd__o21a_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08627_ _08627_/A vssd1 vssd1 vccd1 vccd1 _10791_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06296__B _10905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08558_ _08558_/A vssd1 vssd1 vccd1 vccd1 _10772_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08489_ _08489_/A vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__buf_2
XFILLER_52_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07509_ _07509_/A _07509_/B vssd1 vssd1 vccd1 vccd1 _07510_/B sky130_fd_sc_hd__and2_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10520_ _10531_/B _09121_/X _07715_/C vssd1 vssd1 vccd1 vccd1 _10520_/X sky130_fd_sc_hd__o21a_1
XANTENNA__06655__B2 _06845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451_ _06163_/X _10446_/X _10450_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10953_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08016__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10382_ _10427_/B vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08032__A _08032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09109__B1 _09112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08868__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__B _08819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_3_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 _10840_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10718_ _10737_/CLK _10718_/D vssd1 vssd1 vccd1 vccd1 _10718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09310__B _09396_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08207__A _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10649_ _10832_/CLK _10649_/D vssd1 vssd1 vccd1 vccd1 _10649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07860_ _06193_/A _07849_/X _07850_/X _07859_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ hold10/A sky130_fd_sc_hd__o221ai_4
XFILLER_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07791_ _07791_/A _07791_/B vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__xnor2_1
X_06811_ _06851_/A _06811_/B vssd1 vssd1 vccd1 vccd1 _06813_/A sky130_fd_sc_hd__nand2_2
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _10043_/A vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__clkbuf_2
X_06742_ _06804_/A _06752_/C vssd1 vssd1 vccd1 vccd1 _06743_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09352__A_N _10906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06397__A _10977_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _09430_/A _09430_/B _09460_/X vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__a21o_1
XFILLER_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06673_ _06684_/A _06684_/B vssd1 vssd1 vccd1 vccd1 _06941_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05624_ _10689_/Q vssd1 vssd1 vccd1 vccd1 _08148_/A sky130_fd_sc_hd__clkbuf_2
X_08412_ _10432_/B vssd1 vssd1 vccd1 vccd1 _10495_/A sky130_fd_sc_hd__buf_2
XFILLER_24_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09392_ _09451_/B _09392_/B vssd1 vssd1 vccd1 vccd1 _09393_/B sky130_fd_sc_hd__and2_1
X_08343_ _08037_/A _08351_/B _08341_/Y _08342_/Y _08062_/A vssd1 vssd1 vccd1 vccd1
+ _08343_/X sky130_fd_sc_hd__a311o_1
X_05555_ _10557_/Q _05612_/A vssd1 vssd1 vccd1 vccd1 _05610_/A sky130_fd_sc_hd__or2_1
XFILLER_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08274_ input30/X vssd1 vssd1 vccd1 vccd1 _08274_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05486_ _05910_/B _05470_/B _05495_/A _05455_/X _05485_/Y vssd1 vssd1 vccd1 vccd1
+ _10544_/D sky130_fd_sc_hd__a221o_1
X_07225_ _07217_/Y _07223_/X _07224_/X _07142_/B _07186_/A vssd1 vssd1 vccd1 vccd1
+ _07225_/X sky130_fd_sc_hd__o2111a_1
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07156_ _07132_/A _07132_/B _07286_/A _07133_/A vssd1 vssd1 vccd1 vccd1 _07355_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06107_ _10703_/Q _10702_/Q _08278_/B vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__or3_1
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07087_ _07087_/A _07087_/B vssd1 vssd1 vccd1 vccd1 _07089_/B sky130_fd_sc_hd__nor2_1
X_06038_ _06038_/A vssd1 vssd1 vccd1 vccd1 _06038_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_120_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07989_ _06195_/X _07987_/X _07988_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10661_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09728_ _09665_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09728_/X sky130_fd_sc_hd__and2b_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _09716_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _09713_/B sky130_fd_sc_hd__and2_1
XFILLER_15_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10503_ _06008_/X _10496_/X _10502_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10972_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10434_ _10947_/Q _10440_/B vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__or2_1
XANTENNA__06770__A _07682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__A1 _07539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10365_ _10408_/A vssd1 vssd1 vccd1 vccd1 _10365_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10296_ _10958_/Q _10942_/Q vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__and2b_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09292__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05340_ _05340_/A _05340_/B vssd1 vssd1 vccd1 vccd1 _05340_/X sky130_fd_sc_hd__and2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05271_ _10662_/Q vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__inv_2
XFILLER_127_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_49_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__A1 _06997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ _07567_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07555_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06252__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08961_ _08948_/X _08953_/X _10474_/B _10478_/A vssd1 vssd1 vccd1 vccd1 _08961_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07912_ _10610_/Q _07906_/X _07910_/X _07911_/Y vssd1 vssd1 vccd1 vccd1 _07913_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08892_ _08890_/X _08891_/X _08889_/X vssd1 vssd1 vccd1 vccd1 _08892_/Y sky130_fd_sc_hd__o21ai_1
X_07843_ _07827_/X _05461_/D _07823_/X _07842_/Y vssd1 vssd1 vccd1 vccd1 _10624_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07774_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07775_/S sky130_fd_sc_hd__nor2_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ _09613_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09514_/C sky130_fd_sc_hd__nor2_1
X_06725_ _06725_/A _06725_/B vssd1 vssd1 vccd1 vccd1 _06726_/B sky130_fd_sc_hd__and2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06858__A1 _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06656_ _06656_/A _06656_/B vssd1 vssd1 vccd1 vccd1 _06660_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09444_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09445_/B sky130_fd_sc_hd__and2_1
X_05607_ _10697_/Q vssd1 vssd1 vccd1 vccd1 _08224_/A sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _10895_/Q _10911_/Q vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__and2b_1
XFILLER_40_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06587_ _06587_/A _06587_/B _06587_/C vssd1 vssd1 vccd1 vccd1 _06589_/A sky130_fd_sc_hd__and3_1
XFILLER_33_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08326_ _08025_/A _08058_/X _08325_/X vssd1 vssd1 vccd1 vccd1 _08326_/X sky130_fd_sc_hd__o21ba_1
X_05538_ _10542_/Q vssd1 vssd1 vccd1 vccd1 _05741_/B sky130_fd_sc_hd__inv_2
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06086__A2 _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08257_ _08267_/B _08253_/X _08254_/Y _08256_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08257_/X sky130_fd_sc_hd__a311o_1
X_05469_ _05472_/B vssd1 vssd1 vccd1 vccd1 _05470_/B sky130_fd_sc_hd__buf_2
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08188_ _08188_/A vssd1 vssd1 vccd1 vccd1 _08191_/A sky130_fd_sc_hd__buf_2
XFILLER_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07208_ _07208_/A _07208_/B vssd1 vssd1 vccd1 vccd1 _07209_/B sky130_fd_sc_hd__and2_1
XFILLER_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07139_ _07138_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _07139_/X sky130_fd_sc_hd__and2b_1
XFILLER_106_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10150_ _10478_/A _10068_/B _10070_/B _10074_/A vssd1 vssd1 vccd1 vccd1 _10151_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10081_ _10081_/A _10081_/B _10081_/C vssd1 vssd1 vccd1 vccd1 _10082_/B sky130_fd_sc_hd__or3_1
XFILLER_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09406__A _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08310__A _08837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10983_ _10986_/CLK _10983_/D vssd1 vssd1 vccd1 vccd1 _10983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09141__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06077__A2 _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10417_ _10408_/X _10723_/Q _10414_/X _10416_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10942_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06005__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _09634_/A _06352_/A _10192_/X _10917_/Q vssd1 vssd1 vccd1 vccd1 _10917_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_112_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10279_ _10277_/X _10278_/Y _10279_/S vssd1 vssd1 vccd1 vccd1 _10279_/X sky130_fd_sc_hd__mux2_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09316__A _09316_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06510_ _06510_/A _06510_/B vssd1 vssd1 vccd1 vccd1 _06511_/B sky130_fd_sc_hd__or2_1
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07490_ _07490_/A _07490_/B vssd1 vssd1 vccd1 vccd1 _07509_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_06441_ _06461_/B _06441_/B _06547_/C _06567_/B vssd1 vssd1 vccd1 vccd1 _06442_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09160_ _07981_/A _09123_/X _09127_/X _09159_/X vssd1 vssd1 vccd1 vccd1 _09160_/X
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_55_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10958_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06372_ _06804_/A _06387_/A vssd1 vssd1 vccd1 vccd1 _06375_/A sky130_fd_sc_hd__nand2_2
X_08111_ _08111_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__and2_1
X_05323_ _05830_/A _05831_/B _08342_/A vssd1 vssd1 vccd1 vccd1 _05324_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06068__A2 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09091_ _07393_/Y _08965_/Y _09209_/B vssd1 vssd1 vccd1 vccd1 _09112_/A sky130_fd_sc_hd__a21oi_4
XFILLER_30_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08042_ _08062_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__nor2_2
XANTENNA__05815__A2 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__xor2_2
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ _08944_/A vssd1 vssd1 vccd1 vccd1 _09124_/A sky130_fd_sc_hd__buf_2
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08875_ _10823_/Q vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07826_ _06255_/X _05453_/A _07823_/X _07825_/Y vssd1 vssd1 vccd1 vccd1 _10620_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07757_ _07757_/A _07757_/B vssd1 vssd1 vccd1 vccd1 _07758_/B sky130_fd_sc_hd__xor2_2
XFILLER_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06708_ _06630_/A _06631_/A _06630_/B vssd1 vssd1 vccd1 vccd1 _06717_/B sky130_fd_sc_hd__o21ba_1
XFILLER_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07688_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__xnor2_1
X_09427_ _09427_/A _09427_/B vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__xor2_4
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06639_ _06715_/A _06639_/B vssd1 vssd1 vccd1 vccd1 _06641_/C sky130_fd_sc_hd__and2_1
XFILLER_25_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09358_ _10886_/Q _10902_/Q vssd1 vssd1 vccd1 vccd1 _09359_/A sky130_fd_sc_hd__or2b_1
X_08309_ _08305_/A _08315_/C _08308_/Y vssd1 vssd1 vccd1 vccd1 _08309_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06059__A2 _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09289_ _09289_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__and2_1
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ _10933_/Q _10949_/Q vssd1 vssd1 vccd1 vccd1 _10202_/X sky130_fd_sc_hd__or2b_1
XFILLER_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10133_ _10133_/A _10133_/B vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input34_A io_wbs_m2s_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09136__A _09136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10064_ _10064_/A _10064_/B vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09181__A1 _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10966_ _10968_/CLK _10966_/D vssd1 vssd1 vccd1 vccd1 _10966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10897_ _10909_/CLK _10897_/D vssd1 vssd1 vccd1 vccd1 _10897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05574__A _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10480__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07166_/A sky130_fd_sc_hd__clkbuf_2
X_05941_ _08318_/A _05941_/B vssd1 vssd1 vccd1 vccd1 _05941_/Y sky130_fd_sc_hd__nand2_1
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09046__A _09930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05872_ _05872_/A _05872_/B vssd1 vssd1 vccd1 vccd1 _05872_/X sky130_fd_sc_hd__and2_1
X_08660_ _10369_/A _08971_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08671_/A sky130_fd_sc_hd__and3_1
XANTENNA__09172__B2 _10724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07611_ _07622_/A _07536_/X _07505_/X vssd1 vssd1 vccd1 vccd1 _07611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08591_ input51/X _10253_/A vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__or2_1
XFILLER_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07542_ _07402_/A _07402_/B _07405_/A vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__a21oi_1
X_07473_ _07473_/A _07473_/B vssd1 vssd1 vccd1 vccd1 _07477_/B sky130_fd_sc_hd__and2_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09212_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06424_ _06426_/A _06441_/B _06489_/B _06540_/A vssd1 vssd1 vccd1 vccd1 _06425_/B
+ sky130_fd_sc_hd__and4_1
X_09143_ _10432_/A _09143_/B vssd1 vssd1 vccd1 vccd1 _09143_/Y sky130_fd_sc_hd__nor2_1
X_06355_ _06550_/C vssd1 vssd1 vccd1 vccd1 _06554_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05306_ _10668_/Q _10667_/Q _05350_/B vssd1 vssd1 vccd1 vccd1 _05347_/B sky130_fd_sc_hd__or3_1
XFILLER_135_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08125__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _09067_/X _09073_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10839_/D sky130_fd_sc_hd__o21a_2
X_06286_ _06270_/A _06276_/A _06284_/X _06272_/Y vssd1 vssd1 vccd1 vccd1 _06287_/B
+ sky130_fd_sc_hd__a211oi_1
X_08025_ _08025_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or2_1
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08199__C1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08738__A1 _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09976_ _09977_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _09976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08927_ _08927_/A _08927_/B _08927_/C vssd1 vssd1 vccd1 vccd1 _08927_/X sky130_fd_sc_hd__or3_1
XFILLER_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08858_ _10820_/Q _08847_/X _08919_/B vssd1 vssd1 vccd1 vccd1 _08858_/X sky130_fd_sc_hd__o21a_1
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07809_ hold16/X _07824_/B vssd1 vssd1 vccd1 vccd1 _07809_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08789_ _10813_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08803_/C sky130_fd_sc_hd__xor2_1
XFILLER_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10820_ _10826_/CLK _10820_/D vssd1 vssd1 vccd1 vccd1 _10820_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09403__B _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _10791_/CLK _10751_/D vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10682_ _10682_/CLK _10682_/D vssd1 vssd1 vccd1 vccd1 _10682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07874__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10536__A1 _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10116_ _10109_/A _10109_/B _09626_/A vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__o21ai_1
X_10047_ _09970_/A _09970_/B _09983_/B _09982_/B _09982_/A vssd1 vssd1 vccd1 vccd1
+ _10051_/A sky130_fd_sc_hd__o32a_1
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10949_ _10978_/CLK _10949_/D vssd1 vssd1 vccd1 vccd1 _10949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10348__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06140_ _06140_/A _06145_/B vssd1 vssd1 vccd1 vccd1 _06140_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10194__B _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06071_ _06071_/A _06071_/B _06071_/C _06071_/D vssd1 vssd1 vccd1 vccd1 _06071_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_132_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07784__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08599__B _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__A1 _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09830_ _09977_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09830_/X sky130_fd_sc_hd__and2_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09761_ _09647_/A _09834_/A _09761_/C vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__and3b_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _07622_/A vssd1 vssd1 vccd1 vccd1 _07539_/A sky130_fd_sc_hd__buf_2
X_05924_ _10690_/Q _05892_/B _05895_/X _08146_/A _05923_/X vssd1 vssd1 vccd1 vccd1
+ _05924_/X sky130_fd_sc_hd__o221a_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08712_ _08688_/X _08710_/Y _08711_/X vssd1 vssd1 vccd1 vccd1 _10804_/D sky130_fd_sc_hd__o21a_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09692_ _09692_/A vssd1 vssd1 vccd1 vccd1 _09947_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05855_ _08013_/A _05858_/B _05852_/B vssd1 vssd1 vccd1 vccd1 _05935_/B sky130_fd_sc_hd__o21a_1
XFILLER_82_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08643_ _10796_/Q _08686_/A _08643_/C vssd1 vssd1 vccd1 vccd1 _08648_/B sky130_fd_sc_hd__and3_1
XFILLER_66_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05786_ _05768_/X _05770_/X _05786_/C _05786_/D vssd1 vssd1 vccd1 vccd1 _05787_/B
+ sky130_fd_sc_hd__and4bb_1
X_08574_ _08580_/B _08574_/B _08576_/B vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__and3_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07525_ _07525_/A _07525_/B vssd1 vssd1 vccd1 vccd1 _07526_/B sky130_fd_sc_hd__nand2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07959__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07456_ _07456_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07499_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07387_ _07391_/A _07459_/B _07748_/B _07378_/Y _07397_/A vssd1 vssd1 vccd1 vccd1
+ _07456_/B sky130_fd_sc_hd__a41o_1
X_06407_ _06630_/A _06407_/B vssd1 vssd1 vccd1 vccd1 _06408_/C sky130_fd_sc_hd__xor2_1
XFILLER_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09126_ _09126_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09270_/A sky130_fd_sc_hd__and2_2
X_06338_ _06338_/A vssd1 vssd1 vccd1 vccd1 _06575_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09057_ _10967_/Q vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06269_ _10917_/Q _10900_/Q vssd1 vssd1 vccd1 vccd1 _06270_/B sky130_fd_sc_hd__or2_1
XFILLER_123_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08008_ _08256_/A vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__inv_2
XFILLER_2_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09959_ _09959_/A _09958_/A vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__or2b_1
XANTENNA__05945__A1 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08344__C1 _08258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08895__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10803_ _10803_/CLK _10803_/D vssd1 vssd1 vccd1 vccd1 _10803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10734_ _10768_/CLK _10734_/D vssd1 vssd1 vccd1 vccd1 _10734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10665_ _10811_/CLK _10665_/D vssd1 vssd1 vccd1 vccd1 _10665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10596_ _10958_/CLK _10596_/D vssd1 vssd1 vccd1 vccd1 _10596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10509__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput70 _10856_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput81 _10837_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_122_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05852__A _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05640_ _05910_/B _10543_/Q vssd1 vssd1 vccd1 vccd1 _05641_/B sky130_fd_sc_hd__xnor2_1
XFILLER_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05571_ _10570_/Q _05576_/A vssd1 vssd1 vccd1 vccd1 _05571_/X sky130_fd_sc_hd__xor2_1
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07310_ _07310_/A _07310_/B vssd1 vssd1 vccd1 vccd1 _07312_/B sky130_fd_sc_hd__or2_1
X_08290_ _08297_/B _08253_/X _08288_/Y _08289_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08290_/X sky130_fd_sc_hd__a311o_1
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07241_ _07250_/A _07217_/B _07218_/X vssd1 vssd1 vccd1 vccd1 _07242_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09994__A _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07172_ _07192_/B _07192_/A vssd1 vssd1 vccd1 vccd1 _07185_/A sky130_fd_sc_hd__and2b_1
XFILLER_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06123_ input16/X vssd1 vssd1 vccd1 vccd1 _06124_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_105_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06054_ _05744_/Y _07998_/A _05883_/A _08181_/A _06053_/X vssd1 vssd1 vccd1 vccd1
+ _06054_/X sky130_fd_sc_hd__a221o_1
XFILLER_105_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09813_ _09743_/A _09743_/B _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09814_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_113_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09744_ _09744_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09745_/C sky130_fd_sc_hd__nand2_1
X_06956_ _07663_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__nand2_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05907_ _05907_/A vssd1 vssd1 vccd1 vccd1 _05908_/A sky130_fd_sc_hd__inv_2
XFILLER_100_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09675_ _09733_/B _09675_/B vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06887_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _07801_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05838_ _08025_/A _05838_/B vssd1 vssd1 vccd1 vccd1 _05838_/Y sky130_fd_sc_hd__nand2_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08626_ _08631_/C _08649_/A _08626_/C vssd1 vssd1 vccd1 vccd1 _08627_/A sky130_fd_sc_hd__and3b_1
XFILLER_55_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05769_ _05769_/A vssd1 vssd1 vccd1 vccd1 _05769_/Y sky130_fd_sc_hd__inv_2
X_08557_ _08557_/A _08557_/B _08557_/C vssd1 vssd1 vccd1 vccd1 _08558_/A sky130_fd_sc_hd__and3_1
XFILLER_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08488_ _08488_/A vssd1 vssd1 vccd1 vccd1 _10745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07508_ _07508_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07628_/A sky130_fd_sc_hd__xnor2_2
XFILLER_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07439_ _07439_/A vssd1 vssd1 vccd1 vccd1 _07732_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10450_ _10953_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__or2_1
XFILLER_10_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ _10806_/Q _09168_/A _09112_/A _09103_/Y _09108_/X vssd1 vssd1 vccd1 vccd1
+ _09110_/B sky130_fd_sc_hd__a221o_1
XFILLER_136_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10381_ _10365_/X _10714_/Q _10379_/X _10380_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10933_/D sky130_fd_sc_hd__o221a_1
XFILLER_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08313__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08032__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06040__B1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _10737_/CLK _10717_/D vssd1 vssd1 vccd1 vccd1 _10717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10648_ _10651_/CLK _10648_/D vssd1 vssd1 vccd1 vccd1 _10648_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06008__A _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10579_ _10833_/CLK _10579_/D vssd1 vssd1 vccd1 vccd1 _10579_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_6_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08020__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06810_ _10928_/Q _07570_/A vssd1 vssd1 vccd1 vccd1 _06811_/B sky130_fd_sc_hd__nand2_1
X_07790_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07791_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_45_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06741_ _06741_/A vssd1 vssd1 vccd1 vccd1 _06834_/A sky130_fd_sc_hd__inv_2
X_09460_ _09429_/A _09460_/B vssd1 vssd1 vccd1 vccd1 _09460_/X sky130_fd_sc_hd__and2b_1
X_08411_ _08419_/A _10745_/Q _08992_/A _08410_/X vssd1 vssd1 vccd1 vccd1 _10727_/D
+ sky130_fd_sc_hd__o211a_1
X_06672_ _06672_/A _06672_/B vssd1 vssd1 vccd1 vccd1 _06684_/B sky130_fd_sc_hd__xor2_1
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05623_ _05623_/A _05623_/B vssd1 vssd1 vccd1 vccd1 _05623_/X sky130_fd_sc_hd__and2_1
X_09391_ _09451_/B _09392_/B vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__nor2_2
X_08342_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08342_/Y sky130_fd_sc_hd__nor2_1
X_05554_ _10556_/Q _10555_/Q _05663_/A _05663_/B vssd1 vssd1 vccd1 vccd1 _05612_/A
+ sky130_fd_sc_hd__or4_1
X_08273_ _08273_/A vssd1 vssd1 vccd1 vccd1 _10701_/D sky130_fd_sc_hd__clkbuf_1
X_05485_ _05485_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05485_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07224_ _10981_/Q _07235_/B vssd1 vssd1 vccd1 vccd1 _07224_/X sky130_fd_sc_hd__and2_1
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07155_ _07285_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07286_/A sky130_fd_sc_hd__nor2_1
X_06106_ _10701_/Q _08267_/B vssd1 vssd1 vccd1 vccd1 _08278_/B sky130_fd_sc_hd__or2_1
XFILLER_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09229__A _09229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ _07326_/A _07086_/B _07188_/B _07178_/A vssd1 vssd1 vccd1 vccd1 _07087_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_133_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06037_ _06037_/A vssd1 vssd1 vccd1 vccd1 _08105_/A sky130_fd_sc_hd__clkinv_2
XFILLER_99_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07988_ _07988_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07988_/X sky130_fd_sc_hd__or2_1
XFILLER_59_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09727_ _09727_/A _09727_/B vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06939_ _06939_/A _06939_/B vssd1 vssd1 vccd1 vccd1 _07630_/A sky130_fd_sc_hd__xor2_4
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ _09760_/B vssd1 vssd1 vccd1 vccd1 _09977_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08609_ _08609_/A vssd1 vssd1 vccd1 vccd1 _10786_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09639_/B _09536_/B _09486_/A _09588_/X vssd1 vssd1 vccd1 vccd1 _09590_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07212__A _07415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08027__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10502_ _10502_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10502_/X sky130_fd_sc_hd__or2_1
XFILLER_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10433_ _10472_/B vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10188__A2 _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08250__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10364_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10408_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08043__A _08043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10295_ _10942_/Q _10958_/Q vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__or2b_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08069__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05270_ _10678_/Q vssd1 vssd1 vccd1 vccd1 _08352_/A sky130_fd_sc_hd__buf_2
XFILLER_128_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09018__A0 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08960_ _10068_/A vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__clkbuf_4
X_07911_ _07911_/A vssd1 vssd1 vccd1 vccd1 _07911_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__06004__A0 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08891_ _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08891_/X sky130_fd_sc_hd__and2_1
X_07842_ hold5/X _07828_/X _07829_/X _07841_/Y _07832_/X vssd1 vssd1 vccd1 vccd1 _07842_/Y
+ sky130_fd_sc_hd__o221ai_4
XANTENNA__09741__B2 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__A1 _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07773_ _10508_/A _07773_/B vssd1 vssd1 vccd1 vccd1 _07773_/Y sky130_fd_sc_hd__nand2_1
X_09512_ _10069_/A _09692_/A _09761_/C _09736_/B vssd1 vssd1 vccd1 vccd1 _09513_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_71_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06724_ _06725_/A _06725_/B vssd1 vssd1 vccd1 vccd1 _07796_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09443_ _10967_/Q _09443_/B vssd1 vssd1 vccd1 vccd1 _09534_/C sky130_fd_sc_hd__nand2_1
X_06655_ _06800_/A _06408_/B _06428_/B _06845_/A vssd1 vssd1 vccd1 vccd1 _06656_/B
+ sky130_fd_sc_hd__a22oi_1
X_05606_ _10558_/Q _05610_/A vssd1 vssd1 vccd1 vccd1 _05606_/X sky130_fd_sc_hd__xor2_1
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09374_ _09923_/A _09674_/B _09372_/X _09373_/Y vssd1 vssd1 vccd1 vccd1 _09922_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08325_ _08332_/B _08058_/A _08324_/Y _08120_/X vssd1 vssd1 vccd1 vccd1 _08325_/X
+ sky130_fd_sc_hd__a31o_1
X_06586_ _06591_/A _06591_/B vssd1 vssd1 vccd1 vccd1 _06949_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05537_ _10543_/Q vssd1 vssd1 vccd1 vccd1 _05737_/B sky130_fd_sc_hd__inv_2
X_08256_ _08256_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05468_ _05453_/X _05459_/X _05460_/X _05462_/X _05467_/X vssd1 vssd1 vccd1 vccd1
+ _05472_/B sky130_fd_sc_hd__a2111oi_1
XFILLER_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08187_ _08188_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08196_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07207_ _07208_/A _07208_/B vssd1 vssd1 vccd1 vccd1 _07280_/C sky130_fd_sc_hd__nor2_1
XFILLER_134_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05399_ _10651_/Q _10575_/Q vssd1 vssd1 vccd1 vccd1 _05400_/B sky130_fd_sc_hd__xnor2_1
XFILLER_106_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07138_ _07138_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _07147_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07069_ _07149_/C _07186_/B _07312_/A vssd1 vssd1 vccd1 vccd1 _07070_/B sky130_fd_sc_hd__and3_1
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10080_ _10081_/A _10081_/B _10081_/C vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10982_ _10982_/CLK _10982_/D vssd1 vssd1 vccd1 vccd1 _10982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08038__A _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07877__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08223__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10416_ input18/X _10399_/X _10415_/X vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__a21bo_1
XFILLER_7_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10347_ _09312_/X _06281_/B _10346_/X _10916_/Q vssd1 vssd1 vccd1 vccd1 _10916_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08501__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ _10265_/A _10268_/Y _10265_/B vssd1 vssd1 vccd1 vccd1 _10278_/Y sky130_fd_sc_hd__o21bai_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09316__B _09337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06021__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10478__A _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06440_ _06440_/A vssd1 vssd1 vccd1 vccd1 _06567_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06371_ _06371_/A _06371_/B _06371_/C vssd1 vssd1 vccd1 vccd1 _06387_/A sky130_fd_sc_hd__or3_1
X_08110_ _10533_/A _08086_/X _08109_/X _05728_/X _08166_/A vssd1 vssd1 vccd1 vccd1
+ _08111_/B sky130_fd_sc_hd__o221a_1
X_05322_ _10677_/Q vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__buf_2
X_09090_ _09090_/A vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__clkbuf_2
X_08041_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09992_ _10480_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08943_ _10518_/B vssd1 vssd1 vccd1 vccd1 _08943_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05984__C1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08874_ _10823_/Q _08888_/B vssd1 vssd1 vccd1 vccd1 _08883_/A sky130_fd_sc_hd__and2_1
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09190__A2 _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ _06156_/A _06258_/X _07807_/X _07824_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07825_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_56_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07756_ _07756_/A _07756_/B vssd1 vssd1 vccd1 vccd1 _07757_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09242__A _09242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06707_ _06719_/B _07791_/A _06706_/X vssd1 vssd1 vccd1 vccd1 _06711_/A sky130_fd_sc_hd__o21a_1
XFILLER_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09426_ _10963_/Q _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09427_/B sky130_fd_sc_hd__and3_1
XFILLER_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07687_ _07687_/A _07687_/B vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06638_ _06638_/A _06638_/B vssd1 vssd1 vccd1 vccd1 _06639_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09357_ _10903_/Q _10887_/Q vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__or2b_1
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06569_ _06570_/A _06570_/B vssd1 vssd1 vccd1 vccd1 _06597_/B sky130_fd_sc_hd__nand2_1
X_08308_ _08305_/A _08315_/C _08092_/A vssd1 vssd1 vccd1 vccd1 _08308_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09288_ _10828_/Q _09274_/X _09275_/X _09287_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09289_/B sky130_fd_sc_hd__a32o_1
XFILLER_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08239_ input25/X _08212_/X _08124_/X _08233_/A _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08240_/B sky130_fd_sc_hd__o221a_1
XFILLER_20_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10201_ _07098_/A _10192_/X _10200_/X vssd1 vssd1 vccd1 vccd1 _10899_/D sky130_fd_sc_hd__a21o_1
X_10132_ _10480_/A _10068_/B _10131_/X _10068_/A vssd1 vssd1 vccd1 vccd1 _10133_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09417__A _09417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _10065_/C _10063_/B vssd1 vssd1 vccd1 vccd1 _10064_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09181__A2 _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input27_A io_wbs_m2s_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10965_ _10968_/CLK _10965_/D vssd1 vssd1 vccd1 vccd1 _10965_/Q sky130_fd_sc_hd__dfxtp_1
X_10896_ _10909_/CLK _10896_/D vssd1 vssd1 vccd1 vccd1 _10896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06016__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10003__B2 _09716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__A1 _09930_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05940_ _08315_/B _05940_/B vssd1 vssd1 vccd1 vccd1 _05940_/X sky130_fd_sc_hd__or2_1
XFILLER_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05871_ _05848_/B _05823_/A _06052_/A vssd1 vssd1 vccd1 vccd1 _05872_/B sky130_fd_sc_hd__o21ai_1
XFILLER_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08590_ _09403_/B vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__buf_2
X_07610_ _07610_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__xnor2_2
XFILLER_93_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07541_ _07410_/A _07410_/B _07540_/X vssd1 vssd1 vccd1 vccd1 _07546_/B sky130_fd_sc_hd__o21a_1
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07472_ _07472_/A _07472_/B vssd1 vssd1 vccd1 vccd1 _07473_/B sky130_fd_sc_hd__or2_1
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ _09211_/A _09211_/B vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__nor2_2
XANTENNA__10490__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06423_ _06426_/A _06627_/B _06540_/A _06441_/B vssd1 vssd1 vccd1 vccd1 _06425_/A
+ sky130_fd_sc_hd__a22oi_1
X_09142_ _09142_/A _09142_/B _09142_/C _09142_/D vssd1 vssd1 vccd1 vccd1 _09143_/B
+ sky130_fd_sc_hd__or4_1
X_06354_ _06352_/B _06352_/C _06352_/A vssd1 vssd1 vccd1 vccd1 _06550_/C sky130_fd_sc_hd__o21ai_1
X_05305_ _05353_/A vssd1 vssd1 vccd1 vccd1 _05350_/B sky130_fd_sc_hd__clkbuf_2
X_09073_ _10123_/A _10474_/B _10495_/B _10510_/A _09072_/X vssd1 vssd1 vccd1 vccd1
+ _09073_/X sky130_fd_sc_hd__a221o_1
X_06285_ _06284_/X _06272_/Y _06270_/A _06276_/A vssd1 vssd1 vccd1 vccd1 _06287_/A
+ sky130_fd_sc_hd__o211a_1
X_08024_ input34/X _08015_/X _08023_/Y _08019_/X vssd1 vssd1 vccd1 vccd1 _10674_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09975_ _09975_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__nor2_1
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08926_ _09153_/A _08926_/B vssd1 vssd1 vccd1 vccd1 _10829_/D sky130_fd_sc_hd__nor2_1
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08857_ _08866_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08870_/C sky130_fd_sc_hd__and2_1
XFILLER_85_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07808_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07824_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08788_ _08783_/Y _08784_/X _08787_/X vssd1 vssd1 vccd1 vccd1 _10812_/D sky130_fd_sc_hd__o21a_1
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07739_ _07739_/A _07739_/B vssd1 vssd1 vccd1 vccd1 _07740_/B sky130_fd_sc_hd__xnor2_1
X_10750_ _10791_/CLK _10750_/D vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
X_10681_ _10682_/CLK _10681_/D vssd1 vssd1 vccd1 vccd1 _10681_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10481__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09409_ _09409_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__xnor2_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07937__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08051__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10115_ _10115_/A vssd1 vssd1 vccd1 vccd1 _10115_/X sky130_fd_sc_hd__buf_2
XFILLER_0_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_54_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10813_/CLK sky130_fd_sc_hd__clkbuf_16
X_10046_ _10046_/A _09985_/A vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__or2b_1
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_69_clock _10985_/CLK vssd1 vssd1 vccd1 vccd1 _10984_/CLK sky130_fd_sc_hd__clkbuf_16
X_10948_ _10956_/CLK _10948_/D vssd1 vssd1 vccd1 vccd1 _10948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10879_ _10958_/CLK _10879_/D vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06070_ _06070_/A _06070_/B vssd1 vssd1 vccd1 vccd1 _06071_/D sky130_fd_sc_hd__nand2_1
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05585__A _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10491__A _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09760_ _09834_/B _09760_/B vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__and2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _07715_/D vssd1 vssd1 vccd1 vccd1 _07622_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05923_ _06035_/A _05897_/X _05895_/X _08148_/A _05922_/X vssd1 vssd1 vccd1 vccd1
+ _05923_/X sky130_fd_sc_hd__a221o_1
XFILLER_100_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08711_ _10533_/A _08694_/X _08695_/X _10804_/Q _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08711_/X sky130_fd_sc_hd__o221a_1
X_09691_ _09761_/C vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08642_ _10795_/Q _10794_/Q _10793_/Q _08642_/D vssd1 vssd1 vccd1 vccd1 _08643_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05854_ _05854_/A _05854_/B vssd1 vssd1 vccd1 vccd1 _05858_/B sky130_fd_sc_hd__nor2_1
XFILLER_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05785_ _05785_/A _05785_/B _05785_/C vssd1 vssd1 vccd1 vccd1 _05786_/D sky130_fd_sc_hd__and3_1
X_08573_ _08578_/C _08578_/D vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__nand2_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07524_ _07649_/A vssd1 vssd1 vccd1 vccd1 _07527_/B sky130_fd_sc_hd__inv_2
XFILLER_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07455_ _07455_/A _07455_/B vssd1 vssd1 vccd1 vccd1 _07502_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06406_ _06690_/A _06426_/A _06428_/B vssd1 vssd1 vccd1 vccd1 _06407_/B sky130_fd_sc_hd__and3b_1
XFILLER_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07386_ _07391_/A _07386_/B vssd1 vssd1 vccd1 vccd1 _07397_/A sky130_fd_sc_hd__nor2_2
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _05461_/D _09136_/A _09148_/A _06035_/A _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09125_/X sky130_fd_sc_hd__a221o_1
X_06337_ _06436_/A _06409_/B vssd1 vssd1 vccd1 vccd1 _06872_/A sky130_fd_sc_hd__and2_1
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09056_ _07713_/A _08965_/Y _09036_/X _09052_/X _09055_/X vssd1 vssd1 vccd1 vccd1
+ _09056_/X sky130_fd_sc_hd__a221o_1
X_06268_ _06558_/B _06360_/A _06267_/Y vssd1 vssd1 vccd1 vccd1 _06275_/A sky130_fd_sc_hd__o21ai_1
X_08007_ input26/X _08002_/X _08005_/X _08006_/X vssd1 vssd1 vccd1 vccd1 _10667_/D
+ sky130_fd_sc_hd__o211a_1
X_06199_ _10441_/A vssd1 vssd1 vccd1 vccd1 _07977_/A sky130_fd_sc_hd__buf_2
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07395__A1 _07393_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09958_ _09958_/A _09959_/A vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__or2b_1
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08909_ _08658_/X _08907_/Y _08908_/X vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__a21oi_1
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09889_ _09890_/B _09889_/B vssd1 vssd1 vccd1 vccd1 _09961_/B sky130_fd_sc_hd__and2b_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10802_ _10808_/CLK _10802_/D vssd1 vssd1 vccd1 vccd1 _10802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10733_ _10768_/CLK _10733_/D vssd1 vssd1 vccd1 vccd1 _10733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07855__C1 _07854_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__B _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10664_ _10811_/CLK _10664_/D vssd1 vssd1 vccd1 vccd1 _10664_/Q sky130_fd_sc_hd__dfxtp_1
X_10595_ _10878_/CLK _10595_/D vssd1 vssd1 vccd1 vccd1 _10595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput60 _10847_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[13] sky130_fd_sc_hd__buf_2
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput71 _10857_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[23] sky130_fd_sc_hd__buf_2
XFILLER_96_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput82 _10838_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_122_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10029_ _10029_/A _10029_/B vssd1 vssd1 vccd1 vccd1 _10105_/B sky130_fd_sc_hd__xor2_2
XFILLER_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05570_ _08339_/A vssd1 vssd1 vccd1 vccd1 _05570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ _07235_/C _07235_/B _07515_/A _07239_/Y vssd1 vssd1 vccd1 vccd1 _07246_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07171_ _07196_/A _07184_/B _07170_/X vssd1 vssd1 vccd1 vccd1 _07192_/A sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_41_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06122_ _06122_/A vssd1 vssd1 vccd1 vccd1 _10583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06053_ _10701_/Q _08268_/A vssd1 vssd1 vccd1 vccd1 _06053_/X sky130_fd_sc_hd__xor2_1
XFILLER_98_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _09812_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__xnor2_2
XFILLER_100_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09743_ _09743_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__xor2_1
X_06955_ _07671_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07662_/B sky130_fd_sc_hd__nor2_1
X_05906_ _05906_/A _05906_/B vssd1 vssd1 vccd1 vccd1 _05906_/X sky130_fd_sc_hd__and2_1
XFILLER_67_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09674_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__nand2_1
X_06886_ _06886_/A _06886_/B vssd1 vssd1 vccd1 vccd1 _06891_/A sky130_fd_sc_hd__xor2_4
X_05837_ _08327_/A vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__buf_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08625_ _08600_/X _08628_/C _10791_/Q vssd1 vssd1 vccd1 vccd1 _08626_/C sky130_fd_sc_hd__a21o_1
XFILLER_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08556_ _10771_/Q _08547_/B _10772_/Q vssd1 vssd1 vccd1 vccd1 _08557_/C sky130_fd_sc_hd__a21o_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05768_ _05766_/Y _10569_/Q _10568_/Q _05767_/Y vssd1 vssd1 vccd1 vccd1 _05768_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09250__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _07534_/C _07507_/B vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__nor2_2
X_05699_ _05896_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__inv_2
XANTENNA__07837__C1 _07836_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _08935_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__and2_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07438_ _07570_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _07726_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09054__A1 _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07369_ _07369_/A _07369_/B _07462_/A vssd1 vssd1 vccd1 vccd1 _07370_/B sky130_fd_sc_hd__nor3_1
X_09108_ _08974_/A _09106_/X _09107_/Y _09079_/A _10719_/Q vssd1 vssd1 vccd1 vccd1
+ _09108_/X sky130_fd_sc_hd__a32o_1
XFILLER_108_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ _10526_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10380_/X sky130_fd_sc_hd__a21bo_1
XFILLER_124_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09039_ _05455_/X _09020_/B _06129_/B _05733_/X _09263_/A vssd1 vssd1 vccd1 vccd1
+ _09039_/X sky130_fd_sc_hd__o221a_1
XANTENNA__06114__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05953__A _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08868__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _10737_/CLK _10716_/D vssd1 vssd1 vccd1 vccd1 _10716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10647_ _10673_/CLK _10647_/D vssd1 vssd1 vccd1 vccd1 _10647_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ _10935_/CLK _10578_/D vssd1 vssd1 vccd1 vccd1 _10578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06024__A _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10363__B1 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06740_ _06775_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _06741_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06671_ _06671_/A _06671_/B vssd1 vssd1 vccd1 vccd1 _06684_/A sky130_fd_sc_hd__nor2_1
X_05622_ _10551_/Q _05626_/A vssd1 vssd1 vccd1 vccd1 _05623_/B sky130_fd_sc_hd__nand2_1
X_08410_ _08547_/A _10761_/Q vssd1 vssd1 vccd1 vccd1 _08410_/X sky130_fd_sc_hd__or2_1
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09390_ _09390_/A _09390_/B vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__xnor2_1
XFILLER_17_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08341_ _08332_/A _08332_/B _05570_/X vssd1 vssd1 vccd1 vccd1 _08341_/Y sky130_fd_sc_hd__o21ai_1
X_05553_ _10553_/Q _10552_/Q _05623_/A vssd1 vssd1 vccd1 vccd1 _05663_/B sky130_fd_sc_hd__or3_2
XANTENNA__07819__C1 hold20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08272_ _08270_/X _08272_/B vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__and2b_1
X_05484_ _05482_/X _05470_/B _05495_/A _09020_/A _05483_/Y vssd1 vssd1 vccd1 vccd1
+ _10543_/D sky130_fd_sc_hd__a221o_1
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07223_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07223_/X sky130_fd_sc_hd__and2_1
XFILLER_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07154_ _07296_/A _07309_/A _07309_/B _07153_/Y vssd1 vssd1 vccd1 vccd1 _07285_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08414__A _08414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06105_ _10700_/Q _06105_/B vssd1 vssd1 vccd1 vccd1 _08267_/B sky130_fd_sc_hd__or2_1
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08795__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07085_ _07326_/A _07188_/B _07178_/A _07086_/B vssd1 vssd1 vccd1 vccd1 _07087_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_133_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06036_ _08115_/A _08119_/A _05405_/A _08059_/A _06035_/X vssd1 vssd1 vccd1 vccd1
+ _06036_/X sky130_fd_sc_hd__a221o_1
XFILLER_105_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10354__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07987_ _08015_/A vssd1 vssd1 vccd1 vccd1 _07987_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input1_A io_ba_match vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09726_ _09787_/B _09726_/B vssd1 vssd1 vccd1 vccd1 _09727_/B sky130_fd_sc_hd__xnor2_2
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06938_ _06938_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _07625_/A sky130_fd_sc_hd__xnor2_4
XFILLER_27_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06869_ _06869_/A _06869_/B vssd1 vssd1 vccd1 vccd1 _07761_/B sky130_fd_sc_hd__xnor2_2
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09657_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09713_/A sky130_fd_sc_hd__xor2_1
X_08608_ _08611_/B _08649_/A _08608_/C vssd1 vssd1 vccd1 vccd1 _08609_/A sky130_fd_sc_hd__and3b_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__and2_1
XFILLER_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08539_ _08547_/A _10767_/Q _10768_/Q vssd1 vssd1 vccd1 vccd1 _08540_/C sky130_fd_sc_hd__a21o_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10501_ _10515_/B vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_7_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08324__A _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _10432_/A _10432_/B _10432_/C vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__and3_1
XFILLER_109_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10363_ _08491_/X _07635_/A _09408_/X _10930_/Q vssd1 vssd1 vccd1 vccd1 _10930_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10294_ _07008_/A _10283_/X _10292_/X _10293_/X vssd1 vssd1 vccd1 vccd1 _10908_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06013__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10345__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_9_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06019__A _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06252__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08529__B1 _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07910_/X sky130_fd_sc_hd__clkbuf_1
X_08890_ _10824_/Q _08876_/A _08928_/B vssd1 vssd1 vccd1 vccd1 _08890_/X sky130_fd_sc_hd__o21a_1
XFILLER_68_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07841_ _10874_/Q _07845_/B vssd1 vssd1 vccd1 vccd1 _07841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07772_ _10513_/A _07776_/B _06848_/B _06847_/A vssd1 vssd1 vccd1 vccd1 _07778_/A
+ sky130_fd_sc_hd__a31o_1
X_09511_ _09599_/B vssd1 vssd1 vccd1 vccd1 _09761_/C sky130_fd_sc_hd__clkbuf_2
X_06723_ _06638_/A _06638_/B _06721_/Y _06714_/B _06722_/Y vssd1 vssd1 vccd1 vccd1
+ _06725_/B sky130_fd_sc_hd__o32a_1
XFILLER_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06654_ _06654_/A _06654_/B vssd1 vssd1 vccd1 vccd1 _06700_/B sky130_fd_sc_hd__nor2_1
X_09442_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__nand2_1
X_05605_ _10698_/Q _05605_/B vssd1 vssd1 vccd1 vccd1 _05605_/X sky130_fd_sc_hd__or2_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09373_ _09343_/A _09346_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09373_/Y sky130_fd_sc_hd__o21bai_1
X_06585_ _06585_/A _06585_/B vssd1 vssd1 vccd1 vccd1 _06591_/B sky130_fd_sc_hd__xnor2_1
X_08324_ _08324_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08324_/Y sky130_fd_sc_hd__nand2_1
X_05536_ _05818_/B _05536_/B vssd1 vssd1 vccd1 vccd1 _05652_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08255_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08342_/B sky130_fd_sc_hd__clkbuf_2
X_05467_ _05467_/A _05467_/B _05467_/C _05467_/D vssd1 vssd1 vccd1 vccd1 _05467_/X
+ sky130_fd_sc_hd__or4_4
XANTENNA__09009__B2 _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08186_ _08186_/A vssd1 vssd1 vccd1 vccd1 _10692_/D sky130_fd_sc_hd__clkbuf_1
X_05398_ _05398_/A _05398_/B vssd1 vssd1 vccd1 vccd1 _05487_/A sky130_fd_sc_hd__xnor2_1
X_07206_ _07301_/A _07302_/A _07205_/A vssd1 vssd1 vccd1 vccd1 _07208_/B sky130_fd_sc_hd__o21a_1
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07137_ _07137_/A _07327_/A _07137_/C vssd1 vssd1 vccd1 vccd1 _07139_/B sky130_fd_sc_hd__and3_1
XANTENNA__07983__A _07983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06243__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07068_ _10983_/Q _07197_/B vssd1 vssd1 vccd1 vccd1 _07312_/A sky130_fd_sc_hd__nand2_2
X_06019_ _06019_/A _08212_/A vssd1 vssd1 vccd1 vccd1 _08258_/A sky130_fd_sc_hd__and2_1
XFILLER_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09709_ _09710_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__nor2_1
X_10981_ _10981_/CLK _10981_/D vssd1 vssd1 vccd1 vccd1 _10981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08054__A _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10415_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10415_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07982__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _10355_/A vssd1 vssd1 vccd1 vccd1 _10346_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ _10265_/A _10287_/B _10265_/B vssd1 vssd1 vccd1 vccd1 _10277_/X sky130_fd_sc_hd__o21ba_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06370_ _06409_/B vssd1 vssd1 vccd1 vccd1 _06408_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05321_ _10676_/Q vssd1 vssd1 vccd1 vccd1 _05830_/A sky130_fd_sc_hd__buf_2
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10254__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08040_ _06115_/A _06115_/B _10580_/Q vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__o21a_2
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09991_ _10068_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__nand2_1
XFILLER_115_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08942_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__or2_1
XFILLER_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06212__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _08873_/A _08873_/B vssd1 vssd1 vccd1 vccd1 _08873_/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07725__A1 _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07824_ hold18/X _07824_/B vssd1 vssd1 vccd1 vccd1 _07824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07755_ _07755_/A _07755_/B vssd1 vssd1 vccd1 vccd1 _07756_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06706_ _06719_/A _06627_/B _06719_/C _06841_/A vssd1 vssd1 vccd1 vccd1 _06706_/X
+ sky130_fd_sc_hd__a22o_1
X_07686_ _09409_/A _09409_/B _07666_/A vssd1 vssd1 vccd1 vccd1 _07689_/A sky130_fd_sc_hd__o21a_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09425_ _09424_/A _09418_/A _09677_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__a21o_1
X_06637_ _06638_/A _06638_/B vssd1 vssd1 vccd1 vccd1 _06715_/A sky130_fd_sc_hd__or2_1
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _09356_/A _10888_/Q vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__xnor2_4
X_06568_ _06568_/A _06568_/B _06581_/A vssd1 vssd1 vccd1 vccd1 _06570_/B sky130_fd_sc_hd__and3_1
X_08307_ _05844_/A _08058_/X _08306_/Y _06011_/X vssd1 vssd1 vccd1 vccd1 _08307_/X
+ sky130_fd_sc_hd__o211a_1
X_09287_ _08342_/A _09286_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__mux2_1
X_05519_ _07911_/A _05471_/X _05474_/Y _05442_/Y vssd1 vssd1 vccd1 vccd1 _10567_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06499_ _06561_/B vssd1 vssd1 vccd1 vccd1 _06517_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08238_ _08114_/X _08251_/C _08233_/Y _08237_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08238_/X sky130_fd_sc_hd__o311a_1
XFILLER_119_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08169_ _08169_/A _08169_/B _08169_/C vssd1 vssd1 vccd1 vccd1 _08180_/B sky130_fd_sc_hd__and3_1
XFILLER_119_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ _10197_/Y _10198_/Y _10199_/Y vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _10131_/A _10131_/B _10131_/C vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__and3_1
XANTENNA__08321__B _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10062_ _10062_/A _09338_/X vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__or2b_1
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07716__A1 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05961__A input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08141__A1 _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08049__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10964_ _10968_/CLK _10964_/D vssd1 vssd1 vccd1 vccd1 _10964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10895_ _10909_/CLK _10895_/D vssd1 vssd1 vccd1 vccd1 _10895_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07888__A _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10329_ _10334_/B _10327_/A _10329_/S vssd1 vssd1 vccd1 vccd1 _10330_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09327__B _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06032__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05870_ _05358_/A _05823_/A _05869_/Y vssd1 vssd1 vccd1 vccd1 _05870_/X sky130_fd_sc_hd__o21a_1
XFILLER_94_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07540_ _07540_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07540_/X sky130_fd_sc_hd__or2b_1
XFILLER_35_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07471_ _07471_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _09274_/A vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06422_ _06506_/B vssd1 vssd1 vccd1 vccd1 _06540_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09141_ _09153_/A _09141_/B vssd1 vssd1 vccd1 vccd1 _10843_/D sky130_fd_sc_hd__nor2_4
X_06353_ _06550_/B vssd1 vssd1 vccd1 vccd1 _06554_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05304_ _10666_/Q _05358_/A vssd1 vssd1 vccd1 vccd1 _05353_/A sky130_fd_sc_hd__or2_1
X_09072_ _10936_/Q _10394_/C _10430_/B _10952_/Q vssd1 vssd1 vccd1 vccd1 _09072_/X
+ sky130_fd_sc_hd__a22o_1
X_08023_ _08023_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08023_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06207__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06284_ _10918_/Q _07113_/A vssd1 vssd1 vccd1 vccd1 _06284_/X sky130_fd_sc_hd__and2_1
XFILLER_135_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09974_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__and2_1
XFILLER_131_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08925_ _08658_/X _08923_/Y _08924_/X vssd1 vssd1 vccd1 vccd1 _08926_/B sky130_fd_sc_hd__a21oi_1
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08856_ _10821_/Q _08856_/B vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_36_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07807_ _07850_/A vssd1 vssd1 vccd1 vccd1 _07807_/X sky130_fd_sc_hd__buf_4
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05999_ input41/X vssd1 vssd1 vccd1 vccd1 _10528_/A sky130_fd_sc_hd__clkbuf_4
X_08787_ _06195_/X _08785_/X _08786_/X _10812_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08787_/X sky130_fd_sc_hd__o221a_1
X_07738_ _07738_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07739_/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07669_ _07669_/A vssd1 vssd1 vccd1 vccd1 _07673_/A sky130_fd_sc_hd__inv_2
X_10680_ _10839_/CLK _10680_/D vssd1 vssd1 vccd1 vccd1 _10680_/Q sky130_fd_sc_hd__dfxtp_1
X_09408_ _10115_/A vssd1 vssd1 vccd1 vccd1 _09408_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _10911_/Q _10895_/Q vssd1 vssd1 vccd1 vccd1 _10065_/C sky130_fd_sc_hd__or2b_1
XFILLER_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05956__A _05956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08332__A _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07937__A1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10114_ _10112_/Y _10113_/X _10880_/Q _09406_/X vssd1 vssd1 vccd1 vccd1 _10880_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08986__B _08989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06787__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _10045_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08362__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08362__B2 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09311__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10947_ _10978_/CLK _10947_/D vssd1 vssd1 vccd1 vccd1 _10947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10878_ _10878_/CLK _10878_/D vssd1 vssd1 vccd1 vccd1 _10878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06027__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09338__A _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07928__B2 _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08050__B1 _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _07655_/A vssd1 vssd1 vccd1 vccd1 _07715_/D sky130_fd_sc_hd__clkbuf_2
X_05922_ _08130_/A _05900_/X _05897_/X _05896_/A _05921_/X vssd1 vssd1 vccd1 vccd1
+ _05922_/X sky130_fd_sc_hd__o221a_1
X_08710_ _08725_/B _08710_/B vssd1 vssd1 vccd1 vccd1 _08710_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_79_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09690_ _09690_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09754_/A sky130_fd_sc_hd__xnor2_2
X_05853_ _05340_/A _05854_/B _05852_/Y vssd1 vssd1 vccd1 vccd1 _05853_/X sky130_fd_sc_hd__o21a_1
X_08641_ _08641_/A vssd1 vssd1 vccd1 vccd1 _10795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05784_ _05803_/A _05769_/Y _05780_/Y _08304_/A _05783_/X vssd1 vssd1 vccd1 vccd1
+ _05785_/C sky130_fd_sc_hd__o221a_1
X_08572_ _10777_/Q _08572_/B _10775_/Q vssd1 vssd1 vccd1 vccd1 _08578_/D sky130_fd_sc_hd__and3_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _07525_/B _07523_/B vssd1 vssd1 vccd1 vccd1 _07649_/A sky130_fd_sc_hd__nand2_1
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07454_ _07454_/A _07454_/B _07454_/C vssd1 vssd1 vccd1 vccd1 _07455_/B sky130_fd_sc_hd__or3_1
X_06405_ _06513_/D vssd1 vssd1 vccd1 vccd1 _06428_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07385_ _07378_/Y _07458_/B _09304_/A _07384_/X vssd1 vssd1 vccd1 vccd1 _07386_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09124_ _09124_/A _09124_/B _09124_/C vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__nor3_4
X_06336_ _06522_/B vssd1 vssd1 vccd1 vccd1 _06409_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09055_ _05912_/B _08972_/X _08974_/A _09054_/X vssd1 vssd1 vccd1 vccd1 _09055_/X
+ sky130_fd_sc_hd__o211a_1
X_06267_ _10916_/Q _10899_/Q vssd1 vssd1 vccd1 vccd1 _06267_/Y sky130_fd_sc_hd__nand2_1
X_08006_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08006_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06198_ _09403_/A vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07395__A2 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09957_ _09887_/A _09887_/B _09956_/X vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__a21o_1
XFILLER_106_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08908_ input36/X _08830_/X _08831_/X _10827_/Q vssd1 vssd1 vccd1 vccd1 _08908_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_100_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09888_ _09626_/A _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09889_/B sky130_fd_sc_hd__a21boi_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08835_/Y _08836_/X _08838_/X vssd1 vssd1 vccd1 vccd1 _10818_/D sky130_fd_sc_hd__o21a_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10801_ _10945_/CLK _10801_/D vssd1 vssd1 vccd1 vccd1 _10801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10732_ _10768_/CLK _10732_/D vssd1 vssd1 vccd1 vccd1 _10732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10663_ _10811_/CLK _10663_/D vssd1 vssd1 vccd1 vccd1 _10663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10594_ _10958_/CLK _10594_/D vssd1 vssd1 vccd1 vccd1 _10594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput61 _10848_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput83 _10839_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput72 _10858_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10028_ _10100_/B _10028_/B vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07170_ _07222_/A _07164_/B _07169_/B _07248_/A vssd1 vssd1 vccd1 vccd1 _07170_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08271__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06121_ _08483_/A _06121_/B vssd1 vssd1 vccd1 vccd1 _06122_/A sky130_fd_sc_hd__and2_1
XFILLER_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06052_ _06052_/A vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__buf_2
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09133__A1_N _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09811_ _10493_/A _09811_/B _09811_/C vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__and3_1
XFILLER_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09742_ _09870_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09743_/B sky130_fd_sc_hd__or2_1
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06954_ _07675_/B _07676_/B vssd1 vssd1 vccd1 vccd1 _07670_/B sky130_fd_sc_hd__nand2_1
X_05905_ _05905_/A _05905_/B vssd1 vssd1 vccd1 vccd1 _05906_/B sky130_fd_sc_hd__nand2_1
X_09673_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__or2_1
X_06885_ _06885_/A _06885_/B vssd1 vssd1 vccd1 vccd1 _06886_/B sky130_fd_sc_hd__xnor2_4
X_05836_ _05836_/A _05836_/B vssd1 vssd1 vccd1 vccd1 _05836_/X sky130_fd_sc_hd__and2_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _10791_/Q _08624_/B _08628_/C vssd1 vssd1 vccd1 vccd1 _08631_/C sky130_fd_sc_hd__and3_1
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05767_ _10707_/Q vssd1 vssd1 vccd1 vccd1 _05767_/Y sky130_fd_sc_hd__clkinv_2
X_08555_ _08531_/X _08559_/B _10772_/Q _08531_/A vssd1 vssd1 vccd1 vccd1 _08557_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07506_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07507_/B sky130_fd_sc_hd__and2_1
XFILLER_35_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08147__A _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05698_ _08181_/A _10553_/Q _10552_/Q _08173_/A vssd1 vssd1 vccd1 vccd1 _05717_/B
+ sky130_fd_sc_hd__a22o_1
X_08486_ _10782_/Q _10745_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08487_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09039__C1 _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07437_ _06993_/A _07570_/C _07678_/A vssd1 vssd1 vccd1 vccd1 _07438_/B sky130_fd_sc_hd__o21ai_1
XFILLER_22_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_53_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10878_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07368_ _07369_/B _07462_/A _07369_/A vssd1 vssd1 vccd1 vccd1 _07412_/C sky130_fd_sc_hd__o21a_1
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09107_ _09107_/A _09107_/B vssd1 vssd1 vccd1 vccd1 _09107_/Y sky130_fd_sc_hd__nand2_1
X_06319_ _10924_/Q _10907_/Q vssd1 vssd1 vccd1 vccd1 _06321_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07299_ _07298_/A _07298_/B _07298_/C vssd1 vssd1 vccd1 vccd1 _07300_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09038_ _10715_/Q _08999_/X _09037_/Y _10802_/Q vssd1 vssd1 vccd1 vccd1 _09038_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_132_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_68_clock _10985_/CLK vssd1 vssd1 vccd1 vccd1 _10982_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06040__A2 _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10372__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06067__A2_N _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10737_/CLK _10715_/D vssd1 vssd1 vccd1 vccd1 _10715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ _10646_/CLK _10646_/D vssd1 vssd1 vccd1 vccd1 _10646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10577_ _10652_/CLK _10577_/D vssd1 vssd1 vccd1 vccd1 _10577_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06670_ _06670_/A _06670_/B vssd1 vssd1 vccd1 vccd1 _06671_/B sky130_fd_sc_hd__and2_1
XFILLER_36_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05621_ _10690_/Q vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__05542__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08340_ _05574_/X _08339_/C _05570_/X vssd1 vssd1 vccd1 vccd1 _08340_/Y sky130_fd_sc_hd__a21oi_1
X_05552_ _10551_/Q _05626_/A vssd1 vssd1 vccd1 vccd1 _05623_/A sky130_fd_sc_hd__or2_1
X_08271_ input29/X _08212_/X _08052_/A _08267_/A _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08272_/B sky130_fd_sc_hd__o221a_1
X_05483_ _05483_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05483_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07222_ _07222_/A _07222_/B _07250_/A vssd1 vssd1 vccd1 vccd1 _07233_/B sky130_fd_sc_hd__and3_1
XFILLER_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07153_ _07295_/B _07317_/A _07295_/A vssd1 vssd1 vccd1 vccd1 _07153_/Y sky130_fd_sc_hd__o21ai_1
X_06104_ _10699_/Q _08243_/B vssd1 vssd1 vccd1 vccd1 _06105_/B sky130_fd_sc_hd__or2_1
XFILLER_133_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07084_ _07169_/B vssd1 vssd1 vccd1 vccd1 _07178_/A sky130_fd_sc_hd__clkbuf_2
X_06035_ _06035_/A _07974_/A vssd1 vssd1 vccd1 vccd1 _06035_/X sky130_fd_sc_hd__xor2_1
XFILLER_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07986_ _06191_/X _07965_/X _07985_/Y _07977_/X vssd1 vssd1 vccd1 vccd1 _10660_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09725_ _09779_/A _09779_/B _09661_/X vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06937_ _06937_/A _06937_/B vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__xnor2_4
XFILLER_83_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ _09656_/A _09656_/B vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09261__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08607_ _08498_/X _08550_/X _08597_/B _10786_/Q vssd1 vssd1 vccd1 vccd1 _08608_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06868_ _06868_/A _06868_/B vssd1 vssd1 vccd1 vccd1 _06869_/B sky130_fd_sc_hd__nor2_1
X_05819_ _05907_/A _05909_/A _05908_/B vssd1 vssd1 vccd1 vccd1 _05905_/B sky130_fd_sc_hd__a21o_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _10508_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07774_/A sky130_fd_sc_hd__nand2_1
X_09587_ _09587_/A _09587_/B vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__nand2_1
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08538_ _08567_/D vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ _08469_/A vssd1 vssd1 vccd1 vccd1 _10739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ _10517_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__nor2_2
XFILLER_10_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06125__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ _08491_/X _06855_/A _09408_/X _10929_/Q vssd1 vssd1 vccd1 vccd1 _10929_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10293_ _10351_/A vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05964__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10345__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08226__B1 _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10629_ _10811_/CLK _10629_/D vssd1 vssd1 vccd1 vccd1 _10629_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06035__A _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06252__A2 _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10336__A1 _10291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07840_ _07827_/X _05462_/A _07823_/X _07839_/Y vssd1 vssd1 vccd1 vccd1 _10623_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07771_ _07771_/A _07771_/B vssd1 vssd1 vccd1 vccd1 _07792_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06722_ _06722_/A vssd1 vssd1 vccd1 vccd1 _06722_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09510_ _09555_/B vssd1 vssd1 vccd1 vccd1 _09692_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06653_ _06650_/A _06650_/C _06650_/B vssd1 vssd1 vccd1 vccd1 _06654_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _09441_/A _07689_/A vssd1 vssd1 vccd1 vccd1 _09442_/B sky130_fd_sc_hd__or2b_1
X_05604_ _05604_/A _05604_/B vssd1 vssd1 vccd1 vccd1 _05605_/B sky130_fd_sc_hd__and2_1
X_09372_ _09372_/A _09372_/B _09372_/C vssd1 vssd1 vccd1 vccd1 _09372_/X sky130_fd_sc_hd__or3_1
XFILLER_40_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06584_ _06584_/A _06584_/B vssd1 vssd1 vccd1 vccd1 _06591_/A sky130_fd_sc_hd__or2_1
XFILLER_24_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08323_ _08881_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _10706_/D sky130_fd_sc_hd__nor2_1
X_05535_ _10544_/Q vssd1 vssd1 vccd1 vccd1 _05536_/B sky130_fd_sc_hd__inv_2
XANTENNA__10272__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08254_ _08242_/A _08243_/B _05598_/X vssd1 vssd1 vccd1 vccd1 _08254_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_119_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05466_ _07900_/A _07896_/A _07893_/A _07889_/A vssd1 vssd1 vccd1 vccd1 _05467_/D
+ sky130_fd_sc_hd__or4_1
XANTENNA__08425__A _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08185_ _08185_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__and2_1
XANTENNA__06084__A1_N _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05397_ _05397_/A _05397_/B vssd1 vssd1 vccd1 vccd1 _05398_/B sky130_fd_sc_hd__nor2_1
X_07205_ _07205_/A _07205_/B vssd1 vssd1 vccd1 vccd1 _07302_/A sky130_fd_sc_hd__nand2_1
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08768__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07136_ _07136_/A _07136_/B vssd1 vssd1 vccd1 vccd1 _07138_/A sky130_fd_sc_hd__xnor2_1
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07067_ _07167_/B vssd1 vssd1 vccd1 vccd1 _07186_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06018_ _06023_/B vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10840__D _10840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07969_ _07969_/A vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ _09708_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09710_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10980_ _10980_/CLK _10980_/D vssd1 vssd1 vccd1 vccd1 _10980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09639_ _09588_/A _09639_/B _09696_/A vssd1 vssd1 vccd1 vccd1 _09640_/B sky130_fd_sc_hd__and3b_1
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ _10942_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10414_/X sky130_fd_sc_hd__and2_1
XFILLER_124_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08989__B _08989_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10345_ _09312_/X _07682_/B _10184_/X _10915_/Q vssd1 vssd1 vccd1 vccd1 _10915_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05993__A1 _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ _10287_/C _10287_/D vssd1 vssd1 vccd1 vccd1 _10276_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08931__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05320_ _10645_/Q vssd1 vssd1 vccd1 vccd1 _07922_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08998__A1 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05869__A _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09990_ _09990_/A _09990_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__xnor2_2
XFILLER_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05984__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08941_ _09098_/B vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__buf_2
XFILLER_130_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08872_ _10822_/Q _10821_/Q _10820_/Q _08847_/X _08840_/B vssd1 vssd1 vccd1 vccd1
+ _08873_/B sky130_fd_sc_hd__o41a_1
XFILLER_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07823_ _08557_/A vssd1 vssd1 vccd1 vccd1 _07823_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07754_ _07754_/A _07754_/B vssd1 vssd1 vccd1 vccd1 _07755_/B sky130_fd_sc_hd__xnor2_1
X_07685_ _09329_/A _09329_/B _07674_/A vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__o21a_1
X_06705_ _06719_/A _06719_/C vssd1 vssd1 vccd1 vccd1 _07791_/A sky130_fd_sc_hd__nand2_2
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09424_ _09424_/A _09811_/B _09677_/B vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__nand3_1
X_06636_ _06431_/A _06431_/B _06434_/A vssd1 vssd1 vccd1 vccd1 _06638_/B sky130_fd_sc_hd__o21a_1
XFILLER_25_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06161__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09355_ _10905_/Q _10889_/Q vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__or2b_1
XFILLER_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06567_ _06567_/A _06567_/B vssd1 vssd1 vccd1 vccd1 _06581_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08306_ _08317_/B _08306_/B _08306_/C vssd1 vssd1 vccd1 vccd1 _08306_/Y sky130_fd_sc_hd__nand3_1
X_09286_ _08339_/A _07922_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09286_/X sky130_fd_sc_hd__mux2_1
X_05518_ _05332_/Y _05517_/X _05513_/X _07907_/A vssd1 vssd1 vccd1 vccd1 _10566_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06498_ _10972_/Q vssd1 vssd1 vccd1 vccd1 _06561_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10835__D _10835_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08237_ _08243_/B _08061_/A _08234_/X _08235_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08237_/X sky130_fd_sc_hd__a311o_1
X_05449_ _10647_/Q _05525_/B _05448_/X vssd1 vssd1 vccd1 vccd1 _05490_/A sky130_fd_sc_hd__o21ai_4
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_32_clock_A _10704_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08168_ _08157_/X _08161_/X _08163_/Y _08167_/X vssd1 vssd1 vccd1 vccd1 _10690_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_106_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08099_ _08038_/X _08074_/X _08098_/Y _08044_/X _05905_/A vssd1 vssd1 vccd1 vccd1
+ _08099_/X sky130_fd_sc_hd__a32o_1
XFILLER_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07119_ _10983_/Q _07142_/B vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__and2_1
XFILLER_134_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10130_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08677__B1 _08676_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _10968_/CLK _10963_/D vssd1 vssd1 vccd1 vccd1 _10963_/Q sky130_fd_sc_hd__dfxtp_1
X_10894_ _10909_/CLK _10894_/D vssd1 vssd1 vccd1 vccd1 _10894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10328_ _10312_/A _10310_/X _10320_/A _10327_/Y vssd1 vssd1 vccd1 vccd1 _10334_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10259_ _10243_/A _10250_/X _10245_/B vssd1 vssd1 vccd1 vccd1 _10259_/X sky130_fd_sc_hd__a21o_1
XFILLER_94_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07470_ _07470_/A _07470_/B _07482_/A vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__nor3_1
X_06421_ _06421_/A _06732_/B vssd1 vssd1 vccd1 vccd1 _06506_/B sky130_fd_sc_hd__xnor2_2
X_09140_ _09112_/X _09135_/Y _09139_/X vssd1 vssd1 vccd1 vccd1 _09141_/B sky130_fd_sc_hd__a21oi_1
X_06352_ _06352_/A _06352_/B _06352_/C vssd1 vssd1 vccd1 vccd1 _06550_/B sky130_fd_sc_hd__or3_1
X_05303_ _10665_/Q _10664_/Q _05363_/A vssd1 vssd1 vccd1 vccd1 _05358_/A sky130_fd_sc_hd__or3_2
X_09071_ _09904_/A vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_30_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06283_ _10901_/Q vssd1 vssd1 vccd1 vccd1 _07113_/A sky130_fd_sc_hd__buf_2
X_08022_ input33/X _08015_/X _08021_/Y _08019_/X vssd1 vssd1 vccd1 vccd1 _10673_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08199__A2 _08061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09973_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08924_ input39/X _08830_/X _08831_/X _10829_/Q vssd1 vssd1 vccd1 vccd1 _08924_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08855_ _10821_/Q _08865_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08786_ _08820_/A vssd1 vssd1 vccd1 vccd1 _08786_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07806_ _10160_/A _07804_/Y _07805_/X _10881_/Q vssd1 vssd1 vccd1 vccd1 _07850_/A
+ sky130_fd_sc_hd__a211o_2
X_05998_ _09090_/A vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07737_ _07581_/A _07581_/B _07580_/A vssd1 vssd1 vccd1 vccd1 _07738_/B sky130_fd_sc_hd__o21a_1
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07668_ _07668_/A _07668_/B vssd1 vssd1 vccd1 vccd1 _07669_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09407_ _09402_/X _09405_/X _10868_/Q _09406_/X vssd1 vssd1 vccd1 vccd1 _10868_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06619_ _06668_/A _06668_/B _06618_/X vssd1 vssd1 vccd1 vccd1 _06692_/A sky130_fd_sc_hd__a21o_1
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07599_/X sky130_fd_sc_hd__or2_1
X_09338_ _10912_/Q _10896_/Q vssd1 vssd1 vccd1 vccd1 _09338_/X sky130_fd_sc_hd__or2b_1
XFILLER_21_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09269_ _08318_/A _09268_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09269_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07229__A _07229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09139__B2 _10721_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _10112_/A _10112_/B _09480_/X vssd1 vssd1 vccd1 vccd1 _10113_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input32_A io_wbs_m2s_data[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10044_ hold14/A _09572_/X _10042_/Y _10043_/X vssd1 vssd1 vccd1 vccd1 _10879_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09311__A1 _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07899__A _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946_ _10946_/CLK _10946_/D vssd1 vssd1 vccd1 vccd1 _10946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10877_ _10878_/CLK _10877_/D vssd1 vssd1 vccd1 vccd1 _10877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06027__B _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08523__A _08935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08050__A1 _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ _07678_/A vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05921_ _05726_/A _05902_/Y _05900_/X _10687_/Q _05920_/X vssd1 vssd1 vccd1 vccd1
+ _05921_/X sky130_fd_sc_hd__a221o_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05852_ _08289_/A _05852_/B vssd1 vssd1 vccd1 vccd1 _05852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08640_ _08638_/X _08640_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _08641_/A sky130_fd_sc_hd__and3b_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05783_ _05781_/Y _10566_/Q _10565_/Q _05782_/Y vssd1 vssd1 vccd1 vccd1 _05783_/X
+ sky130_fd_sc_hd__o22a_1
X_08571_ _08572_/B _08565_/X _10777_/Q vssd1 vssd1 vccd1 vccd1 _08574_/B sky130_fd_sc_hd__a21o_1
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07522_ _07522_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07523_/B sky130_fd_sc_hd__or2_1
XFILLER_62_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07453_ _07454_/B _07454_/C _07454_/A vssd1 vssd1 vccd1 vccd1 _07455_/A sky130_fd_sc_hd__o21ai_1
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06404_ _06461_/B vssd1 vssd1 vccd1 vccd1 _06426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09123_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09123_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07384_ _07384_/A _07384_/B vssd1 vssd1 vccd1 vccd1 _07384_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08813__B1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06335_ _06515_/B vssd1 vssd1 vccd1 vccd1 _06522_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _05905_/A _08995_/X _09053_/X _08981_/A vssd1 vssd1 vccd1 vccd1 _09054_/X
+ sky130_fd_sc_hd__a211o_1
X_06266_ _10916_/Q _10899_/Q vssd1 vssd1 vccd1 vccd1 _06360_/A sky130_fd_sc_hd__xnor2_2
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08005_ _08244_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08005_/X sky130_fd_sc_hd__or2_1
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06197_ _06197_/A _06204_/B vssd1 vssd1 vccd1 vccd1 _06197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07991__B _08021_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _09886_/B _09956_/B vssd1 vssd1 vccd1 vccd1 _09956_/X sky130_fd_sc_hd__and2b_1
XFILLER_112_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08907_/Y sky130_fd_sc_hd__xnor2_1
X_09887_ _09887_/A _09887_/B vssd1 vssd1 vccd1 vccd1 _09890_/B sky130_fd_sc_hd__xor2_1
XFILLER_58_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08838_ input26/X _08785_/X _08786_/X _10818_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08838_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08769_ _08766_/Y _08767_/X _08768_/X vssd1 vssd1 vccd1 vccd1 _10810_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10800_ _10803_/CLK _10800_/D vssd1 vssd1 vccd1 vccd1 _10800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10731_ _10768_/CLK _10731_/D vssd1 vssd1 vccd1 vccd1 _10731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10662_ _10811_/CLK _10662_/D vssd1 vssd1 vccd1 vccd1 _10662_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06128__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _10958_/CLK _10593_/D vssd1 vssd1 vccd1 vccd1 _10593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05967__A input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06026__A_N _10581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06798__A _06845_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput62 _10849_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput73 _10859_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[25] sky130_fd_sc_hd__buf_2
Xoutput84 _10840_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_48_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10027_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__or2_1
XFILLER_49_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_clock_A _10981_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08099__B2 _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09296__A0 _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10929_ _10930_/CLK _10929_/D vssd1 vssd1 vccd1 vccd1 _10929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08271__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06120_ input16/X _06019_/A _06120_/S vssd1 vssd1 vccd1 vccd1 _06121_/B sky130_fd_sc_hd__mux2_1
X_06051_ _08130_/A vssd1 vssd1 vccd1 vccd1 _09104_/A sky130_fd_sc_hd__clkinv_2
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09810_ _09810_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09811_/C sky130_fd_sc_hd__nand2_1
XFILLER_87_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09741_ _10480_/A _10129_/B _10122_/B _10478_/A vssd1 vssd1 vccd1 vccd1 _09742_/B
+ sky130_fd_sc_hd__a22oi_1
X_06953_ _06769_/A _06460_/B _06558_/X vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08326__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05904_ _05904_/A _05904_/B vssd1 vssd1 vccd1 vccd1 _05904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09672_ _09670_/Y _09672_/B vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__and2b_1
X_06884_ _06884_/A _06884_/B vssd1 vssd1 vccd1 vccd1 _06886_/A sky130_fd_sc_hd__or2_2
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05835_ _08025_/A _05838_/B _08027_/A vssd1 vssd1 vccd1 vccd1 _05836_/B sky130_fd_sc_hd__o21ai_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08623_ _10790_/Q _10789_/Q _08623_/C _08623_/D vssd1 vssd1 vccd1 vccd1 _08628_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_55_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05766_ _10708_/Q vssd1 vssd1 vccd1 vccd1 _05766_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__09287__A0 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _08583_/A _08554_/B vssd1 vssd1 vccd1 vccd1 _10771_/D sky130_fd_sc_hd__nor2_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07505_ _07505_/A _07505_/B vssd1 vssd1 vccd1 vccd1 _07505_/X sky130_fd_sc_hd__and2_1
X_05697_ _05885_/A vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__clkinv_2
X_08485_ _09090_/A vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07436_ _07727_/A _07433_/A _07729_/B _07713_/A vssd1 vssd1 vccd1 vccd1 _07445_/B
+ sky130_fd_sc_hd__a22o_1
X_07367_ _07412_/B _07367_/B vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _06050_/X _08995_/A _09105_/X _09107_/B vssd1 vssd1 vccd1 vccd1 _09106_/X
+ sky130_fd_sc_hd__a211o_1
X_06318_ _06755_/A _06729_/A vssd1 vssd1 vccd1 vccd1 _06318_/X sky130_fd_sc_hd__or2_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09037_ _09037_/A _09079_/A vssd1 vssd1 vccd1 vccd1 _09037_/Y sky130_fd_sc_hd__nor2_1
X_07298_ _07298_/A _07298_/B _07298_/C vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__and3_1
XANTENNA__10843__D _10843_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06249_ _10613_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06249_/X sky130_fd_sc_hd__or2_1
XANTENNA__08014__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09939_ _09940_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__or2_1
XFILLER_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10935_/CLK _10714_/D vssd1 vssd1 vccd1 vccd1 _10714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10645_ _10676_/CLK _10645_/D vssd1 vssd1 vccd1 vccd1 _10645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09169__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09345__A_N _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10576_ _10652_/CLK _10576_/D vssd1 vssd1 vccd1 vccd1 _10576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_114_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__A2 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09632__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05620_ _10692_/Q vssd1 vssd1 vccd1 vccd1 _05885_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09269__A0 _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09351__B _10906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08248__A _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05551_ _10550_/Q _10549_/Q _05630_/A vssd1 vssd1 vccd1 vccd1 _05626_/A sky130_fd_sc_hd__or3_1
XFILLER_17_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05482_ _10574_/Q vssd1 vssd1 vccd1 vccd1 _05482_/X sky130_fd_sc_hd__clkbuf_4
X_08270_ _08263_/X _08276_/B _08266_/Y _08269_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08270_/X sky130_fd_sc_hd__o311a_1
XFILLER_60_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07221_ _07250_/A _07217_/B _07218_/X _07242_/B vssd1 vssd1 vccd1 vccd1 _07233_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_118_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07152_ _07309_/A _07152_/B _07322_/A vssd1 vssd1 vccd1 vccd1 _07317_/A sky130_fd_sc_hd__and3_1
XFILLER_20_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06103_ _10698_/Q _10697_/Q _10696_/Q _08218_/B vssd1 vssd1 vccd1 vccd1 _08243_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_106_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07083_ _07083_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07169_/B sky130_fd_sc_hd__xnor2_2
X_06034_ _10686_/Q vssd1 vssd1 vccd1 vccd1 _08115_/A sky130_fd_sc_hd__inv_2
XFILLER_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07985_ _07985_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _07985_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09724_ _09724_/A _09723_/Y vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__or2b_1
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06936_ _06936_/A _06936_/B vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__xnor2_4
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06867_ _06866_/B _06867_/B vssd1 vssd1 vccd1 vccd1 _06868_/B sky130_fd_sc_hd__and2b_1
X_09655_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09656_/B sky130_fd_sc_hd__nor2_1
X_05818_ _05818_/A _05818_/B vssd1 vssd1 vccd1 vccd1 _05908_/B sky130_fd_sc_hd__nor2_1
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08606_ _10786_/Q _10785_/Q _08617_/B vssd1 vssd1 vccd1 vccd1 _08611_/B sky130_fd_sc_hd__and3_1
XFILLER_43_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ _06845_/A vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__buf_2
X_09586_ _09639_/B _09834_/B _09642_/A _09696_/A vssd1 vssd1 vccd1 vccd1 _09587_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__07062__A _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05749_ _05749_/A _10564_/Q vssd1 vssd1 vccd1 vccd1 _05749_/X sky130_fd_sc_hd__and2_1
X_08537_ _10291_/S _08686_/A _08462_/A vssd1 vssd1 vccd1 vccd1 _08567_/D sky130_fd_sc_hd__a21oi_1
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10838__D _10838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _08477_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__or2_1
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07419_ _07416_/A _07727_/B _07713_/B _07567_/A vssd1 vssd1 vccd1 vccd1 _07419_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08399_ _08408_/A _10756_/Q vssd1 vssd1 vccd1 vccd1 _08399_/X sky130_fd_sc_hd__or2_1
X_10430_ _10495_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__nand2_2
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10361_ _08491_/X _06853_/B _10355_/X _10928_/Q vssd1 vssd1 vccd1 vccd1 _10928_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10292_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10292_/X sky130_fd_sc_hd__xor2_1
XFILLER_2_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05964__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10345__A2 _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05980__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10628_ _10811_/CLK _10628_/D vssd1 vssd1 vccd1 vccd1 _10628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10559_ _10700_/CLK _10559_/D vssd1 vssd1 vccd1 vccd1 _10559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06788__A1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06035__B _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09627__A _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05874__B _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07770_ _06864_/A _06864_/B _06863_/A vssd1 vssd1 vccd1 vccd1 _07771_/B sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_52_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10819_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06721_ _06721_/A vssd1 vssd1 vccd1 vccd1 _06721_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06986__A _06997_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08162__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09440_ _10869_/Q _09408_/X _09438_/Y _09439_/X vssd1 vssd1 vccd1 vccd1 _10869_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06652_ _06702_/B _06652_/B vssd1 vssd1 vccd1 vccd1 _06893_/A sky130_fd_sc_hd__xnor2_4
X_05603_ _10558_/Q _05610_/A _10559_/Q vssd1 vssd1 vccd1 vccd1 _05604_/B sky130_fd_sc_hd__o21ai_1
X_09371_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09372_/C sky130_fd_sc_hd__nor2_1
X_06583_ _06568_/A _06459_/B _06576_/B _10973_/Q vssd1 vssd1 vccd1 vccd1 _06584_/B
+ sky130_fd_sc_hd__a22oi_1
Xclkbuf_leaf_67_clock _10981_/CLK vssd1 vssd1 vccd1 vccd1 _10980_/CLK sky130_fd_sc_hd__clkbuf_16
X_08322_ _08314_/Y _08086_/X _08157_/A _08320_/X _08321_/X vssd1 vssd1 vccd1 vccd1
+ _08323_/B sky130_fd_sc_hd__o221a_1
X_05534_ _09107_/A _10544_/Q vssd1 vssd1 vccd1 vccd1 _05652_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08253_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05465_ _07885_/A _07882_/A _07878_/A _07875_/A vssd1 vssd1 vccd1 vccd1 _05467_/C
+ sky130_fd_sc_hd__or4_1
X_07204_ _07204_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07205_/B sky130_fd_sc_hd__nand2_1
X_08184_ input19/X _08123_/X _08109_/X _08180_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08185_/B sky130_fd_sc_hd__o221a_1
XFILLER_119_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05396_ _10652_/Q _05452_/A vssd1 vssd1 vccd1 vccd1 _05397_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06226__A _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07135_ _07135_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07136_/B sky130_fd_sc_hd__nor2_1
X_07066_ _07066_/A _07066_/B vssd1 vssd1 vccd1 vccd1 _07167_/B sky130_fd_sc_hd__xnor2_2
X_06017_ _10341_/A _09124_/B _09098_/A vssd1 vssd1 vccd1 vccd1 _06023_/B sky130_fd_sc_hd__or3_4
XFILLER_0_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07968_ _08971_/B _08989_/A vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09707_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__or2_1
X_06919_ _06748_/X _06940_/B _06918_/X vssd1 vssd1 vccd1 vccd1 _06939_/B sky130_fd_sc_hd__a21oi_4
X_07899_ _07899_/A vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09638_ _09769_/A _09744_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__and3_1
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09569_ _09527_/A _09527_/B _09568_/X vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__a21bo_1
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06136__A _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05690__A1 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _10408_/X _10722_/Q _10410_/X _10411_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10941_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10344_ _10344_/A vssd1 vssd1 vccd1 vccd1 _10914_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08351__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10275_ _10940_/Q _10956_/Q vssd1 vssd1 vccd1 vccd1 _10287_/D sky130_fd_sc_hd__or2b_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07958__A0 _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08940_ _09142_/D vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_130_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08871_ _08871_/A _08871_/B vssd1 vssd1 vccd1 vccd1 _08871_/Y sky130_fd_sc_hd__nand2_1
X_07822_ _06255_/X _05455_/X _06257_/X _07821_/Y vssd1 vssd1 vccd1 vccd1 hold22/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_97_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07605__A _07708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _07753_/A _07753_/B vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08280__A1_N _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ _06885_/A _06885_/B _06642_/A vssd1 vssd1 vccd1 vccd1 _06876_/B sky130_fd_sc_hd__a21oi_2
X_07684_ _07681_/A _07681_/B _09314_/A vssd1 vssd1 vccd1 vccd1 _09329_/B sky130_fd_sc_hd__o21ba_1
XFILLER_64_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _09423_/A vssd1 vssd1 vccd1 vccd1 _09677_/B sky130_fd_sc_hd__clkinv_2
X_06635_ _06719_/B _06635_/B vssd1 vssd1 vccd1 vccd1 _06638_/A sky130_fd_sc_hd__xnor2_1
X_09354_ _09372_/A _09734_/A _09674_/A vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__or3_1
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08305_ _08305_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08306_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08436__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06566_ _06571_/B _06571_/C _06571_/A vssd1 vssd1 vccd1 vccd1 _06570_/A sky130_fd_sc_hd__a21bo_1
XFILLER_33_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05517_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05517_/X sky130_fd_sc_hd__clkbuf_1
X_09285_ _09285_/A vssd1 vssd1 vccd1 vccd1 _10862_/D sky130_fd_sc_hd__buf_2
XFILLER_21_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06497_ _06502_/B _06515_/B vssd1 vssd1 vccd1 vccd1 _06517_/C sky130_fd_sc_hd__and2_1
XFILLER_138_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08236_ _08236_/A vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__clkbuf_2
X_05448_ _10647_/Q _05525_/B _05318_/X _07925_/A _05447_/X vssd1 vssd1 vccd1 vccd1
+ _05448_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08167_ input17/X _08164_/X _08165_/X _08158_/X _08394_/A vssd1 vssd1 vccd1 vccd1
+ _08167_/X sky130_fd_sc_hd__o221a_1
XFILLER_4_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05379_ _10657_/Q _05383_/A vssd1 vssd1 vccd1 vccd1 _05380_/B sky130_fd_sc_hd__and2_1
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07118_ _07150_/A _07135_/B _07117_/X vssd1 vssd1 vccd1 vccd1 _07145_/A sky130_fd_sc_hd__o21ai_1
X_08098_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08098_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07049_ _07473_/A _07463_/B vssd1 vssd1 vccd1 vccd1 _07464_/A sky130_fd_sc_hd__nor2_1
X_10060_ _10491_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10962_ _10962_/CLK _10962_/D vssd1 vssd1 vccd1 vccd1 _10962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10893_ _10909_/CLK _10893_/D vssd1 vssd1 vccd1 vccd1 _10893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10327_ _10327_/A vssd1 vssd1 vccd1 vccd1 _10327_/Y sky130_fd_sc_hd__inv_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10258_ _10243_/A _10249_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10258_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10189_ _10931_/Q _10947_/Q vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__and2b_1
XFILLER_39_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06083__A1_N _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06420_ _06420_/A _06420_/B vssd1 vssd1 vccd1 vccd1 _06732_/B sky130_fd_sc_hd__xnor2_2
XFILLER_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06351_ _06895_/A vssd1 vssd1 vccd1 vccd1 _06365_/B sky130_fd_sc_hd__clkinv_2
X_05302_ _10663_/Q _05362_/B vssd1 vssd1 vccd1 vccd1 _05363_/A sky130_fd_sc_hd__or2_1
X_09070_ _09834_/A vssd1 vssd1 vccd1 vccd1 _09904_/A sky130_fd_sc_hd__clkbuf_2
X_06282_ _06352_/A _06352_/B vssd1 vssd1 vccd1 vccd1 _06371_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08021_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09972_ _09971_/Y _09906_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__a21o_1
X_08923_ _08927_/C _08923_/B vssd1 vssd1 vccd1 vccd1 _08923_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08356__B1 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07159__A1 _07229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08854_ _08814_/X _08852_/X _08853_/X vssd1 vssd1 vccd1 vccd1 _10820_/D sky130_fd_sc_hd__o21a_1
XFILLER_69_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05997_ _09403_/A vssd1 vssd1 vccd1 vccd1 _09090_/A sky130_fd_sc_hd__clkbuf_2
X_08785_ _08819_/A vssd1 vssd1 vccd1 vccd1 _08785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07805_ _10160_/A _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _07805_/X sky130_fd_sc_hd__and3b_1
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07736_ _07729_/A _07728_/B _07565_/B _07563_/X vssd1 vssd1 vccd1 vccd1 _07738_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10466__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07667_ _07678_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08166__A _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09406_ _10192_/A vssd1 vssd1 vccd1 vccd1 _09406_/X sky130_fd_sc_hd__buf_2
XFILLER_52_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06618_ _06618_/A _06618_/B vssd1 vssd1 vccd1 vccd1 _06618_/X sky130_fd_sc_hd__and2_1
X_07598_ _07598_/A vssd1 vssd1 vccd1 vccd1 _07598_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10846__D _10846_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06549_ _06549_/A _06549_/B vssd1 vssd1 vccd1 vccd1 _06571_/B sky130_fd_sc_hd__nor2_1
X_09337_ _09387_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__or2_2
XFILLER_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09268_ _08317_/A _07911_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09268_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06117__C _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ _07998_/A _08306_/B _08217_/X _08228_/B _06011_/X vssd1 vssd1 vccd1 vccd1
+ _08219_/X sky130_fd_sc_hd__o221a_1
XFILLER_126_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08292__C1 _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ _08209_/A _09226_/S _09203_/A _09198_/X vssd1 vssd1 vccd1 vccd1 _09199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06414__A _10905_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _10112_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _10112_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10043_ _10043_/A vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_input25_A io_wbs_m2s_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07858__C1 _07857_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10945_ _10945_/CLK _10945_/D vssd1 vssd1 vccd1 vccd1 _10945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10876_ _10878_/CLK _10876_/D vssd1 vssd1 vccd1 vccd1 _10876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05884__A1 _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06308__B _10906_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08035__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ _06037_/A _05904_/Y _05902_/Y _10686_/Q _05919_/X vssd1 vssd1 vccd1 vccd1
+ _05920_/X sky130_fd_sc_hd__o221a_1
XFILLER_100_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05851_ _05851_/A _10669_/Q _05857_/B vssd1 vssd1 vccd1 vccd1 _05852_/B sky130_fd_sc_hd__or3_1
XFILLER_67_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08570_ _08572_/B _08565_/X _08569_/Y vssd1 vssd1 vccd1 vccd1 _10776_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05782_ _10704_/Q vssd1 vssd1 vccd1 vccd1 _05782_/Y sky130_fd_sc_hd__inv_2
XFILLER_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_75_clock_A clkbuf_3_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06994__A _10909_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07521_ _07657_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07648_/B sky130_fd_sc_hd__or2_1
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07452_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07454_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09066__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07383_ _07459_/B _07748_/B _07381_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07384_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_06403_ _10976_/Q vssd1 vssd1 vccd1 vccd1 _06461_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09122_ _09113_/X _09120_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06334_ _06371_/A _06334_/B vssd1 vssd1 vccd1 vccd1 _06515_/B sky130_fd_sc_hd__xor2_2
XFILLER_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09053_ _05453_/A _08978_/A _06129_/B _08098_/A _09179_/A vssd1 vssd1 vccd1 vccd1
+ _09053_/X sky130_fd_sc_hd__o221a_1
X_06265_ _10915_/Q _10898_/Q vssd1 vssd1 vccd1 vccd1 _06558_/B sky130_fd_sc_hd__nand2_2
XFILLER_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08004_ input25/X _08002_/X _08003_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10666_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06234__A _07977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06196_ _10597_/Q vssd1 vssd1 vccd1 vccd1 _06197_/A sky130_fd_sc_hd__inv_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09955_ _09955_/A _09955_/B vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__xnor2_1
XFILLER_131_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08906_ _08889_/X _08891_/X _08896_/X _08905_/X vssd1 vssd1 vccd1 vccd1 _08907_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09886_ _09956_/B _09886_/B vssd1 vssd1 vccd1 vccd1 _09887_/B sky130_fd_sc_hd__xnor2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08837_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09280__A _09280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08768_ _06187_/X _08694_/X _08695_/X _10810_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08768_/X sky130_fd_sc_hd__o221a_1
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08699_ _10803_/Q _08732_/B vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__and2_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07719_ _07391_/A _07391_/B _07588_/B _07596_/A _07718_/Y vssd1 vssd1 vccd1 vccd1
+ _07720_/B sky130_fd_sc_hd__a32o_1
X_10730_ _10768_/CLK _10730_/D vssd1 vssd1 vccd1 vccd1 _10730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10661_ _10695_/CLK _10661_/D vssd1 vssd1 vccd1 vccd1 _10661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10592_ _10958_/CLK _10592_/D vssd1 vssd1 vccd1 vccd1 _10592_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05967__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput52 _10581_/Q vssd1 vssd1 vccd1 vccd1 io_motor_irq sky130_fd_sc_hd__buf_2
Xoutput74 _10860_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[26] sky130_fd_sc_hd__buf_2
Xoutput85 _10841_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_122_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput63 _10850_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[16] sky130_fd_sc_hd__buf_2
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10928_ _10930_/CLK _10928_/D vssd1 vssd1 vccd1 vccd1 _10928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ _10862_/CLK _10859_/D vssd1 vssd1 vccd1 vccd1 _10859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08534__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08271__A2 _08212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06050_ _10655_/Q vssd1 vssd1 vccd1 vccd1 _06050_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _09930_/C vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06952_ _06952_/A _06952_/B vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__nor2_1
.ends

