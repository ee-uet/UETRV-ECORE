* NGSPICE file created from Motor_Top.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

.subckt Motor_Top clock io_ba_match io_motor_irq io_pwm_high io_pwm_low io_qei_ch_a
+ io_qei_ch_b io_wbs_ack_o io_wbs_data_o[0] io_wbs_data_o[10] io_wbs_data_o[11] io_wbs_data_o[12]
+ io_wbs_data_o[13] io_wbs_data_o[14] io_wbs_data_o[15] io_wbs_data_o[16] io_wbs_data_o[17]
+ io_wbs_data_o[18] io_wbs_data_o[19] io_wbs_data_o[1] io_wbs_data_o[20] io_wbs_data_o[21]
+ io_wbs_data_o[22] io_wbs_data_o[23] io_wbs_data_o[24] io_wbs_data_o[25] io_wbs_data_o[26]
+ io_wbs_data_o[27] io_wbs_data_o[28] io_wbs_data_o[29] io_wbs_data_o[2] io_wbs_data_o[30]
+ io_wbs_data_o[31] io_wbs_data_o[3] io_wbs_data_o[4] io_wbs_data_o[5] io_wbs_data_o[6]
+ io_wbs_data_o[7] io_wbs_data_o[8] io_wbs_data_o[9] io_wbs_m2s_addr[0] io_wbs_m2s_addr[10]
+ io_wbs_m2s_addr[11] io_wbs_m2s_addr[12] io_wbs_m2s_addr[13] io_wbs_m2s_addr[14]
+ io_wbs_m2s_addr[15] io_wbs_m2s_addr[1] io_wbs_m2s_addr[2] io_wbs_m2s_addr[3] io_wbs_m2s_addr[4]
+ io_wbs_m2s_addr[5] io_wbs_m2s_addr[6] io_wbs_m2s_addr[7] io_wbs_m2s_addr[8] io_wbs_m2s_addr[9]
+ io_wbs_m2s_data[0] io_wbs_m2s_data[10] io_wbs_m2s_data[11] io_wbs_m2s_data[12] io_wbs_m2s_data[13]
+ io_wbs_m2s_data[14] io_wbs_m2s_data[15] io_wbs_m2s_data[16] io_wbs_m2s_data[17]
+ io_wbs_m2s_data[18] io_wbs_m2s_data[19] io_wbs_m2s_data[1] io_wbs_m2s_data[20] io_wbs_m2s_data[21]
+ io_wbs_m2s_data[22] io_wbs_m2s_data[23] io_wbs_m2s_data[24] io_wbs_m2s_data[25]
+ io_wbs_m2s_data[26] io_wbs_m2s_data[27] io_wbs_m2s_data[28] io_wbs_m2s_data[29]
+ io_wbs_m2s_data[2] io_wbs_m2s_data[30] io_wbs_m2s_data[31] io_wbs_m2s_data[3] io_wbs_m2s_data[4]
+ io_wbs_m2s_data[5] io_wbs_m2s_data[6] io_wbs_m2s_data[7] io_wbs_m2s_data[8] io_wbs_m2s_data[9]
+ io_wbs_m2s_sel[0] io_wbs_m2s_sel[1] io_wbs_m2s_sel[2] io_wbs_m2s_sel[3] io_wbs_m2s_stb
+ io_wbs_m2s_we reset vccd1 vssd1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05903_ _06038_/A _05906_/A vssd1 vssd1 vccd1 vccd1 _05904_/B sky130_fd_sc_hd__and2_1
X_09671_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__nand2_1
X_06883_ _06883_/A _06883_/B vssd1 vssd1 vccd1 vccd1 _06884_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05834_ _05834_/A _05844_/C vssd1 vssd1 vccd1 vccd1 _05838_/B sky130_fd_sc_hd__or2_1
XFILLER_94_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08622_ _10790_/Q _08617_/X _08621_/Y vssd1 vssd1 vccd1 vccd1 _10790_/D sky130_fd_sc_hd__o21a_1
XFILLER_39_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08553_ _10771_/Q _08553_/B vssd1 vssd1 vccd1 vccd1 _08554_/B sky130_fd_sc_hd__xor2_1
X_05765_ _05750_/X _05765_/B _05765_/C _05765_/D vssd1 vssd1 vccd1 vccd1 _05787_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_36_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07504_ _07504_/A _07504_/B _07535_/A vssd1 vssd1 vccd1 vccd1 _07505_/B sky130_fd_sc_hd__or3_1
X_08484_ _08484_/A vssd1 vssd1 vccd1 vccd1 _10744_/D sky130_fd_sc_hd__clkbuf_1
X_05696_ _08173_/A _10552_/Q _05694_/Y _08160_/A vssd1 vssd1 vccd1 vccd1 _05798_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07435_ _07727_/A _07713_/A _07728_/B _07729_/B vssd1 vssd1 vccd1 vccd1 _07714_/S
+ sky130_fd_sc_hd__nand4_1
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09039__B2 _05733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07366_ _07366_/A _07366_/B _07366_/C vssd1 vssd1 vccd1 vccd1 _07367_/B sky130_fd_sc_hd__and3_1
XFILLER_148_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06317_ _06317_/A _06317_/B vssd1 vssd1 vccd1 vccd1 _06729_/A sky130_fd_sc_hd__nand2_2
X_09105_ _05462_/A _09148_/A _07969_/A _09104_/Y vssd1 vssd1 vccd1 vccd1 _09105_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07297_ _07310_/A _07297_/B vssd1 vssd1 vccd1 vccd1 _07298_/C sky130_fd_sc_hd__xnor2_1
X_09036_ _09209_/B vssd1 vssd1 vccd1 vccd1 _09036_/X sky130_fd_sc_hd__clkbuf_2
X_06248_ input36/X _06238_/X _06246_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10612_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06179_ _10593_/Q vssd1 vssd1 vccd1 vccd1 _06180_/A sky130_fd_sc_hd__inv_2
XANTENNA__10357__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09275__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09938_ _10482_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _09940_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09869_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09933_/A sky130_fd_sc_hd__o21ai_2
XFILLER_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09214__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10713_ _10804_/CLK _10713_/D vssd1 vssd1 vccd1 vccd1 _10713_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08238__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10644_ _10865_/CLK _10644_/D vssd1 vssd1 vccd1 vccd1 _10644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10575_ _10651_/CLK _10575_/D vssd1 vssd1 vccd1 vccd1 _10575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output56_A _10834_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__and3_1
XFILLER_37_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10520__B1 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05550_ _10548_/Q _05629_/B vssd1 vssd1 vccd1 vccd1 _05630_/A sky130_fd_sc_hd__or2_1
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05481_ _05912_/B _05470_/B _05495_/A _08994_/A _05480_/Y vssd1 vssd1 vccd1 vccd1
+ _10542_/D sky130_fd_sc_hd__a221o_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07220_ _07102_/A _07215_/B _07249_/B _07248_/A vssd1 vssd1 vccd1 vccd1 _07242_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_60_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05888__A _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07151_ _07151_/A _07394_/A _07151_/C vssd1 vssd1 vccd1 vccd1 _07322_/A sky130_fd_sc_hd__and3_1
XFILLER_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06102_ _10695_/Q _08208_/B vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__or2_1
XFILLER_157_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07082_ _09356_/A _07060_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _07083_/B sky130_fd_sc_hd__o21ai_2
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06033_ _08096_/A vssd1 vssd1 vccd1 vccd1 _06033_/X sky130_fd_sc_hd__buf_4
XFILLER_161_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07984_ _08015_/A vssd1 vssd1 vccd1 vccd1 _07985_/B sky130_fd_sc_hd__clkbuf_4
X_09723_ _09723_/A _09723_/B _09723_/C vssd1 vssd1 vccd1 vccd1 _09723_/Y sky130_fd_sc_hd__nand3_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06935_ _06935_/A _06935_/B vssd1 vssd1 vccd1 vccd1 _07609_/A sky130_fd_sc_hd__xnor2_4
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09654_ _09867_/A _09717_/A vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06866_ _06867_/B _06866_/B vssd1 vssd1 vccd1 vccd1 _06868_/A sky130_fd_sc_hd__and2b_1
XFILLER_82_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08439__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _08498_/X _08617_/B _08604_/Y _08630_/A vssd1 vssd1 vccd1 vccd1 _10785_/D
+ sky130_fd_sc_hd__a211oi_1
X_05817_ _06065_/A _09078_/A _05816_/X vssd1 vssd1 vccd1 vccd1 _05909_/A sky130_fd_sc_hd__o21a_1
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09585_ _10968_/Q _09642_/A _09492_/A _10967_/Q vssd1 vssd1 vccd1 vccd1 _09587_/A
+ sky130_fd_sc_hd__a22o_1
X_06797_ _06882_/A _06836_/A vssd1 vssd1 vccd1 vccd1 _06823_/A sky130_fd_sc_hd__xnor2_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05748_ _10703_/Q vssd1 vssd1 vccd1 vccd1 _05749_/A sky130_fd_sc_hd__inv_2
X_08536_ _08624_/B vssd1 vssd1 vccd1 vccd1 _08686_/A sky130_fd_sc_hd__buf_4
XFILLER_70_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05679_ _08304_/A _05580_/X _05583_/Y _05803_/A _05678_/X vssd1 vssd1 vccd1 vccd1
+ _05679_/X sky130_fd_sc_hd__o221a_1
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08467_ _08572_/B _10739_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08468_/B sky130_fd_sc_hd__mux2_1
XFILLER_11_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07418_ _07732_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07418_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08398_ _10198_/A vssd1 vssd1 vccd1 vccd1 _08408_/A sky130_fd_sc_hd__clkbuf_1
X_07349_ _07349_/A _07349_/B _07349_/C vssd1 vssd1 vccd1 vccd1 _07350_/B sky130_fd_sc_hd__nor3_1
XANTENNA__10854__D _10854_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10360_ _08491_/X _06818_/A _10355_/X _10927_/Q vssd1 vssd1 vccd1 vccd1 _10927_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07994__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09019_ _08998_/X _09001_/X _09018_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10835_/D
+ sky130_fd_sc_hd__o31a_4
X_10291_ _10289_/X _10300_/B _10291_/S vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05964__C input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08349__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10627_ _10657_/CLK _10627_/D vssd1 vssd1 vccd1 vccd1 _10627_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08226__A2 _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06237__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10558_ _10562_/CLK _10558_/D vssd1 vssd1 vccd1 vccd1 _10558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10489_ _10489_/A _10489_/B vssd1 vssd1 vccd1 vccd1 _10489_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08531__B _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06720_ _06720_/A _06720_/B vssd1 vssd1 vccd1 vccd1 _06725_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07163__A _07415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06651_ _06648_/A _06648_/B _06654_/A vssd1 vssd1 vccd1 vccd1 _06652_/B sky130_fd_sc_hd__o21ba_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05602_ _05602_/A _05602_/B vssd1 vssd1 vccd1 vccd1 _05602_/X sky130_fd_sc_hd__and2_1
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09370_ _09606_/B _09607_/A _09369_/X vssd1 vssd1 vccd1 vccd1 _09674_/B sky130_fd_sc_hd__a21oi_2
X_06582_ _06581_/B _06581_/C _06581_/A vssd1 vssd1 vccd1 vccd1 _06593_/B sky130_fd_sc_hd__o21ai_1
XFILLER_91_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08321_ _08321_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08321_/X sky130_fd_sc_hd__or2_1
XFILLER_33_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05533_ _10545_/Q vssd1 vssd1 vccd1 vccd1 _05547_/A sky130_fd_sc_hd__inv_2
X_08252_ _08243_/A _08251_/C _05598_/X vssd1 vssd1 vccd1 vccd1 _08252_/Y sky130_fd_sc_hd__a21oi_1
X_05464_ _10647_/Q _10646_/Q _07922_/A _07919_/A vssd1 vssd1 vccd1 vccd1 _05467_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__07610__B _07706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07203_ _07204_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07205_/A sky130_fd_sc_hd__or2_1
XFILLER_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08183_ _05883_/A _08043_/A _08179_/Y _08038_/A _08182_/Y vssd1 vssd1 vccd1 vccd1
+ _08185_/A sky130_fd_sc_hd__a221o_1
X_05395_ _10576_/Q vssd1 vssd1 vccd1 vccd1 _05452_/A sky130_fd_sc_hd__inv_2
XANTENNA__06228__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07134_ _07134_/A _07134_/B vssd1 vssd1 vccd1 vccd1 _07295_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09818__A _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07065_ _09381_/A _07056_/A _07056_/B vssd1 vssd1 vccd1 vccd1 _07066_/B sky130_fd_sc_hd__a21oi_2
XFILLER_160_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06016_ input8/X _08048_/A vssd1 vssd1 vccd1 vccd1 _09098_/A sky130_fd_sc_hd__or2_1
XFILLER_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07967_ _07967_/A _09013_/A vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09706_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__nand2_1
X_06918_ _10515_/A _07682_/B _06918_/C vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__and3_1
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07898_ _07898_/A _07898_/B vssd1 vssd1 vccd1 vccd1 _10638_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08153__A1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08153__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09637_ _09834_/B _09692_/A vssd1 vssd1 vccd1 vccd1 _09647_/A sky130_fd_sc_hd__and2_2
XFILLER_83_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10849__D _10849_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06849_ _06900_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _06860_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09568_ _09568_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _09568_/X sky130_fd_sc_hd__or2b_1
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08519_ _10797_/Q _08514_/X _08517_/X _10760_/Q vssd1 vssd1 vccd1 vccd1 _10760_/D
+ sky130_fd_sc_hd__a22o_1
X_09499_ _09542_/B _09499_/B _09499_/C vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__nand3_1
XFILLER_24_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06417__A _09356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07947__S _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06219__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10412_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09447__B _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10343_ _10343_/A _10343_/B vssd1 vssd1 vccd1 vccd1 _10344_/A sky130_fd_sc_hd__and2_1
XFILLER_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05978__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10274_ _10956_/Q _10940_/Q vssd1 vssd1 vccd1 vccd1 _10287_/C sky130_fd_sc_hd__or2b_1
XANTENNA__06152__A _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05991__A _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10402__A _10939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07958__A1 _08119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08870_ _08844_/A _08870_/B _08870_/C _08870_/D vssd1 vssd1 vccd1 vccd1 _08871_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_97_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06997__A _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07821_ _06151_/A _06258_/X _07807_/X _07820_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07821_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07752_ _07586_/A _07586_/B _07751_/X vssd1 vssd1 vccd1 vccd1 _07753_/B sky130_fd_sc_hd__o21ai_1
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06703_ _06893_/A _06893_/B _06702_/X vssd1 vssd1 vccd1 vccd1 _06885_/B sky130_fd_sc_hd__a21o_2
XFILLER_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07683_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__and2_1
X_09422_ _09422_/A _09422_/B vssd1 vssd1 vccd1 vccd1 _09423_/A sky130_fd_sc_hd__xnor2_1
X_06634_ _06634_/A _06634_/B vssd1 vssd1 vccd1 vccd1 _06635_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09353_ _09371_/B _09353_/B vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__or2_1
X_06565_ _06564_/A _06564_/B _06584_/A vssd1 vssd1 vccd1 vccd1 _06571_/A sky130_fd_sc_hd__o21ai_1
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08304_ _08304_/A vssd1 vssd1 vccd1 vccd1 _08305_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05516_ _05337_/B _05510_/X _05513_/X _07903_/A vssd1 vssd1 vccd1 vccd1 _10565_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09284_ _09289_/A _09284_/B vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__and2_2
X_06496_ _06496_/A vssd1 vssd1 vccd1 vccd1 _06521_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05447_ _07922_/A _05324_/X _05318_/X _07925_/A _05446_/X vssd1 vssd1 vccd1 vccd1
+ _05447_/X sky130_fd_sc_hd__o221a_1
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08235_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05378_ _10658_/Q _05380_/A vssd1 vssd1 vccd1 vccd1 _05378_/Y sky130_fd_sc_hd__xnor2_1
X_08166_ _08166_/A vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__buf_4
XFILLER_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07117_ _10984_/Q _07125_/A _07222_/B _10983_/Q vssd1 vssd1 vccd1 vccd1 _07117_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ _08092_/X _08094_/X _08105_/B _08096_/X vssd1 vssd1 vccd1 vccd1 _08097_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07048_ _07048_/A _07048_/B vssd1 vssd1 vccd1 vccd1 _07463_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10203__B_N _10933_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08999_ _09079_/A vssd1 vssd1 vccd1 vccd1 _08999_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08126__A1 _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08126__B2 _08117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05316__A _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10961_ _10962_/CLK _10961_/D vssd1 vssd1 vccd1 vccd1 _10961_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10892_ _10909_/CLK _10892_/D vssd1 vssd1 vccd1 vccd1 _10892_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06147__A _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05986__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10704_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10326_ _10325_/X _10318_/Y _10316_/B vssd1 vssd1 vccd1 vccd1 _10327_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10652_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _10257_/A _10257_/B vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10188_ _07539_/A _10043_/A _10184_/X _10897_/Q vssd1 vssd1 vccd1 vccd1 _10897_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06350_ _06457_/A vssd1 vssd1 vccd1 vccd1 _06895_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05301_ _07991_/A _05369_/A vssd1 vssd1 vccd1 vccd1 _05362_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06281_ _06338_/A _06281_/B vssd1 vssd1 vccd1 vccd1 _06352_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08020_ input32/X _08015_/X _08018_/Y _08019_/X vssd1 vssd1 vccd1 vccd1 _10672_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_71_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09971_ _09971_/A vssd1 vssd1 vccd1 vccd1 _09971_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _08927_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07159__A2 _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08853_ input29/X _08785_/X _08786_/X _10820_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08853_/X sky130_fd_sc_hd__o221a_1
XFILLER_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07804_ _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _07804_/Y sky130_fd_sc_hd__nor2_1
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08784_ _08773_/A _08778_/B _08803_/B _08688_/A vssd1 vssd1 vccd1 vccd1 _08784_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08108__A1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05996_ _08201_/A vssd1 vssd1 vccd1 vccd1 _09403_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08108__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07735_ _07735_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__xnor2_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__nand2_2
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _09757_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09405_/X sky130_fd_sc_hd__or2_1
XFILLER_164_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06617_ _06672_/A _06672_/B _06616_/Y vssd1 vssd1 vccd1 vccd1 _06668_/B sky130_fd_sc_hd__a21o_1
XFILLER_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07597_ _07751_/A _07597_/B vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__xor2_2
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09336_ _09336_/A _09336_/B vssd1 vssd1 vccd1 vccd1 _09417_/A sky130_fd_sc_hd__xor2_2
X_06548_ _06567_/A _06547_/C _06567_/B _06568_/A vssd1 vssd1 vccd1 vccd1 _06549_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_166_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09267_ _09267_/A vssd1 vssd1 vccd1 vccd1 _10859_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08292__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06479_ _06479_/A _06479_/B vssd1 vssd1 vccd1 vccd1 _06480_/B sky130_fd_sc_hd__and2_1
XFILLER_126_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08218_ _08218_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08228_/B sky130_fd_sc_hd__nor2_1
XFILLER_166_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _07871_/A _09136_/A _09148_/A _08208_/A _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09198_/X sky130_fd_sc_hd__a221o_1
XFILLER_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08149_ _08169_/C vssd1 vssd1 vccd1 vccd1 _08149_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08910__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10111_ _10039_/Y _10042_/B _10040_/A vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__a21o_1
XFILLER_1_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10042_ _10042_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10042_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input18_A io_wbs_m2s_data[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10944_ _10945_/CLK _10944_/D vssd1 vssd1 vccd1 vccd1 _10944_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__08357__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10875_ _10879_/CLK _10875_/D vssd1 vssd1 vccd1 vccd1 _10875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08283__B1 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08092__A _08092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ _10309_/A vssd1 vssd1 vccd1 vccd1 _10309_/Y sky130_fd_sc_hd__inv_2
XFILLER_113_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08338__A1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05850_ _10668_/Q _05863_/B vssd1 vssd1 vccd1 vccd1 _05857_/B sky130_fd_sc_hd__or2_1
XFILLER_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05781_ _08315_/B vssd1 vssd1 vccd1 vccd1 _05781_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07520_ _07661_/A _07668_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__or3_1
XANTENNA__08267__A _08267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07451_ _07598_/A _07451_/B vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__xor2_1
XFILLER_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06402_ _06441_/B _06409_/B vssd1 vssd1 vccd1 vccd1 _06690_/A sky130_fd_sc_hd__and2_2
X_07382_ _07382_/A vssd1 vssd1 vccd1 vccd1 _09304_/A sky130_fd_sc_hd__inv_2
XFILLER_148_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09121_ _10518_/B vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__clkbuf_2
X_06333_ _06371_/B _06371_/C _06804_/A vssd1 vssd1 vccd1 vccd1 _06334_/B sky130_fd_sc_hd__o21a_1
XFILLER_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06264_ _10917_/Q _10900_/Q vssd1 vssd1 vccd1 vccd1 _06270_/A sky130_fd_sc_hd__nand2_1
X_09052_ _10716_/Q _08999_/X _09037_/Y _08701_/A vssd1 vssd1 vccd1 vccd1 _09052_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08003_ _08235_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08003_/X sky130_fd_sc_hd__or2_1
XFILLER_129_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06195_ input20/X vssd1 vssd1 vccd1 vccd1 _06195_/X sky130_fd_sc_hd__buf_4
XFILLER_132_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10384__A1 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09954_ _09953_/Y _09878_/B _09882_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09955_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08905_ hold12/A _10825_/Q _10824_/Q _08876_/A _08902_/B vssd1 vssd1 vccd1 vccd1
+ _08905_/X sky130_fd_sc_hd__o41a_1
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _09883_/Y _09809_/B _09884_/X vssd1 vssd1 vccd1 vccd1 _09886_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__10136__A1 _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08825_/A _08828_/Y _08841_/C _08688_/A vssd1 vssd1 vccd1 vccd1 _08836_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08767_ _08758_/A _08761_/Y _08804_/C _08688_/A vssd1 vssd1 vccd1 vccd1 _08767_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05979_ _05958_/X _05975_/X _05978_/Y vssd1 vssd1 vccd1 vccd1 _10573_/D sky130_fd_sc_hd__o21a_1
XFILLER_72_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07718_ _07718_/A vssd1 vssd1 vccd1 vccd1 _07718_/Y sky130_fd_sc_hd__inv_2
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10500__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08698_ _08698_/A vssd1 vssd1 vccd1 vccd1 _08732_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _07649_/A _07649_/B vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__xnor2_1
XFILLER_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10660_ _10665_/CLK _10660_/D vssd1 vssd1 vccd1 vccd1 _10660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09319_ _09536_/B vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10591_ _10970_/CLK _10591_/D vssd1 vssd1 vccd1 vccd1 _10591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08624__B _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05967__C input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput53 _05956_/X vssd1 vssd1 vccd1 vccd1 io_pwm_high sky130_fd_sc_hd__buf_2
Xoutput64 _10851_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[17] sky130_fd_sc_hd__buf_2
XFILLER_150_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput75 _10861_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[27] sky130_fd_sc_hd__buf_2
XFILLER_1_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput86 _10842_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[8] sky130_fd_sc_hd__buf_2
XFILLER_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10025_ _10097_/A _10025_/B vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__xnor2_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10839__CLK _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10927_ _10929_/CLK _10927_/D vssd1 vssd1 vccd1 vccd1 _10927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10858_ _10858_/CLK _10858_/D vssd1 vssd1 vccd1 vccd1 _10858_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_108_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10790_/CLK _10789_/D vssd1 vssd1 vccd1 vccd1 _10789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08550__A _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07166__A _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _06951_/A _06951_/B vssd1 vssd1 vccd1 vccd1 _06952_/B sky130_fd_sc_hd__and2_1
XFILLER_67_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05902_ _08119_/A _05904_/A vssd1 vssd1 vccd1 vccd1 _05902_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09670_ _09671_/A _09671_/B vssd1 vssd1 vccd1 vccd1 _09670_/Y sky130_fd_sc_hd__nor2_1
X_06882_ _06882_/A _06882_/B vssd1 vssd1 vccd1 vccd1 _06883_/B sky130_fd_sc_hd__and2_1
XFILLER_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08621_ _10790_/Q _08617_/X _08630_/A vssd1 vssd1 vccd1 vccd1 _08621_/Y sky130_fd_sc_hd__a21oi_1
X_05833_ _10675_/Q vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08552_ _08586_/A vssd1 vssd1 vccd1 vccd1 _08583_/A sky130_fd_sc_hd__clkbuf_2
X_05764_ _05764_/A _05791_/A _05789_/A vssd1 vssd1 vccd1 vccd1 _05765_/D sky130_fd_sc_hd__and3_1
X_07503_ _07503_/A vssd1 vssd1 vccd1 vccd1 _07606_/A sky130_fd_sc_hd__inv_2
X_08483_ _08483_/A _08483_/B vssd1 vssd1 vccd1 vccd1 _08484_/A sky130_fd_sc_hd__and2_1
XFILLER_51_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08495__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05695_ _08169_/B vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__buf_2
XFILLER_62_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07434_ _07434_/A vssd1 vssd1 vccd1 vccd1 _07729_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07365_ _07366_/A _07366_/B _07366_/C vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__a21oi_1
XFILLER_149_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09104_ _09104_/A _09104_/B vssd1 vssd1 vccd1 vccd1 _09104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06316_ _10925_/Q _10908_/Q vssd1 vssd1 vccd1 vccd1 _06317_/B sky130_fd_sc_hd__or2_1
XFILLER_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07296_ _07296_/A _07296_/B vssd1 vssd1 vccd1 vccd1 _07297_/B sky130_fd_sc_hd__or2_1
XFILLER_164_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09035_ _09037_/A _09035_/B _09211_/B vssd1 vssd1 vccd1 vccd1 _09209_/B sky130_fd_sc_hd__or3_2
X_06247_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06247_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06178_ input47/X vssd1 vssd1 vccd1 vccd1 _06178_/X sky130_fd_sc_hd__buf_4
XFILLER_104_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08970__A1 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _09937_/A vssd1 vssd1 vccd1 vccd1 _10123_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _09868_/A _09868_/B vssd1 vssd1 vccd1 vccd1 _09870_/C sky130_fd_sc_hd__nor2_1
XFILLER_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _08819_/A vssd1 vssd1 vccd1 vccd1 _08819_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__07804__A _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09859_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09937_/A sky130_fd_sc_hd__xnor2_4
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08619__B _08649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ _10804_/CLK _10712_/D vssd1 vssd1 vccd1 vccd1 _10712_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10643_ _10643_/CLK _10643_/D vssd1 vssd1 vccd1 vccd1 _10643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10574_ _10651_/CLK _10574_/D vssd1 vssd1 vccd1 vccd1 _10574_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05994__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08370__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07749__C1 _07393_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10405__A _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08961__B2 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05775__A1 _06113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10008_ _10009_/A _10009_/B _10009_/C vssd1 vssd1 vccd1 vccd1 _10081_/A sky130_fd_sc_hd__a21oi_1
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10140__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05480_ _05480_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07150_ _07150_/A _07150_/B vssd1 vssd1 vccd1 vccd1 _07151_/C sky130_fd_sc_hd__xnor2_1
XFILLER_157_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06101_ _10694_/Q _10693_/Q _08191_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__or3_1
XFILLER_173_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07081_ _07149_/C vssd1 vssd1 vccd1 vccd1 _07326_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06032_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__buf_2
XFILLER_161_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07983_ _07983_/A vssd1 vssd1 vccd1 vccd1 _08015_/A sky130_fd_sc_hd__buf_2
XFILLER_141_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09722_ _09723_/A _09723_/B _09723_/C vssd1 vssd1 vccd1 vccd1 _09724_/A sky130_fd_sc_hd__a21oi_1
X_06934_ _06934_/A _06934_/B vssd1 vssd1 vccd1 vccd1 _06966_/A sky130_fd_sc_hd__xor2_4
X_09653_ _09653_/A _09600_/A vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__or2b_1
X_06865_ _06821_/A _06821_/B _06824_/A vssd1 vssd1 vccd1 vccd1 _06866_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08604_ _08600_/X _08597_/B _08498_/X vssd1 vssd1 vccd1 vccd1 _08604_/Y sky130_fd_sc_hd__a21oi_1
X_05816_ _06065_/A _05454_/A _05911_/A vssd1 vssd1 vccd1 vccd1 _05816_/X sky130_fd_sc_hd__a21o_1
X_09584_ _09767_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09594_/A sky130_fd_sc_hd__or2_1
XFILLER_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06796_ _06796_/A _06796_/B vssd1 vssd1 vccd1 vccd1 _06836_/A sky130_fd_sc_hd__xor2_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10291_/S sky130_fd_sc_hd__buf_2
X_05747_ _08282_/A _10563_/Q _10562_/Q _05746_/Y vssd1 vssd1 vccd1 vccd1 _05747_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08466_ _10776_/Q vssd1 vssd1 vccd1 vccd1 _08572_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05678_ _05771_/A _05588_/X _05580_/X _08304_/A _05677_/X vssd1 vssd1 vccd1 vccd1
+ _05678_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07417_ _07417_/A vssd1 vssd1 vccd1 vccd1 _07713_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08397_ _08419_/A vssd1 vssd1 vccd1 vccd1 _08397_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07348_ _07489_/A _07481_/B vssd1 vssd1 vccd1 vccd1 _07482_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07443__A1 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07443__B2 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07279_ _07302_/A _07279_/B _07344_/A vssd1 vssd1 vccd1 vccd1 _07289_/A sky130_fd_sc_hd__nor3_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09018_ _07442_/X _09015_/X _10537_/C vssd1 vssd1 vccd1 vccd1 _09018_/X sky130_fd_sc_hd__mux2_1
X_10290_ _10287_/D _10278_/Y _10287_/C vssd1 vssd1 vccd1 vccd1 _10300_/B sky130_fd_sc_hd__a21bo_1
XFILLER_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08171__A2 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05989__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10626_ _10657_/CLK _10626_/D vssd1 vssd1 vccd1 vccd1 _10626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10557_ _10562_/CLK _10557_/D vssd1 vssd1 vccd1 vccd1 _10557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10488_ _05958_/X _10475_/X _10487_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10967_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06650_ _06650_/A _06650_/B _06650_/C vssd1 vssd1 vccd1 vccd1 _06654_/A sky130_fd_sc_hd__and3_1
XFILLER_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05601_ _10560_/Q _05604_/A vssd1 vssd1 vccd1 vccd1 _05602_/B sky130_fd_sc_hd__nand2_1
XFILLER_92_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06581_ _06581_/A _06581_/B _06581_/C vssd1 vssd1 vccd1 vccd1 _06593_/A sky130_fd_sc_hd__or3_1
XFILLER_91_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08320_ _08263_/A _08327_/B _08316_/Y _08319_/X _08062_/X vssd1 vssd1 vccd1 vccd1
+ _08320_/X sky130_fd_sc_hd__o32a_1
X_05532_ _10547_/Q vssd1 vssd1 vccd1 vccd1 _05549_/A sky130_fd_sc_hd__inv_2
XFILLER_33_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08251_ _08251_/A _08251_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08277_/C sky130_fd_sc_hd__and3_1
X_05463_ _07914_/A _07911_/A _07907_/A _07903_/A vssd1 vssd1 vccd1 vccd1 _05467_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_119_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07202_ _07201_/Y _07187_/B _07190_/A vssd1 vssd1 vccd1 vccd1 _07204_/B sky130_fd_sc_hd__a21oi_1
XFILLER_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08182_ _08263_/A _08180_/Y _08189_/B _08258_/A vssd1 vssd1 vccd1 vccd1 _08182_/Y
+ sky130_fd_sc_hd__o31ai_1
X_05394_ _10621_/Q vssd1 vssd1 vccd1 vccd1 _05462_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_146_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07133_ _07133_/A _07133_/B vssd1 vssd1 vccd1 vccd1 _07134_/B sky130_fd_sc_hd__nor2_1
XFILLER_118_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07064_ _10984_/Q vssd1 vssd1 vccd1 vccd1 _07149_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_134_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06015_ input7/X _07967_/A input4/X input9/X vssd1 vssd1 vccd1 vccd1 _08048_/A sky130_fd_sc_hd__or4b_1
XANTENNA__08925__A1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07966_ _08414_/A _08939_/C vssd1 vssd1 vccd1 vccd1 _08971_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09705_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09707_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06917_ _06917_/A _06918_/C vssd1 vssd1 vccd1 vccd1 _06940_/B sky130_fd_sc_hd__xnor2_2
X_07897_ _10606_/Q _07888_/X _07892_/X _07896_/Y vssd1 vssd1 vccd1 vccd1 _07898_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09689_/A sky130_fd_sc_hd__xor2_4
X_06848_ _06848_/A _06848_/B vssd1 vssd1 vccd1 vccd1 _06862_/A sky130_fd_sc_hd__xnor2_1
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_66_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09567_ _09567_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09570_/A sky130_fd_sc_hd__xor2_1
XFILLER_128_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06779_ _06779_/A _06779_/B vssd1 vssd1 vccd1 vccd1 _06781_/B sky130_fd_sc_hd__xnor2_1
XFILLER_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08518_ _10796_/Q _08514_/X _08517_/X _10759_/Q vssd1 vssd1 vccd1 vccd1 _10759_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09498_ _09458_/A _09458_/C _09458_/B vssd1 vssd1 vccd1 vccd1 _09499_/C sky130_fd_sc_hd__a21bo_1
XFILLER_23_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ _10771_/Q _10734_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08450_/B sky130_fd_sc_hd__mux2_1
XFILLER_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10411_ _06182_/X _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10411_/X sky130_fd_sc_hd__a21bo_1
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10342_ input16/X _10415_/A _10342_/S vssd1 vssd1 vccd1 vccd1 _10343_/B sky130_fd_sc_hd__mux2_1
XFILLER_152_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10273_ _06997_/B _10115_/X _10271_/X _10272_/Y vssd1 vssd1 vccd1 vccd1 _10906_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08916__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input48_A io_wbs_m2s_sel[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08301__C1 _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06327__B _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10609_ _10643_/CLK _10609_/D vssd1 vssd1 vccd1 vccd1 _10609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_156_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07820_ _10869_/Q _07824_/B vssd1 vssd1 vccd1 vccd1 _07820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_111_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07751_ _07751_/A _07597_/B vssd1 vssd1 vccd1 vccd1 _07751_/X sky130_fd_sc_hd__or2b_1
XFILLER_38_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06702_ _06652_/B _06702_/B vssd1 vssd1 vccd1 vccd1 _06702_/X sky130_fd_sc_hd__and2b_1
X_07682_ _07682_/A _07682_/B _09303_/B vssd1 vssd1 vccd1 vccd1 _09313_/B sky130_fd_sc_hd__and3_2
XANTENNA__06146__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09422_/B sky130_fd_sc_hd__nor2_1
X_06633_ _06633_/A _06633_/B vssd1 vssd1 vccd1 vccd1 _06634_/B sky130_fd_sc_hd__or2_1
X_09352_ _10906_/Q _10890_/Q vssd1 vssd1 vccd1 vccd1 _09353_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07621__B _07702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06564_ _06564_/A _06564_/B _06584_/A vssd1 vssd1 vccd1 vccd1 _06571_/C sky130_fd_sc_hd__or3_1
XFILLER_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08303_ _08303_/A vssd1 vssd1 vccd1 vccd1 _10704_/D sky130_fd_sc_hd__clkbuf_1
X_05515_ _05340_/X _05510_/X _05513_/X _07900_/A vssd1 vssd1 vccd1 vccd1 _10564_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09283_ hold1/X _09274_/X _09275_/X _09282_/X _09270_/X vssd1 vssd1 vccd1 vccd1 _09284_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06495_ _06502_/B _06502_/C vssd1 vssd1 vccd1 vccd1 _06496_/A sky130_fd_sc_hd__and2_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08234_ _08228_/A _08228_/B _08232_/A vssd1 vssd1 vccd1 vccd1 _08234_/X sky130_fd_sc_hd__a21o_1
X_05446_ _07919_/A _05326_/X _05324_/X _10645_/Q _05445_/X vssd1 vssd1 vccd1 vccd1
+ _05446_/X sky130_fd_sc_hd__a221o_1
XFILLER_165_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08733__A _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08165_ _08355_/B vssd1 vssd1 vccd1 vccd1 _08165_/X sky130_fd_sc_hd__clkbuf_2
X_05377_ _06039_/A _05383_/A vssd1 vssd1 vccd1 vccd1 _05380_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07116_ _10984_/Q _07229_/B vssd1 vssd1 vccd1 vccd1 _07135_/B sky130_fd_sc_hd__nand2_1
X_08096_ _08096_/A vssd1 vssd1 vccd1 vccd1 _08096_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07047_ _07472_/A _07472_/B vssd1 vssd1 vccd1 vccd1 _07473_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08998_ _08062_/X _08972_/X _08974_/X _08997_/X vssd1 vssd1 vccd1 vccd1 _08998_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__07084__A _07169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _07949_/A vssd1 vssd1 vccd1 vccd1 _10651_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10960_ _10962_/CLK _10960_/D vssd1 vssd1 vccd1 vccd1 _10960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09619_ _09619_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09620_/B sky130_fd_sc_hd__xnor2_1
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10891_ _10926_/CLK _10891_/D vssd1 vssd1 vccd1 vccd1 _10891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09087__A0 _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05986__B input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06163__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06073__B1 _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10325_ _10944_/Q _10960_/Q vssd1 vssd1 vccd1 vccd1 _10325_/X sky130_fd_sc_hd__or2b_1
XFILLER_98_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09474__A _09475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10256_ _10954_/Q _10938_/Q vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__and2b_1
XFILLER_106_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07706__B _07706_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10187_ _09379_/B _10181_/X _10184_/X _10896_/Q vssd1 vssd1 vccd1 vccd1 _10896_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06983__D _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05300_ _10661_/Q _10660_/Q _05886_/A vssd1 vssd1 vccd1 vccd1 _05369_/A sky130_fd_sc_hd__nor3_2
X_06280_ _06558_/B _06360_/A vssd1 vssd1 vccd1 vccd1 _06281_/B sky130_fd_sc_hd__xor2_2
XFILLER_147_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07169__A _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06064__B1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09983_/A sky130_fd_sc_hd__or2_1
XFILLER_171_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ _08921_/A _08921_/B vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__nor2_1
XFILLER_143_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06801__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08356__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _08870_/B _08852_/B vssd1 vssd1 vccd1 vccd1 _08852_/X sky130_fd_sc_hd__xor2_1
XFILLER_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07616__B _09898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07803_ _07803_/A _07803_/B vssd1 vssd1 vccd1 vccd1 _10117_/B sky130_fd_sc_hd__xnor2_4
X_08783_ _08773_/A _08778_/B _08803_/B vssd1 vssd1 vccd1 vccd1 _08783_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05995_ input51/X vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__inv_4
XFILLER_73_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07734_ _07734_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07735_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07632__A _07715_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07665_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__or2_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ _09402_/A _09402_/B _09402_/C vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__a21oi_1
X_06616_ _06616_/A _06616_/B vssd1 vssd1 vccd1 vccd1 _06616_/Y sky130_fd_sc_hd__nor2_1
X_07596_ _07596_/A _07718_/A vssd1 vssd1 vccd1 vccd1 _07597_/B sky130_fd_sc_hd__xnor2_2
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09335_ _09316_/A _09337_/B _09334_/X vssd1 vssd1 vccd1 vccd1 _09336_/B sky130_fd_sc_hd__o21ai_2
X_06547_ _06568_/A _10973_/Q _06547_/C _06567_/B vssd1 vssd1 vccd1 vccd1 _06549_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09266_ _09289_/A _09266_/B vssd1 vssd1 vccd1 vccd1 _09267_/A sky130_fd_sc_hd__and2_2
XANTENNA__08292__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06478_ _06478_/A _06478_/B vssd1 vssd1 vccd1 vccd1 _06480_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08292__B2 _08287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08217_ _08216_/X _08218_/B _08058_/A vssd1 vssd1 vccd1 vccd1 _08217_/X sky130_fd_sc_hd__a21bo_1
X_05429_ _07882_/A _05353_/X _05350_/X _10635_/Q _05428_/X vssd1 vssd1 vccd1 vccd1
+ _05429_/X sky130_fd_sc_hd__a221o_1
XFILLER_154_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09197_ _09113_/A _09196_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08148_ _08148_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08169_/C sky130_fd_sc_hd__and2_1
XFILLER_135_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06055__B1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08075_/A _08075_/B _05733_/X vssd1 vssd1 vccd1 vccd1 _08079_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09294__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ _10110_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__xnor2_1
XFILLER_171_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07807__A _07850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10041_ _09964_/X _09967_/B _09965_/A vssd1 vssd1 vccd1 vccd1 _10042_/B sky130_fd_sc_hd__a21o_1
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10943_ _10958_/CLK _10943_/D vssd1 vssd1 vccd1 vccd1 _10943_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10874_ _10879_/CLK _10874_/D vssd1 vssd1 vccd1 vccd1 _10874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08035__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10308_ _10298_/A _10301_/Y _10297_/A vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__a21o_1
XFILLER_113_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output79_A _10864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ _10246_/C _10238_/X _08514_/A vssd1 vssd1 vccd1 vccd1 _10239_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_6_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05780_ _10566_/Q vssd1 vssd1 vccd1 vccd1 _05780_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07450_ _07450_/A _07551_/B vssd1 vssd1 vccd1 vccd1 _07451_/B sky130_fd_sc_hd__xor2_2
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06401_ _06845_/A _06627_/B vssd1 vssd1 vccd1 vccd1 _06630_/A sky130_fd_sc_hd__and2_1
X_07381_ _07381_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07458_/B sky130_fd_sc_hd__xnor2_1
XFILLER_148_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09120_ _09114_/X _09117_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__o21a_1
X_06332_ _06388_/A vssd1 vssd1 vccd1 vccd1 _06804_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ _09042_/X _09050_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10837_/D sky130_fd_sc_hd__o21a_2
X_06263_ _10918_/Q _10901_/Q vssd1 vssd1 vccd1 vccd1 _06263_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ _08015_/A vssd1 vssd1 vccd1 vccd1 _08002_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__08026__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06194_ _06191_/X _06183_/X _06193_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10596_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07627__A _07715_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09953_/Y sky130_fd_sc_hd__inv_2
XFILLER_103_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__nor2_1
XFILLER_100_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09812_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09884_/X sky130_fd_sc_hd__and2b_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08825_/A _08828_/Y _08841_/C vssd1 vssd1 vccd1 vccd1 _08835_/Y sky130_fd_sc_hd__a21oi_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08766_ _08758_/A _08761_/Y _08804_/C vssd1 vssd1 vccd1 vccd1 _08766_/Y sky130_fd_sc_hd__a21oi_1
X_05978_ _05286_/B _05975_/X _05977_/X vssd1 vssd1 vccd1 vccd1 _05978_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_100_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10703_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07720_/A sky130_fd_sc_hd__xnor2_2
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _08688_/X _08693_/Y _08696_/X vssd1 vssd1 vccd1 vccd1 _10802_/D sky130_fd_sc_hd__o21a_1
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07648_ _07655_/A _07648_/B vssd1 vssd1 vccd1 vccd1 _07649_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07579_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__or2_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_65_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10968_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09318_ _09443_/B vssd1 vssd1 vccd1 vccd1 _09536_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10590_ _10968_/CLK _10590_/D vssd1 vssd1 vccd1 vccd1 _10590_/Q sky130_fd_sc_hd__dfxtp_1
X_09249_ _09249_/A vssd1 vssd1 vccd1 vccd1 _10856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08017__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09214__A0 _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09736__B _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput54 _05954_/X vssd1 vssd1 vccd1 vccd1 io_pwm_low sky130_fd_sc_hd__buf_2
XFILLER_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput65 _10852_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[18] sky130_fd_sc_hd__buf_2
Xoutput76 _10862_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[28] sky130_fd_sc_hd__buf_2
Xoutput87 _10843_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[9] sky130_fd_sc_hd__buf_2
XFILLER_89_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input30_A io_wbs_m2s_data[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _09828_/B _09830_/X _10095_/B vssd1 vssd1 vccd1 vccd1 _10025_/B sky130_fd_sc_hd__a21boi_1
XFILLER_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ _10926_/CLK _10926_/D vssd1 vssd1 vccd1 vccd1 _10926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10857_ _10857_/CLK _10857_/D vssd1 vssd1 vccd1 vccd1 _10857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10788_/CLK _10788_/D vssd1 vssd1 vccd1 vccd1 _10788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10138__A _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09205__A0 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06950_ _06950_/A _06952_/A vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__xnor2_1
XFILLER_140_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05901_ _10654_/Q vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__buf_2
X_06881_ _06881_/A _06881_/B vssd1 vssd1 vccd1 vccd1 _06932_/B sky130_fd_sc_hd__xor2_4
X_08620_ _08620_/A vssd1 vssd1 vccd1 vccd1 _10789_/D sky130_fd_sc_hd__clkbuf_1
X_05832_ _08342_/A _05836_/A _05827_/Y vssd1 vssd1 vccd1 vccd1 _05947_/B sky130_fd_sc_hd__a21oi_1
XFILLER_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08278__A _08278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08551_ _10198_/A _08550_/X _08462_/A vssd1 vssd1 vccd1 vccd1 _08586_/A sky130_fd_sc_hd__a21o_1
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05763_ _08228_/A _10558_/Q _10557_/Q _05744_/Y vssd1 vssd1 vccd1 vccd1 _05789_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_63_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07502_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07503_/A sky130_fd_sc_hd__xnor2_2
XFILLER_74_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08482_ _10781_/Q _10744_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08483_/B sky130_fd_sc_hd__mux2_1
X_05694_ _10551_/Q vssd1 vssd1 vccd1 vccd1 _05694_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07910__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07433_ _07433_/A vssd1 vssd1 vccd1 vccd1 _07728_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07364_ _07410_/A _07364_/B vssd1 vssd1 vccd1 vccd1 _07366_/C sky130_fd_sc_hd__nand2_1
XFILLER_149_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ _09113_/A _09102_/X _10518_/B vssd1 vssd1 vccd1 vccd1 _09103_/Y sky130_fd_sc_hd__o21ai_1
X_06315_ _10925_/Q _09344_/B vssd1 vssd1 vccd1 vccd1 _06317_/A sky130_fd_sc_hd__nand2_1
XFILLER_149_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07295_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07296_/B sky130_fd_sc_hd__and2_1
X_09034_ _09023_/X _09025_/X _09033_/X _06137_/X vssd1 vssd1 vccd1 vccd1 _10836_/D
+ sky130_fd_sc_hd__o31a_4
X_06246_ _10612_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06246_/X sky130_fd_sc_hd__or2_1
XFILLER_164_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09747__A1 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05481__A1 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06177_ _06172_/X _06158_/X _06175_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10592_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09936_ _10009_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09572__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _09867_/A _09867_/B _09937_/A _09867_/D vssd1 vssd1 vccd1 vccd1 _09868_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_112_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08817_/A _08817_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08818_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07804__B _10117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10511__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09798_ _09432_/A _09735_/B _09735_/A vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__o21a_1
XFILLER_73_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ _06172_/X _08728_/X _08729_/X _08748_/X vssd1 vssd1 vccd1 vccd1 _08749_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10711_ _10851_/CLK _10711_/D vssd1 vssd1 vccd1 vccd1 _10711_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10642_ _10643_/CLK _10642_/D vssd1 vssd1 vccd1 vccd1 _10642_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08238__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10573_ _10651_/CLK _10573_/D vssd1 vssd1 vccd1 vccd1 _10573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10007_ _10077_/B _10007_/B vssd1 vssd1 vccd1 vccd1 _10009_/C sky130_fd_sc_hd__nand2_1
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10421__A _10944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08098__A _08098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10140__B _10140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10909_/CLK _10909_/D vssd1 vssd1 vccd1 vccd1 _10909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08229__A1 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08229__B2 _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06100_ _10692_/Q _10691_/Q _10690_/Q _08160_/B vssd1 vssd1 vccd1 vccd1 _08191_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_146_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07080_ _07070_/A _07070_/B _07298_/A vssd1 vssd1 vccd1 vccd1 _07089_/A sky130_fd_sc_hd__a21bo_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06031_ _10582_/Q vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__buf_2
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10315__B _10944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07982_ _06187_/X _07965_/X _07981_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10659_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_114_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09721_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09723_/C sky130_fd_sc_hd__xnor2_1
X_06933_ _06935_/A _06935_/B _06932_/X vssd1 vssd1 vccd1 vccd1 _06934_/B sky130_fd_sc_hd__a21o_2
XFILLER_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09652_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09662_/B sky130_fd_sc_hd__and2_1
X_06864_ _06864_/A _06864_/B vssd1 vssd1 vccd1 vccd1 _06867_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05815_ _05405_/A _05482_/X _05814_/X vssd1 vssd1 vccd1 vccd1 _05911_/A sky130_fd_sc_hd__o21ai_1
X_08603_ _08603_/A vssd1 vssd1 vccd1 vccd1 _10784_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09583_ _10969_/Q _09744_/B _09671_/A vssd1 vssd1 vccd1 vccd1 _09584_/B sky130_fd_sc_hd__a21boi_1
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06795_ _06763_/A _06763_/B _06766_/A vssd1 vssd1 vccd1 vccd1 _06796_/B sky130_fd_sc_hd__a21oi_1
XFILLER_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08534_ _10251_/S _10768_/Q _10767_/Q vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__and3_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05746_ _08277_/B vssd1 vssd1 vccd1 vccd1 _05746_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08465_ _08465_/A vssd1 vssd1 vccd1 vccd1 _10738_/D sky130_fd_sc_hd__clkbuf_1
X_05677_ _08285_/A _05590_/X _05588_/X _05771_/A _05676_/X vssd1 vssd1 vccd1 vccd1
+ _05677_/X sky130_fd_sc_hd__o221a_1
X_07416_ _07416_/A vssd1 vssd1 vccd1 vccd1 _07732_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08396_ _08383_/X _10739_/Q _08394_/X _08395_/X vssd1 vssd1 vccd1 vccd1 _10721_/D
+ sky130_fd_sc_hd__o211a_1
X_07347_ _07347_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07481_/B sky130_fd_sc_hd__xor2_1
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09567__A _09567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07278_ _07308_/A _07319_/A _07308_/C vssd1 vssd1 vccd1 vccd1 _07344_/A sky130_fd_sc_hd__o21ai_4
XFILLER_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09017_ _10523_/A vssd1 vssd1 vccd1 vccd1 _10537_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_06229_ _10605_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06229_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_62_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10506__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09919_ _10057_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _10056_/C sky130_fd_sc_hd__nand2_1
XFILLER_101_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05335__A _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10625_ _10657_/CLK _10625_/D vssd1 vssd1 vccd1 vccd1 _10625_/Q sky130_fd_sc_hd__dfxtp_1
X_10556_ _10665_/CLK _10556_/D vssd1 vssd1 vccd1 vccd1 _10556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10487_/X sky130_fd_sc_hd__or2_1
XFILLER_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05600_ _10699_/Q vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_92_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06580_ _06594_/A _06594_/B _06579_/Y vssd1 vssd1 vccd1 vccd1 _06607_/B sky130_fd_sc_hd__o21bai_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05531_ _10554_/Q vssd1 vssd1 vccd1 vccd1 _05663_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08250_ _08157_/X _08245_/Y _08247_/Y _08249_/X vssd1 vssd1 vccd1 vccd1 _10699_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05462_ _05462_/A _05462_/B _05462_/C _05462_/D vssd1 vssd1 vccd1 vccd1 _05462_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07201_ _07201_/A vssd1 vssd1 vccd1 vccd1 _07201_/Y sky130_fd_sc_hd__inv_2
X_08181_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08189_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05393_ _10621_/Q _05393_/B vssd1 vssd1 vccd1 vccd1 _05393_/X sky130_fd_sc_hd__and2_1
XFILLER_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07132_ _07132_/A _07132_/B vssd1 vssd1 vccd1 vccd1 _07285_/A sky130_fd_sc_hd__xnor2_1
XFILLER_119_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07063_ _07086_/B _07188_/B vssd1 vssd1 vccd1 vccd1 _07070_/A sky130_fd_sc_hd__and2_1
XFILLER_133_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06014_ input50/X input48/X vssd1 vssd1 vccd1 vccd1 _10341_/A sky130_fd_sc_hd__nand2_2
XANTENNA__07189__A1 _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07635__A _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07965_ _08034_/B vssd1 vssd1 vccd1 vccd1 _07965_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09704_ _09644_/A _09769_/C _09703_/X vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__o21a_1
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06916_ _06916_/A _06916_/B vssd1 vssd1 vccd1 vccd1 _06918_/C sky130_fd_sc_hd__nor2_2
XFILLER_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07896_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07896_/Y sky130_fd_sc_hd__inv_2
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09635_ _10873_/Q _09572_/X _09631_/X _09634_/Y vssd1 vssd1 vccd1 vccd1 _10873_/D
+ sky130_fd_sc_hd__a22o_1
X_06847_ _06847_/A _06847_/B vssd1 vssd1 vccd1 vccd1 _06848_/B sky130_fd_sc_hd__nor2_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09566_ _09566_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__xnor2_1
X_06778_ _06792_/A _06778_/B vssd1 vssd1 vccd1 vccd1 _06781_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08517_ _10177_/A vssd1 vssd1 vccd1 vccd1 _08517_/X sky130_fd_sc_hd__clkbuf_4
X_05729_ _10546_/Q vssd1 vssd1 vccd1 vccd1 _05729_/Y sky130_fd_sc_hd__inv_2
X_09497_ _09542_/A _09496_/C _09496_/A vssd1 vssd1 vccd1 vccd1 _09499_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08448_ _08448_/A vssd1 vssd1 vccd1 vccd1 _10733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08379_ _08367_/X _10733_/Q _07865_/X _08378_/X vssd1 vssd1 vccd1 vccd1 _10715_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10410_ _10941_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10410_/X sky130_fd_sc_hd__and2_1
XFILLER_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _10341_/A _10341_/B _10341_/C vssd1 vssd1 vccd1 vccd1 _10342_/S sky130_fd_sc_hd__or3_1
XFILLER_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10272_ _10287_/A _10271_/B _09480_/X vssd1 vssd1 vccd1 vccd1 _10272_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_105_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08377__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _10643_/CLK _10608_/D vssd1 vssd1 vccd1 vccd1 _10608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10411__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10539_ _08974_/X _08969_/Y _09036_/X _06137_/X vssd1 vssd1 vccd1 vccd1 _10987_/D
+ sky130_fd_sc_hd__o31a_2
XFILLER_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07158__C _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09654__B _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07750_ _07750_/A _07750_/B vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__xor2_1
XFILLER_38_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06701_ _06903_/A _06903_/B _06700_/X vssd1 vssd1 vccd1 vccd1 _06893_/B sky130_fd_sc_hd__a21o_2
X_07681_ _07681_/A _07681_/B vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_10_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09420_ _09420_/A _10885_/Q vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__and2_1
X_06632_ _06633_/A _06633_/B vssd1 vssd1 vccd1 vccd1 _06634_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08286__A _08287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09351_ _10890_/Q _10906_/Q vssd1 vssd1 vccd1 vccd1 _09371_/B sky130_fd_sc_hd__and2b_1
X_06563_ _10974_/Q _10973_/Q _06575_/B _06587_/A vssd1 vssd1 vccd1 vccd1 _06584_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ _08300_/X _08302_/B vssd1 vssd1 vccd1 vccd1 _08303_/A sky130_fd_sc_hd__and2b_1
X_05514_ _05343_/Y _05510_/X _05513_/X _07896_/A vssd1 vssd1 vccd1 vccd1 _10563_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09282_ _08027_/A _09281_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09282_/X sky130_fd_sc_hd__mux2_1
XFILLER_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06494_ _10971_/Q vssd1 vssd1 vccd1 vccd1 _06502_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_08233_ _08233_/A _08233_/B vssd1 vssd1 vccd1 vccd1 _08233_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05445_ _07914_/A _05329_/X _05326_/X _10644_/Q _05444_/X vssd1 vssd1 vccd1 vccd1
+ _05445_/X sky130_fd_sc_hd__o221a_1
XFILLER_165_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08164_ _08248_/A vssd1 vssd1 vccd1 vccd1 _08164_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05376_ _10626_/Q vssd1 vssd1 vccd1 vccd1 _05461_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07115_ _07222_/B vssd1 vssd1 vccd1 vccd1 _07229_/B sky130_fd_sc_hd__buf_2
XFILLER_162_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08095_ _08095_/A _08095_/B vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10056__A _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06253__B _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07046_ _07421_/A _07046_/B vssd1 vssd1 vccd1 vccd1 _07472_/B sky130_fd_sc_hd__xnor2_1
XFILLER_47_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09571__A2 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08997_ _05813_/A _08976_/X _08994_/X _08996_/Y _09078_/B vssd1 vssd1 vccd1 vccd1
+ _08997_/X sky130_fd_sc_hd__a221o_1
XFILLER_102_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07948_ _07955_/A _07948_/B vssd1 vssd1 vccd1 vccd1 _07949_/A sky130_fd_sc_hd__or2_1
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07879_ hold6/X _07870_/X _07874_/X _07878_/Y vssd1 vssd1 vccd1 vccd1 _07880_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09618_ _09618_/A _09618_/B _09618_/C vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__or3_1
XFILLER_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10890_ _10909_/CLK _10890_/D vssd1 vssd1 vccd1 vccd1 _10890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09549_ _09549_/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09610_/C sky130_fd_sc_hd__xor2_4
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08643__B _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05968__A_N input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10324_ _10324_/A _10334_/A vssd1 vssd1 vccd1 vccd1 _10330_/A sky130_fd_sc_hd__or2_1
XANTENNA__06073__B2 _08082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10255_ _10938_/Q _10954_/Q vssd1 vssd1 vccd1 vccd1 _10257_/A sky130_fd_sc_hd__and2b_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10186_ _07570_/A _10181_/X _10184_/X _10895_/Q vssd1 vssd1 vccd1 vccd1 _10895_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07869__A_N _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07169__B _07169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06064__A1 _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06064__B2 _09104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08927_/C sky130_fd_sc_hd__nand2_1
XFILLER_112_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08851_ _08847_/X _08815_/B _08845_/Y vssd1 vssd1 vccd1 vccd1 _08852_/B sky130_fd_sc_hd__a21o_1
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08210__C1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07564__A1 _07563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07802_ _07802_/A _07802_/B vssd1 vssd1 vccd1 vccd1 _07803_/B sky130_fd_sc_hd__xnor2_2
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05994_ _07880_/A _05994_/B vssd1 vssd1 vccd1 vccd1 _10576_/D sky130_fd_sc_hd__nor2_1
XFILLER_111_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08782_ _10812_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08803_/B sky130_fd_sc_hd__xor2_2
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07733_ _07733_/A _07733_/B vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07664_ _07665_/A _07665_/B vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__nand2_1
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09403_ _09403_/A _09403_/B vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__nand2_4
XFILLER_164_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06615_ _06681_/A _06674_/C _06674_/A vssd1 vssd1 vccd1 vccd1 _06672_/B sky130_fd_sc_hd__a21bo_1
X_07595_ _07397_/A _07397_/B _07594_/X vssd1 vssd1 vccd1 vccd1 _07718_/A sky130_fd_sc_hd__a21oi_2
XFILLER_34_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ _10883_/Q _07098_/A vssd1 vssd1 vccd1 vccd1 _09334_/X sky130_fd_sc_hd__or2b_1
X_06546_ _06546_/A _06602_/A vssd1 vssd1 vccd1 vccd1 _06618_/A sky130_fd_sc_hd__xnor2_2
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09265_ _10824_/Q _09243_/X _09244_/X _09264_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09266_/B sky130_fd_sc_hd__a32o_1
X_06477_ _06477_/A _06477_/B vssd1 vssd1 vccd1 vccd1 _06478_/B sky130_fd_sc_hd__and2_1
XFILLER_166_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08216_ _08218_/A vssd1 vssd1 vccd1 vccd1 _08216_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05428_ _07878_/A _05358_/X _05353_/X _10634_/Q _05427_/X vssd1 vssd1 vccd1 vccd1
+ _05428_/X sky130_fd_sc_hd__o221a_1
XFILLER_166_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09196_ _09114_/A _09195_/X _10500_/B vssd1 vssd1 vccd1 vccd1 _09196_/X sky130_fd_sc_hd__o21a_1
XFILLER_135_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ _08150_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08147_/X sky130_fd_sc_hd__or2_1
XFILLER_112_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05359_ _10632_/Q vssd1 vssd1 vccd1 vccd1 _07875_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06055__B2 _09104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08078_ _08073_/X _08076_/X _08077_/X vssd1 vssd1 vccd1 vccd1 _10682_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07029_ _07044_/A _07030_/C _07417_/A _07021_/A vssd1 vssd1 vccd1 vccd1 _07031_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ _10040_/A _10039_/Y vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__or2b_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07823__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10942_ _10942_/CLK _10942_/D vssd1 vssd1 vccd1 vccd1 _10942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10873_ _10879_/CLK _10873_/D vssd1 vssd1 vccd1 vccd1 _10873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06174__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08035__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _10307_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10424__A _10945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10238_ _10236_/X _10237_/Y _10279_/S vssd1 vssd1 vccd1 vccd1 _10238_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10169_ _07098_/A _10167_/X _08517_/X _10883_/Q vssd1 vssd1 vccd1 vccd1 _10883_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06400_ _06441_/B vssd1 vssd1 vccd1 vccd1 _06845_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_90_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07380_ _07459_/B _07490_/A _07327_/X vssd1 vssd1 vccd1 vccd1 _07381_/B sky130_fd_sc_hd__a21bo_1
XFILLER_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06331_ _06342_/A _06342_/B vssd1 vssd1 vccd1 vccd1 _06388_/A sky130_fd_sc_hd__xnor2_1
XFILLER_148_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09379__B _09379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ _10484_/A _10474_/B _10495_/B _10506_/A _09049_/X vssd1 vssd1 vccd1 vccd1
+ _09050_/X sky130_fd_sc_hd__a221o_1
X_06262_ _06262_/A _06262_/B vssd1 vssd1 vccd1 vccd1 _06305_/A sky130_fd_sc_hd__nand2_2
XFILLER_163_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08001_ input24/X _07987_/X _08000_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10665_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06193_ _06193_/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06193_/Y sky130_fd_sc_hd__nand2_1
XFILLER_156_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09952_ _09952_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__xnor2_2
XFILLER_116_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08903_ hold1/X _08919_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__nor2_1
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09883_/A vssd1 vssd1 vccd1 vccd1 _09883_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08834_ _10818_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08841_/C sky130_fd_sc_hd__xor2_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08765_ _10810_/Q _08801_/B vssd1 vssd1 vccd1 vccd1 _08804_/C sky130_fd_sc_hd__xor2_2
X_05977_ _08445_/A vssd1 vssd1 vccd1 vccd1 _05977_/X sky130_fd_sc_hd__buf_2
XFILLER_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _07442_/X _07574_/B _07715_/X vssd1 vssd1 vccd1 vccd1 _07717_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08696_ _06147_/X _08694_/X _08695_/X _10802_/Q _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08696_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07647_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _09532_/A sky130_fd_sc_hd__xnor2_4
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07578_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07580_/A sky130_fd_sc_hd__nand2_1
XFILLER_80_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _09736_/B _09388_/A vssd1 vssd1 vccd1 vccd1 _09396_/B sky130_fd_sc_hd__nand2_1
X_06529_ _06527_/A _06489_/B _06540_/A _06600_/A vssd1 vssd1 vccd1 vccd1 _06529_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _09259_/A _09248_/B vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__and2_2
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09226_/S sky130_fd_sc_hd__buf_2
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08640__C _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput55 _10987_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_ack_o sky130_fd_sc_hd__buf_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 _10853_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[19] sky130_fd_sc_hd__buf_2
Xoutput77 _10863_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[29] sky130_fd_sc_hd__buf_2
XFILLER_150_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10023_ _10023_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _10095_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08649__A _08649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input23_A io_wbs_m2s_data[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_57_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09150__B1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10925_ _10925_/CLK _10925_/D vssd1 vssd1 vccd1 vccd1 _10925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10856_ _10856_/CLK _10856_/D vssd1 vssd1 vccd1 vccd1 _10856_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08384__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ _10788_/CLK _10787_/D vssd1 vssd1 vccd1 vccd1 _10787_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07728__A _07728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05900_ _05900_/A _05900_/B vssd1 vssd1 vccd1 vccd1 _05900_/X sky130_fd_sc_hd__and2_1
XFILLER_67_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06880_ _07799_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _06934_/A sky130_fd_sc_hd__xor2_4
XFILLER_39_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08192__A1 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08192__B2 _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05831_ _08027_/A _05831_/B _05831_/C vssd1 vssd1 vccd1 vccd1 _05836_/A sky130_fd_sc_hd__or3_1
XFILLER_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05762_ _05746_/Y _10562_/Q _10561_/Q _05751_/Y _05761_/X vssd1 vssd1 vccd1 vccd1
+ _05791_/A sky130_fd_sc_hd__o221a_1
XFILLER_48_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08550_ _08661_/A vssd1 vssd1 vccd1 vccd1 _08550_/X sky130_fd_sc_hd__clkbuf_2
X_07501_ _07501_/A _07505_/A vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__and2_1
X_08481_ _08481_/A vssd1 vssd1 vccd1 vccd1 _10743_/D sky130_fd_sc_hd__clkbuf_1
X_05693_ _05693_/A vssd1 vssd1 vccd1 vccd1 _08173_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08495__A2 _08491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07432_ _07563_/A vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_161_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10974__D _10974_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07363_ _07361_/Y _07363_/B _07363_/C vssd1 vssd1 vccd1 vccd1 _07364_/B sky130_fd_sc_hd__nand3b_1
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09102_ _09114_/A _09101_/X _09118_/A vssd1 vssd1 vccd1 vccd1 _09102_/X sky130_fd_sc_hd__o21a_1
X_06314_ _10908_/Q vssd1 vssd1 vccd1 vccd1 _09344_/B sky130_fd_sc_hd__clkbuf_2
X_07294_ _07309_/A _07309_/C _07309_/B vssd1 vssd1 vccd1 vccd1 _07310_/A sky130_fd_sc_hd__a21oi_1
XFILLER_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06245_ input35/X _06238_/X _06244_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10611_/D
+ sky130_fd_sc_hd__o211a_1
X_09033_ _07726_/A _09032_/X _10537_/C vssd1 vssd1 vccd1 vccd1 _09033_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07638__A _07715_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06176_ _10343_/A vssd1 vssd1 vccd1 vccd1 _06176_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_144_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09935_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08707__B1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _09931_/A _09937_/A _10139_/S _09736_/B vssd1 vssd1 vccd1 vccd1 _09868_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08183__A1 _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08183__B2 _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ _08817_/A _08817_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08817_/X sky130_fd_sc_hd__and3_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _09797_/A _09797_/B vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__xnor2_4
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ _10807_/Q vssd1 vssd1 vccd1 vccd1 _08748_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_38_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08679_ _10801_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08679_/X sky130_fd_sc_hd__and2_1
XFILLER_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _10860_/CLK _10710_/D vssd1 vssd1 vccd1 vccd1 _10710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _10643_/CLK _10641_/D vssd1 vssd1 vccd1 vccd1 _10641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10572_ _10855_/CLK _10572_/D vssd1 vssd1 vccd1 vccd1 _10572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07997__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08174__A1 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08174__B2 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10007_/B sky130_fd_sc_hd__or2_1
XFILLER_92_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10908_ _10925_/CLK _10908_/D vssd1 vssd1 vccd1 vccd1 _10908_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10839_ _10977_/CLK _10839_/D vssd1 vssd1 vccd1 vccd1 _10839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08229__A2 _08074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07437__B1 _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09938__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06030_ _10581_/Q _06020_/X _06029_/X vssd1 vssd1 vccd1 vccd1 _10581_/D sky130_fd_sc_hd__o21a_1
XFILLER_173_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07981_ _07981_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07981_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_64_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10962_/CLK sky130_fd_sc_hd__clkbuf_16
X_09720_ _09716_/Y _09718_/Y _09719_/X vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__o21a_1
XFILLER_101_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06932_ _06890_/B _06932_/B vssd1 vssd1 vccd1 vccd1 _06932_/X sky130_fd_sc_hd__and2b_1
XFILLER_67_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08289__A _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09651_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09662_/A sky130_fd_sc_hd__nor2_1
XFILLER_110_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06863_ _06863_/A _06863_/B vssd1 vssd1 vccd1 vccd1 _06864_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08602_ _08617_/B _08649_/A _08602_/C vssd1 vssd1 vccd1 vccd1 _08603_/A sky130_fd_sc_hd__and3b_1
X_05814_ _05408_/Y _05643_/A _05813_/X vssd1 vssd1 vccd1 vccd1 _05814_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09582_ _10970_/Q _09744_/A vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__nand2_2
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06794_ _06832_/A _06794_/B vssd1 vssd1 vccd1 vccd1 _06796_/A sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_79_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10967_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__07921__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ _08881_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _10767_/D sky130_fd_sc_hd__nor2_1
X_05745_ _10702_/Q vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__clkinv_2
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08464_ _08477_/A _08464_/B vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__or2_1
X_05676_ _08277_/A _05593_/X _05590_/X _08285_/A _05675_/X vssd1 vssd1 vccd1 vccd1
+ _05676_/X sky130_fd_sc_hd__a221o_1
XFILLER_50_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07415_ _07415_/A _07472_/A _07415_/C _07434_/A vssd1 vssd1 vccd1 vccd1 _07428_/A
+ sky130_fd_sc_hd__or4b_1
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08395_ _08395_/A _10755_/Q vssd1 vssd1 vccd1 vccd1 _08395_/X sky130_fd_sc_hd__or2_1
X_07346_ _07488_/B _07529_/A _07488_/A vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__o21ai_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07277_ _07277_/A _07277_/B vssd1 vssd1 vccd1 vccd1 _07308_/C sky130_fd_sc_hd__xnor2_2
XFILLER_164_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09016_ _09016_/A _09016_/B vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__or2_1
X_06228_ input28/X _06225_/X _06227_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10604_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_124_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06159_ _10589_/Q vssd1 vssd1 vccd1 vccd1 _06160_/A sky130_fd_sc_hd__inv_2
XFILLER_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _10031_/A sky130_fd_sc_hd__xnor2_2
XFILLER_120_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09849_ _09901_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09851_/C sky130_fd_sc_hd__xor2_1
XFILLER_19_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10624_ _10655_/CLK _10624_/D vssd1 vssd1 vccd1 vccd1 _10624_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10555_ _10665_/CLK _10555_/D vssd1 vssd1 vccd1 vccd1 _10555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06182__A input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ _06147_/X _10475_/X _10484_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10966_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_154_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05530_ _10567_/Q vssd1 vssd1 vccd1 vccd1 _05769_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05461_ _05461_/A _05461_/B _05461_/C _05461_/D vssd1 vssd1 vccd1 vccd1 _05462_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_159_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07200_ _07200_/A _07200_/B vssd1 vssd1 vccd1 vccd1 _07204_/A sky130_fd_sc_hd__xnor2_1
XFILLER_159_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05392_ _05392_/A _05392_/B vssd1 vssd1 vccd1 vccd1 _05393_/B sky130_fd_sc_hd__nor2_1
X_08180_ _08180_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _08180_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07131_ _07377_/A _07229_/B _07147_/A vssd1 vssd1 vccd1 vccd1 _07132_/B sky130_fd_sc_hd__and3_1
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07062_ _07164_/B vssd1 vssd1 vccd1 vccd1 _07188_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_161_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06013_ _06008_/X _05975_/X _06012_/Y vssd1 vssd1 vccd1 vccd1 _10579_/D sky130_fd_sc_hd__o21a_1
XFILLER_173_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10193__B2 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07964_ _07964_/A vssd1 vssd1 vccd1 vccd1 _08034_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09703_ _09703_/A _09703_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__or3b_1
XFILLER_68_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06915_ _06915_/A _06915_/B _06942_/A vssd1 vssd1 vccd1 vccd1 _06916_/B sky130_fd_sc_hd__nor3_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07895_ _07898_/A _07895_/B vssd1 vssd1 vccd1 vccd1 _10637_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09634_ _09634_/A _09686_/B vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06846_ _10508_/A _07784_/B _06845_/C vssd1 vssd1 vccd1 vccd1 _06847_/B sky130_fd_sc_hd__a21oi_1
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09565_ _09625_/A _09625_/B _09626_/A vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__o21a_1
X_06777_ _06900_/A _07783_/B _06775_/C vssd1 vssd1 vccd1 vccd1 _06778_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10248__A2 _10935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08516_ _10795_/Q _08514_/X _08509_/X _10758_/Q vssd1 vssd1 vccd1 vccd1 _10758_/D
+ sky130_fd_sc_hd__a22o_1
X_05728_ _06037_/A vssd1 vssd1 vccd1 vccd1 _05728_/X sky130_fd_sc_hd__buf_2
X_09496_ _09496_/A _09542_/A _09496_/C vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__nand3_1
XFILLER_12_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08447_ _08460_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08448_/A sky130_fd_sc_hd__or2_1
X_05659_ _05896_/A _05628_/X _05626_/X _08148_/A _05658_/X vssd1 vssd1 vccd1 vccd1
+ _05659_/X sky130_fd_sc_hd__o221a_1
XFILLER_12_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08378_ _08381_/A _10749_/Q vssd1 vssd1 vccd1 vccd1 _08378_/X sky130_fd_sc_hd__or2_1
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07329_ _07562_/A _07327_/X _07511_/A _07328_/Y vssd1 vssd1 vccd1 vccd1 _07333_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10517__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10340_ _10914_/Q vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10420__A2 _10724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10271_ _10287_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10271_/X sky130_fd_sc_hd__or2_1
XFILLER_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08657__A _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07561__A _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_4_0_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__B2 _08297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_6_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 _10682_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_159_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10607_ _10643_/CLK _10607_/D vssd1 vssd1 vccd1 vccd1 _10607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10427__A _10946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10538_ _07592_/A _10522_/A _10537_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10986_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10469_ _10961_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10469_/X sky130_fd_sc_hd__or2_1
XFILLER_124_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07040__A1 _07416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10357__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07591__A2 _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06700_ _06665_/B _06700_/B vssd1 vssd1 vccd1 vccd1 _06700_/X sky130_fd_sc_hd__and2b_1
XFILLER_77_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07680_ _07680_/A _07680_/B vssd1 vssd1 vccd1 vccd1 _07681_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06631_ _06631_/A _06631_/B vssd1 vssd1 vccd1 vccd1 _06633_/B sky130_fd_sc_hd__xnor2_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09350_ _09371_/A _09372_/B vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__or2_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06562_ _06585_/A _06585_/B _06573_/C vssd1 vssd1 vccd1 vccd1 _06564_/B sky130_fd_sc_hd__and3_1
XFILLER_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08301_ input32/X _08248_/A _08052_/A _08297_/A _08175_/A vssd1 vssd1 vccd1 vccd1
+ _08302_/B sky130_fd_sc_hd__o221a_1
X_05513_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05513_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09281_ _08332_/A _07919_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09281_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06493_ _06527_/A _06513_/D _06493_/C vssd1 vssd1 vccd1 vccd1 _06510_/A sky130_fd_sc_hd__and3_1
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08251_/C sky130_fd_sc_hd__nor2_2
X_05444_ _10643_/Q _05329_/X _05438_/X _07911_/A _05443_/X vssd1 vssd1 vccd1 vccd1
+ _05444_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06815__A _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ _08158_/X _08169_/C _08162_/Y vssd1 vssd1 vccd1 vccd1 _08163_/Y sky130_fd_sc_hd__a21oi_1
X_05375_ _10627_/Q vssd1 vssd1 vccd1 vccd1 _05461_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07114_ _07216_/B vssd1 vssd1 vccd1 vccd1 _07222_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08094_ _08098_/A _08095_/B vssd1 vssd1 vccd1 vccd1 _08094_/X sky130_fd_sc_hd__or2_1
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07045_ _07573_/A _07434_/A _07509_/A vssd1 vssd1 vccd1 vccd1 _07046_/B sky130_fd_sc_hd__and3_1
XFILLER_162_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08359__A1 _05528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06550__A _10971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10166__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ _05721_/Y _06212_/B _08995_/X vssd1 vssd1 vccd1 vccd1 _08996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07947_ input41/X _05279_/A _07964_/A vssd1 vssd1 vccd1 vccd1 _07948_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07878_ _07878_/A vssd1 vssd1 vccd1 vccd1 _07878_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09617_ _09545_/B _09617_/B vssd1 vssd1 vccd1 vccd1 _09618_/C sky130_fd_sc_hd__and2b_1
XFILLER_71_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06829_ _06882_/A _06883_/A _06882_/B vssd1 vssd1 vccd1 vccd1 _06884_/A sky130_fd_sc_hd__and3_1
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09548_ _09432_/A _09508_/B _09508_/A vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__o21ai_4
XFILLER_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _09479_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09479_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10323_ _10945_/Q _10961_/Q vssd1 vssd1 vccd1 vccd1 _10334_/A sky130_fd_sc_hd__and2b_1
XANTENNA__06073__A2 _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10254_ _07061_/A _10253_/A _10253_/Y _08563_/X vssd1 vssd1 vccd1 vccd1 _10904_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10185_ _09920_/B _10181_/X _10184_/X _10894_/Q vssd1 vssd1 vccd1 vccd1 _10894_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10396__A1 _10937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06064__A2 _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08850_ _10820_/Q _08865_/B vssd1 vssd1 vccd1 vccd1 _08870_/B sky130_fd_sc_hd__xor2_1
XFILLER_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07801_ _07801_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__xnor2_1
X_08781_ _08778_/X _08779_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10811_/D sky130_fd_sc_hd__o21a_1
X_05993_ _05992_/X _09107_/A _05993_/S vssd1 vssd1 vccd1 vccd1 _05994_/B sky130_fd_sc_hd__mux2_1
XFILLER_78_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07732_ _07732_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07733_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08297__A _08297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07663_ _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07665_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10977__D _10977_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09402_ _09402_/A _09402_/B _09402_/C vssd1 vssd1 vccd1 vccd1 _09402_/X sky130_fd_sc_hd__and3_1
X_06614_ _06614_/A _06614_/B _06614_/C vssd1 vssd1 vccd1 vccd1 _06674_/A sky130_fd_sc_hd__nand3_1
XFILLER_111_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07594_ _07396_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07594_/X sky130_fd_sc_hd__and2b_1
XFILLER_81_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09333_ _09333_/A _09333_/B vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__nor2_2
X_06545_ _06545_/A _06520_/X vssd1 vssd1 vccd1 vccd1 _06546_/A sky130_fd_sc_hd__or2b_1
XFILLER_34_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09264_ _05844_/A _09262_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09264_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06476_ _06688_/A _06688_/B vssd1 vssd1 vccd1 vccd1 _06658_/A sky130_fd_sc_hd__or2b_1
XANTENNA__07679__B1_N _07519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08215_ _08215_/A vssd1 vssd1 vccd1 vccd1 _10695_/D sky130_fd_sc_hd__clkbuf_1
X_05427_ _07875_/A _05360_/X _05358_/X _10633_/Q _05426_/X vssd1 vssd1 vccd1 vccd1
+ _05427_/X sky130_fd_sc_hd__a221o_1
X_09195_ _10946_/Q _09143_/Y _09194_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09195_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_5_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09856__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08146_ _08146_/A vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__buf_2
X_05358_ _05358_/A _05358_/B vssd1 vssd1 vccd1 vccd1 _05358_/X sky130_fd_sc_hd__and2_1
XANTENNA__10387__A1 _10935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06055__A2 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08077_ _10526_/A _08047_/X _08052_/X _08075_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08077_/X sky130_fd_sc_hd__o221a_1
XFILLER_150_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05289_ _05279_/A _05454_/A _05400_/A vssd1 vssd1 vccd1 vccd1 _05289_/Y sky130_fd_sc_hd__a21oi_1
X_07028_ _07028_/A _07028_/B vssd1 vssd1 vccd1 vccd1 _07417_/A sky130_fd_sc_hd__xnor2_2
XFILLER_162_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08979_ hold10/A _09020_/B vssd1 vssd1 vccd1 vccd1 _08979_/X sky130_fd_sc_hd__or2_1
XFILLER_75_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10941_ _10945_/CLK _10941_/D vssd1 vssd1 vccd1 vccd1 _10941_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08000__A _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10872_ _10970_/CLK _10872_/D vssd1 vssd1 vccd1 vccd1 _10872_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08670__A _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_53_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ _10959_/Q _10943_/Q vssd1 vssd1 vccd1 vccd1 _10307_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08991__A1 _10799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10237_ _10225_/A _10228_/Y _10225_/B vssd1 vssd1 vccd1 vccd1 _10237_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10168_ _07394_/X _10167_/X _08517_/X _10882_/Q vssd1 vssd1 vccd1 vccd1 _10882_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10099_ _10100_/A _10100_/B _10100_/C vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__a21o_1
XANTENNA__05534__A _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06330_ _10930_/Q _07112_/A vssd1 vssd1 vccd1 vccd1 _06342_/B sky130_fd_sc_hd__xnor2_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06365__A _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06261_ _10919_/Q _10902_/Q vssd1 vssd1 vccd1 vccd1 _06262_/B sky130_fd_sc_hd__or2_1
XFILLER_117_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08000_ _08000_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08000_/X sky130_fd_sc_hd__or2_1
XFILLER_129_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06192_ _10596_/Q vssd1 vssd1 vccd1 vccd1 _06193_/A sky130_fd_sc_hd__inv_2
XFILLER_117_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08982__A1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09951_ _09671_/A _10023_/B _09949_/Y _10027_/A vssd1 vssd1 vccd1 vccd1 _09952_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_89_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08902_ hold1/X _08902_/B vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__and2_1
XFILLER_98_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _09882_/A _09882_/B vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__xor2_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07924__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ _08829_/X _08832_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10817_/D sky130_fd_sc_hd__o21a_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08762_/X _08763_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10809_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05976_ input51/X vssd1 vssd1 vccd1 vccd1 _08445_/A sky130_fd_sc_hd__buf_4
XFILLER_122_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07715_ _09379_/B _07571_/B _07715_/C _07715_/D vssd1 vssd1 vccd1 vccd1 _07715_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_66_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08695_ _08820_/A vssd1 vssd1 vccd1 vccd1 _08695_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07646_ _07647_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07170__B1 _07169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07577_ _07577_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07579_/B sky130_fd_sc_hd__xnor2_1
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05720__A1 _08082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09316_ _09316_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09388_/A sky130_fd_sc_hd__xor2_2
X_06528_ _06785_/A _06540_/A vssd1 vssd1 vccd1 vccd1 _06528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_166_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09247_ hold4/A _09243_/X _09244_/X _09246_/X _09239_/X vssd1 vssd1 vccd1 vccd1 _09248_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_167_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06459_ _10977_/Q _06459_/B vssd1 vssd1 vccd1 vccd1 _06670_/A sky130_fd_sc_hd__nand2_1
XFILLER_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09178_ _09113_/A _09177_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09178_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08490__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _08132_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08129_/X sky130_fd_sc_hd__or2_1
XFILLER_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10244__B _10937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput56 _10834_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[0] sky130_fd_sc_hd__buf_2
XFILLER_122_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput67 _10835_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[1] sky130_fd_sc_hd__buf_2
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput78 _10836_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[2] sky130_fd_sc_hd__buf_2
XFILLER_150_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10022_ _10022_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _10029_/A sky130_fd_sc_hd__nand2_1
XFILLER_76_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10532__A1 _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input16_A io_wbs_m2s_data[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09150__A1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10924_ _10930_/CLK _10924_/D vssd1 vssd1 vccd1 vccd1 _10924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _10855_/CLK _10855_/D vssd1 vssd1 vccd1 vccd1 _10855_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10786_ _10788_/CLK _10786_/D vssd1 vssd1 vccd1 vccd1 _10786_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08110__C1 _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05830_ _05830_/A vssd1 vssd1 vccd1 vccd1 _08027_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10170__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05761_ _05749_/A _10564_/Q _10563_/Q _08282_/A vssd1 vssd1 vccd1 vccd1 _05761_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_82_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05950__A1 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07500_ _07504_/B _07535_/A _07504_/A vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__o21ai_2
X_08480_ _08483_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08481_/A sky130_fd_sc_hd__and2_1
X_05692_ _05692_/A vssd1 vssd1 vccd1 vccd1 _05693_/A sky130_fd_sc_hd__inv_2
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07431_ _07562_/A vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07362_ _07363_/B _07363_/C _07361_/Y vssd1 vssd1 vccd1 vccd1 _07410_/A sky130_fd_sc_hd__a21bo_1
XFILLER_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09101_ _10938_/Q _10369_/B _09100_/Y _08968_/A vssd1 vssd1 vccd1 vccd1 _09101_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06313_ _06313_/A _06313_/B vssd1 vssd1 vccd1 vccd1 _06755_/A sky130_fd_sc_hd__nand2_2
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07293_ _07317_/A vssd1 vssd1 vccd1 vccd1 _07309_/C sky130_fd_sc_hd__inv_2
X_09032_ _10504_/A _09031_/X _09087_/S vssd1 vssd1 vccd1 vccd1 _09032_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06244_ _10611_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06244_/X sky130_fd_sc_hd__or2_1
XFILLER_148_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06175_ _06175_/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10211__B1 _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09934_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _10009_/A sky130_fd_sc_hd__or2_1
XFILLER_86_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input8_A io_wbs_m2s_addr[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09865_ _09867_/D vssd1 vssd1 vccd1 vccd1 _10139_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_100_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10514__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _10816_/Q _08856_/B vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__xor2_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _09372_/C _09733_/B _09372_/B vssd1 vssd1 vccd1 vccd1 _09797_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06194__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08747_ _08759_/A _08747_/B _08778_/A vssd1 vssd1 vccd1 vccd1 _08747_/X sky130_fd_sc_hd__and3b_1
XFILLER_27_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05959_ input50/X input48/X vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__and2_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08678_/A vssd1 vssd1 vccd1 vccd1 _08698_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08485__A _09090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05902__A _08119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07629_ _07662_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07630_/B sky130_fd_sc_hd__nor2_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10640_ _10640_/CLK _10640_/D vssd1 vssd1 vccd1 vccd1 _10640_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06436__C _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _10855_/CLK _10571_/D vssd1 vssd1 vccd1 vccd1 _10571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07829__A _07850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09199__A1 _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10505__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10005_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05932__B2 _08233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10907_ _10929_/CLK _10907_/D vssd1 vssd1 vccd1 vccd1 _10907_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10838_ _10856_/CLK _10838_/D vssd1 vssd1 vccd1 vccd1 _10838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07437__A1 _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10769_ _10833_/CLK _10769_/D vssd1 vssd1 vccd1 vccd1 _10769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07980_ _06182_/X _07965_/X _07979_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10658_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06931_ _06936_/A _06936_/B _06930_/Y vssd1 vssd1 vccd1 vccd1 _06935_/B sky130_fd_sc_hd__a21o_2
XFILLER_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09650_ _09620_/A _09648_/X _09649_/X vssd1 vssd1 vccd1 vccd1 _09779_/A sky130_fd_sc_hd__a21o_1
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06862_ _06862_/A _06862_/B vssd1 vssd1 vccd1 vccd1 _06863_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_83_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08601_ _10783_/Q _08600_/X _10784_/Q vssd1 vssd1 vccd1 vccd1 _08602_/C sky130_fd_sc_hd__a21o_1
XFILLER_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05813_ _05813_/A _10574_/Q vssd1 vssd1 vccd1 vccd1 _05813_/X sky130_fd_sc_hd__xor2_1
X_09581_ _09638_/C _09703_/A vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__nor2_1
XFILLER_94_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06793_ _06833_/A _06793_/B vssd1 vssd1 vccd1 vccd1 _06794_/B sky130_fd_sc_hd__and2_1
XANTENNA__05923__A1 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08532_ _08531_/X _08547_/A _10767_/Q vssd1 vssd1 vccd1 vccd1 _08533_/B sky130_fd_sc_hd__mux2_1
XFILLER_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05744_ _08218_/A vssd1 vssd1 vccd1 vccd1 _05744_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10985__D _10985_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08463_ _10775_/Q _10738_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08464_/B sky130_fd_sc_hd__mux2_1
X_05675_ _08277_/B _05596_/X _05593_/X _08277_/A _05674_/X vssd1 vssd1 vccd1 vccd1
+ _05675_/X sky130_fd_sc_hd__o221a_1
XFILLER_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ _07414_/A _07051_/A vssd1 vssd1 vccd1 vccd1 _07430_/A sky130_fd_sc_hd__or2b_1
X_08394_ _08394_/A vssd1 vssd1 vccd1 vccd1 _08394_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07345_ _07345_/A _07345_/B vssd1 vssd1 vccd1 vccd1 _07488_/A sky130_fd_sc_hd__xor2_1
XFILLER_148_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_137_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07276_ _07318_/B _07324_/A _07318_/A vssd1 vssd1 vccd1 vccd1 _07319_/A sky130_fd_sc_hd__a21oi_2
XFILLER_148_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _10502_/A _09012_/X _09087_/S vssd1 vssd1 vccd1 vccd1 _09015_/X sky130_fd_sc_hd__mux2_1
X_06227_ _10604_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06227_/X sky130_fd_sc_hd__or2_1
XFILLER_117_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09305__A_N _10898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06158_ _06204_/B vssd1 vssd1 vccd1 vccd1 _06158_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06089_ _06089_/A _06089_/B _06089_/C _06089_/D vssd1 vssd1 vccd1 vccd1 _06089_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_77_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09917_ _09855_/A _09855_/B _09852_/A vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__a21o_1
XFILLER_104_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09848_ _09848_/A _09848_/B _09848_/C vssd1 vssd1 vccd1 vccd1 _09901_/B sky130_fd_sc_hd__and3_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08561__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09787_/A sky130_fd_sc_hd__nand2_1
XFILLER_85_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09104__A _09104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07419__A1 _07416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10623_ _10653_/CLK _10623_/D vssd1 vssd1 vccd1 vccd1 _10623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10554_ _10554_/CLK _10554_/D vssd1 vssd1 vccd1 vccd1 _10554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10485_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10485_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_2_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_78_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05460_ _07871_/A _05460_/B _05460_/C _05460_/D vssd1 vssd1 vccd1 vccd1 _05460_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05391_ _06038_/A _05391_/B vssd1 vssd1 vccd1 vccd1 _05392_/B sky130_fd_sc_hd__and2_1
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07130_ _07134_/A _07133_/A _07133_/B _07123_/B _07144_/A vssd1 vssd1 vccd1 vccd1
+ _07132_/A sky130_fd_sc_hd__o32ai_4
XFILLER_119_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07061_ _07061_/A _07061_/B vssd1 vssd1 vccd1 vccd1 _07164_/B sky130_fd_sc_hd__xnor2_4
XFILLER_146_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06012_ _06011_/X _05993_/S _05977_/X vssd1 vssd1 vccd1 vccd1 _06012_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09032__A0 _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09583__A1 _10969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07963_ _07963_/A vssd1 vssd1 vccd1 vccd1 _10655_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09702_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__xor2_1
X_06914_ _06914_/A _06914_/B vssd1 vssd1 vccd1 vccd1 _06939_/A sky130_fd_sc_hd__xnor2_4
XFILLER_56_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07894_ _10605_/Q _07888_/X _07892_/X _07893_/Y vssd1 vssd1 vccd1 vccd1 _07895_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09633_ _09631_/A _09631_/B _09631_/C vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__o21a_1
XFILLER_83_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06845_ _06845_/A _07784_/B _06845_/C vssd1 vssd1 vccd1 vccd1 _06847_/A sky130_fd_sc_hd__and3_1
XFILLER_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09566_/A sky130_fd_sc_hd__xor2_1
X_06776_ _06776_/A vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08515_ _08638_/B _08514_/X _08509_/X _10757_/Q vssd1 vssd1 vccd1 vccd1 _10757_/D
+ sky130_fd_sc_hd__a22o_1
X_05727_ _08130_/A _05739_/B _05549_/A _08117_/A vssd1 vssd1 vccd1 vccd1 _05732_/C
+ sky130_fd_sc_hd__a22o_1
X_09495_ _09610_/A _09492_/A _09494_/D _09494_/B vssd1 vssd1 vccd1 vccd1 _09496_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_169_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08446_ _10770_/Q _10733_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08447_/B sky130_fd_sc_hd__mux2_1
X_05658_ _05631_/X _05657_/X _05628_/X _05896_/A vssd1 vssd1 vccd1 vccd1 _05658_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08377_ _08367_/X _10732_/Q _07865_/X _08376_/X vssd1 vssd1 vccd1 vccd1 _10714_/D
+ sky130_fd_sc_hd__o211a_1
X_05589_ _10703_/Q vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07328_ _07326_/A _07394_/A _07327_/X _07086_/B vssd1 vssd1 vccd1 vccd1 _07328_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07259_ _07197_/A _07076_/B _07197_/C vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__a21oi_1
XFILLER_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10270_ _10287_/B _10268_/A _10279_/S vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10533__A _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08003__A _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08301__A2 _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08673__A _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_63_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10914_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10606_ _10822_/CLK _10606_/D vssd1 vssd1 vccd1 vccd1 _10606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06076__B1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10537_ _10537_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10537_/X sky130_fd_sc_hd__or3_1
XFILLER_128_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_78_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10881_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10468_ _06195_/X _10459_/X _10467_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10960_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10399_ _10399_/A vssd1 vssd1 vccd1 vccd1 _10399_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_69_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06630_ _06630_/A _06630_/B vssd1 vssd1 vccd1 vccd1 _06631_/B sky130_fd_sc_hd__or2_1
XFILLER_53_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06561_ _06587_/B _06561_/B _06561_/C vssd1 vssd1 vccd1 vccd1 _06573_/C sky130_fd_sc_hd__and3b_1
XFILLER_33_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08300_ _08263_/X _08315_/C _08296_/Y _08299_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08300_/X sky130_fd_sc_hd__o311a_1
X_05512_ _05348_/X _05510_/X _05506_/X _07893_/A vssd1 vssd1 vccd1 vccd1 _10562_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09280_ _09280_/A vssd1 vssd1 vccd1 vccd1 _10861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06492_ _06567_/A _06515_/B vssd1 vssd1 vccd1 vccd1 _06493_/C sky130_fd_sc_hd__nand2_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08231_ _08227_/X _08229_/X _08230_/X vssd1 vssd1 vccd1 vccd1 _10697_/D sky130_fd_sc_hd__o21a_1
X_05443_ _10642_/Q _05438_/X _05442_/Y vssd1 vssd1 vccd1 vccd1 _05443_/X sky130_fd_sc_hd__o21ba_1
XFILLER_60_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08162_ _08158_/X _08169_/C _08067_/X vssd1 vssd1 vccd1 vccd1 _08162_/Y sky130_fd_sc_hd__o21ai_1
X_05374_ _05374_/A _05374_/B vssd1 vssd1 vccd1 vccd1 _05374_/X sky130_fd_sc_hd__and2_1
XFILLER_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07113_ _07113_/A _07113_/B vssd1 vssd1 vccd1 vccd1 _07216_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06067__B1 _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08093_ _08093_/A vssd1 vssd1 vccd1 vccd1 _08098_/A sky130_fd_sc_hd__buf_2
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07927__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ _07044_/A vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05290__A1 _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08995_ _08995_/A vssd1 vssd1 vccd1 vccd1 _08995_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_07946_ _07946_/A vssd1 vssd1 vccd1 vccd1 _10650_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07877_ _07880_/A _07877_/B vssd1 vssd1 vccd1 vccd1 _10632_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09616_ _09652_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09619_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06828_ _06828_/A _06828_/B vssd1 vssd1 vccd1 vccd1 _06882_/B sky130_fd_sc_hd__nand2_1
XFILLER_141_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09547_ _09676_/A _09547_/B vssd1 vssd1 vccd1 vccd1 _09549_/A sky130_fd_sc_hd__xnor2_4
X_06759_ _06759_/A _06759_/B vssd1 vssd1 vccd1 vccd1 _06779_/B sky130_fd_sc_hd__nor2_1
XFILLER_93_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09478_ _09438_/A _09438_/B _09477_/X vssd1 vssd1 vccd1 vccd1 _09479_/B sky130_fd_sc_hd__a21oi_1
XFILLER_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08429_ _10772_/Q _10771_/Q _08547_/B vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__and3_1
XANTENNA__10528__A _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10322_ _10961_/Q _10945_/Q vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__and2b_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10253_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10253_/Y sky130_fd_sc_hd__nand2_1
XFILLER_121_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10184_ _10355_/A vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__buf_2
XFILLER_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input46_A io_wbs_m2s_data[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07572__A _09379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05820__A _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07747__A _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07800_ _06934_/A _06934_/B _07799_/Y vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__a21oi_1
X_08780_ _08992_/A vssd1 vssd1 vccd1 vccd1 _08780_/X sky130_fd_sc_hd__clkbuf_4
X_05992_ input45/X _05992_/B vssd1 vssd1 vccd1 vccd1 _05992_/X sky130_fd_sc_hd__xor2_1
XFILLER_111_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07731_ _07731_/A _07731_/B vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07662_ _07662_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07663_/B sky130_fd_sc_hd__nor2_1
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09401_ _09437_/A _09401_/B vssd1 vssd1 vccd1 vccd1 _09402_/C sky130_fd_sc_hd__or2_1
X_06613_ _06614_/A _06614_/B _06614_/C vssd1 vssd1 vccd1 vccd1 _06674_/C sky130_fd_sc_hd__a21o_1
XFILLER_81_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07593_ _07593_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _07596_/A sky130_fd_sc_hd__xnor2_2
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09332_ _10900_/Q _10884_/Q vssd1 vssd1 vccd1 vccd1 _09333_/B sky130_fd_sc_hd__and2b_1
X_06544_ _06544_/A _06544_/B vssd1 vssd1 vccd1 vccd1 _06622_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09263_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09287_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06475_ _06666_/B _06671_/A _06666_/A vssd1 vssd1 vccd1 vccd1 _06688_/B sky130_fd_sc_hd__a21bo_1
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08214_ _08211_/X _08214_/B vssd1 vssd1 vccd1 vccd1 _08215_/A sky130_fd_sc_hd__and2b_1
X_05426_ _07871_/A _05363_/X _05360_/X _10632_/Q _05425_/X vssd1 vssd1 vccd1 vccd1
+ _05426_/X sky130_fd_sc_hd__o221a_1
X_09194_ _10962_/Q _09194_/B vssd1 vssd1 vccd1 vccd1 _09194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ _08145_/A vssd1 vssd1 vccd1 vccd1 _10688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05357_ _06052_/A _05848_/B _10665_/Q vssd1 vssd1 vccd1 vccd1 _05358_/B sky130_fd_sc_hd__o21ai_1
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08076_ _08038_/X _08074_/X _08075_/Y _08044_/X _06065_/X vssd1 vssd1 vccd1 vccd1
+ _08076_/X sky130_fd_sc_hd__a32o_1
X_05288_ _06065_/A _05283_/Y _05287_/Y vssd1 vssd1 vccd1 vccd1 _05400_/A sky130_fd_sc_hd__a21o_1
XFILLER_136_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07027_ _09344_/B _07007_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _07028_/B sky130_fd_sc_hd__o21ai_1
XFILLER_115_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08978_ _08978_/A vssd1 vssd1 vccd1 vccd1 _09020_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__05905__A _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07929_ _08284_/A _07929_/B vssd1 vssd1 vccd1 vccd1 _10647_/D sky130_fd_sc_hd__nor2_1
XFILLER_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _10940_/CLK _10940_/D vssd1 vssd1 vccd1 vccd1 _10940_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _10970_/CLK _10871_/D vssd1 vssd1 vccd1 vccd1 _10871_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10305_ _10943_/Q _10959_/Q vssd1 vssd1 vccd1 vccd1 _10307_/A sky130_fd_sc_hd__and2b_1
XFILLER_113_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10236_ _10225_/A _10246_/B _10225_/B vssd1 vssd1 vccd1 vccd1 _10236_/X sky130_fd_sc_hd__o21ba_1
XFILLER_106_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10167_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10167_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07951__A0 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08398__A _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10098_ _10098_/A _10098_/B vssd1 vssd1 vccd1 vccd1 _10100_/C sky130_fd_sc_hd__or2_1
XFILLER_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06047__A1_N _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08259__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06260_ _10919_/Q _10902_/Q vssd1 vssd1 vccd1 vccd1 _06262_/A sky130_fd_sc_hd__nand2_1
XFILLER_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06191_ input19/X vssd1 vssd1 vccd1 vccd1 _06191_/X sky130_fd_sc_hd__buf_4
XFILLER_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09950_ _09744_/A _09949_/A _09830_/X vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__o21a_1
XFILLER_144_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08901_ _09154_/A vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__buf_4
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09811_/B _09452_/A _09452_/B _10097_/A vssd1 vssd1 vccd1 vccd1 _09882_/B
+ sky130_fd_sc_hd__a31o_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08832_ input25/X _08830_/X _08831_/X hold3/A vssd1 vssd1 vccd1 vccd1 _08832_/X sky130_fd_sc_hd__a22o_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05975_ _05993_/S vssd1 vssd1 vccd1 vccd1 _05975_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08763_ _06182_/X _08728_/X _08729_/X _10809_/Q vssd1 vssd1 vccd1 vccd1 _08763_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07714_ _07713_/B _07713_/Y _07714_/S vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _08819_/A vssd1 vssd1 vccd1 vccd1 _08694_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07940__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07645_ _07645_/A _07645_/B vssd1 vssd1 vccd1 vccd1 _07647_/B sky130_fd_sc_hd__xnor2_4
XFILLER_81_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07576_ _07576_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06556__A _10971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09315_ _10899_/Q _10883_/Q vssd1 vssd1 vccd1 vccd1 _09337_/B sky130_fd_sc_hd__xor2_4
X_06527_ _06527_/A vssd1 vssd1 vccd1 vccd1 _06785_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ _05851_/A _09245_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09246_/X sky130_fd_sc_hd__mux2_1
X_06458_ _06458_/A _06458_/B vssd1 vssd1 vccd1 vccd1 _06646_/A sky130_fd_sc_hd__xnor2_1
XFILLER_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05484__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05409_ _10617_/Q vssd1 vssd1 vccd1 vccd1 _08994_/A sky130_fd_sc_hd__clkbuf_2
X_09177_ _09114_/A _09176_/X _10500_/B vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__o21a_1
X_06389_ _06412_/A _06389_/B vssd1 vssd1 vccd1 vccd1 _06502_/C sky130_fd_sc_hd__xnor2_2
XFILLER_135_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08128_ _08128_/A vssd1 vssd1 vccd1 vccd1 _10686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08059_ _08059_/A _08082_/D vssd1 vssd1 vccd1 vccd1 _08072_/B sky130_fd_sc_hd__nand2_1
XFILLER_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput57 _10844_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[10] sky130_fd_sc_hd__buf_2
Xoutput68 _10854_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[20] sky130_fd_sc_hd__buf_2
XFILLER_89_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput79 _10864_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[30] sky130_fd_sc_hd__buf_2
X_10021_ _10021_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__or2_1
XFILLER_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09107__A _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08011__A _08268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07850__A _07850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10923_ _10930_/CLK _10923_/D vssd1 vssd1 vccd1 vccd1 _10923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10854_ _10857_/CLK _10854_/D vssd1 vssd1 vccd1 vccd1 _10854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10785_ _10788_/CLK _10785_/D vssd1 vssd1 vccd1 vccd1 _10785_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10219_ _10216_/X _10217_/X _10329_/S vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__mux2_1
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05760_ _08232_/A _10559_/Q _10558_/Q _08228_/A vssd1 vssd1 vccd1 vccd1 _05764_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_36_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05691_ _08169_/A vssd1 vssd1 vccd1 vccd1 _05692_/A sky130_fd_sc_hd__buf_2
XFILLER_63_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ _07430_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__xnor2_2
X_07361_ _07406_/A _07361_/B vssd1 vssd1 vccd1 vccd1 _07361_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_50_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06312_ _10926_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _06313_/B sky130_fd_sc_hd__or2_1
X_09100_ _10954_/Q _09124_/A vssd1 vssd1 vccd1 vccd1 _09100_/Y sky130_fd_sc_hd__nor2_1
X_07292_ _07326_/A _07076_/B _07390_/B _07563_/A vssd1 vssd1 vccd1 vccd1 _07298_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08591__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09031_ _10482_/A _09030_/X _09086_/S vssd1 vssd1 vccd1 vccd1 _09031_/X sky130_fd_sc_hd__mux2_1
X_06243_ input34/X _06238_/X _06242_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10610_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06174_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06193_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07000__A _09920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10211__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09933_ _09933_/A _09933_/B vssd1 vssd1 vccd1 vccd1 _09935_/B sky130_fd_sc_hd__xor2_1
XFILLER_132_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _09864_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09867_/D sky130_fd_sc_hd__xnor2_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08815_ hold13/X _08815_/B vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__nand2_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09795_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09883_/A sky130_fd_sc_hd__xor2_4
XFILLER_86_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08746_ _08743_/Y _08744_/X _08740_/X _08741_/X vssd1 vssd1 vccd1 vccd1 _08747_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05958_ _10531_/A vssd1 vssd1 vccd1 vccd1 _05958_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07670__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08670_/X _08675_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10800_/D sky130_fd_sc_hd__o21a_1
XANTENNA__07143__A1 _10985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05889_ _10659_/Q _05891_/A _05886_/B _05886_/A vssd1 vssd1 vccd1 vccd1 _05889_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08340__B1 _05570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07628_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _07698_/A sky130_fd_sc_hd__xor2_4
XFILLER_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07559_ _07724_/A _07559_/B vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__or2_1
X_10570_ _10855_/CLK _10570_/D vssd1 vssd1 vccd1 vccd1 _10570_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _09229_/A vssd1 vssd1 vccd1 vccd1 _10853_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09199__A2 _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08006__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10271__A _10287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10004_ _09940_/B _10078_/A _10003_/X vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__o21a_1
XFILLER_67_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08676__A _08992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10906_ _10925_/CLK _10906_/D vssd1 vssd1 vccd1 vccd1 _10906_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05696__B2 _08160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10837_ _10848_/CLK _10837_/D vssd1 vssd1 vccd1 vccd1 _10837_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10768_ _10770_/CLK _10768_/D vssd1 vssd1 vccd1 vccd1 _10768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10699_ _10704_/CLK _10699_/D vssd1 vssd1 vccd1 vccd1 _10699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06930_ _06930_/A _06930_/B vssd1 vssd1 vccd1 vccd1 _06930_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10181__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06861_ _06862_/A _06862_/B vssd1 vssd1 vccd1 vccd1 _06863_/A sky130_fd_sc_hd__and2_1
XFILLER_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08600_ _08600_/A vssd1 vssd1 vccd1 vccd1 _08600_/X sky130_fd_sc_hd__clkbuf_2
X_05812_ _10649_/Q vssd1 vssd1 vccd1 vccd1 _05813_/A sky130_fd_sc_hd__buf_4
X_09580_ _10970_/Q _09744_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__nand2_1
X_06792_ _06792_/A _06792_/B vssd1 vssd1 vccd1 vccd1 _06793_/B sky130_fd_sc_hd__or2_1
XFILLER_83_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08531_ _08531_/A _08661_/A vssd1 vssd1 vccd1 vccd1 _08531_/X sky130_fd_sc_hd__or2_1
X_05743_ _08224_/B vssd1 vssd1 vccd1 vccd1 _08218_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08322__B1 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05674_ _05598_/X _05599_/X _05596_/X _10701_/Q _05673_/X vssd1 vssd1 vccd1 vccd1
+ _05674_/X sky130_fd_sc_hd__a221o_1
XFILLER_24_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08462_ _08462_/A vssd1 vssd1 vccd1 vccd1 _08477_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ _07549_/A _07413_/B vssd1 vssd1 vccd1 vccd1 _07598_/A sky130_fd_sc_hd__and2_1
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08393_ _08383_/X _10738_/Q _08380_/X _08392_/X vssd1 vssd1 vccd1 vccd1 _10720_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_11_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07344_ _07344_/A _07344_/B vssd1 vssd1 vccd1 vccd1 _07345_/A sky130_fd_sc_hd__and2_1
XFILLER_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09210__A _09274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07275_ _07275_/A _07275_/B vssd1 vssd1 vccd1 vccd1 _07318_/A sky130_fd_sc_hd__xnor2_1
XFILLER_164_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06226_ _06253_/B vssd1 vssd1 vccd1 vccd1 _06236_/B sky130_fd_sc_hd__clkbuf_1
X_09014_ _09016_/A _10341_/C vssd1 vssd1 vccd1 vccd1 _09087_/S sky130_fd_sc_hd__or2_2
XFILLER_117_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06157_ _05958_/X _06131_/X _06156_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10588_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09050__A1 _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09050__B2 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06088_ _05778_/Y _10679_/Q _07985_/A _08180_/A _06087_/X vssd1 vssd1 vccd1 vccd1
+ _06089_/D sky130_fd_sc_hd__a221o_1
XFILLER_160_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09916_ _09916_/A _09916_/B vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09847_ _09716_/Y _09780_/X _09781_/Y _09718_/Y vssd1 vssd1 vccd1 vccd1 _09848_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09851_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _09827_/A sky130_fd_sc_hd__nor2_2
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _08831_/A vssd1 vssd1 vccd1 vccd1 _08729_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10622_ _10653_/CLK _10622_/D vssd1 vssd1 vccd1 vccd1 _10622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10553_ _10554_/CLK _10553_/D vssd1 vssd1 vccd1 vccd1 _10553_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10266__A _10938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10484_ _10484_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10484_/X sky130_fd_sc_hd__or2_1
XFILLER_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09041__A1 _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10187__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05390_ _10653_/Q vssd1 vssd1 vccd1 vccd1 _06038_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07060_ _07112_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07061_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06011_ _06011_/A vssd1 vssd1 vccd1 vccd1 _06011_/X sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_44_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07962_ _08443_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _07963_/A sky130_fd_sc_hd__or2_1
XFILLER_99_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09701_ _09844_/A _09701_/B vssd1 vssd1 vccd1 vccd1 _09773_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06913_ _06913_/A _06923_/B vssd1 vssd1 vccd1 vccd1 _06914_/B sky130_fd_sc_hd__xnor2_2
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07893_ _07893_/A vssd1 vssd1 vccd1 vccd1 _07893_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09632_ _09757_/A vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06844_ _10510_/A _07783_/B _06844_/C vssd1 vssd1 vccd1 vccd1 _06845_/C sky130_fd_sc_hd__and3_1
XFILLER_83_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05733__A _08082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09563_ _09563_/A _09563_/B vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06775_ _06775_/A _06776_/A _06775_/C vssd1 vssd1 vccd1 vccd1 _06792_/A sky130_fd_sc_hd__and3_1
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08514_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08514_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05726_ _05726_/A vssd1 vssd1 vccd1 vccd1 _08117_/A sky130_fd_sc_hd__buf_2
X_09494_ _09610_/A _09494_/B _09696_/A _09494_/D vssd1 vssd1 vccd1 vccd1 _09542_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_63_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08445_ _08445_/A vssd1 vssd1 vccd1 vccd1 _08460_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05657_ _10687_/Q _05631_/B _05632_/Y _05726_/A _05656_/X vssd1 vssd1 vccd1 vccd1
+ _05657_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05588_ _05588_/A _05588_/B vssd1 vssd1 vccd1 vccd1 _05588_/X sky130_fd_sc_hd__and2_1
X_08376_ _08381_/A _10748_/Q vssd1 vssd1 vccd1 vccd1 _08376_/X sky130_fd_sc_hd__or2_1
XFILLER_149_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07327_ _07327_/A vssd1 vssd1 vccd1 vccd1 _07327_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_109_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07258_ _07258_/A _07258_/B vssd1 vssd1 vccd1 vccd1 _07273_/A sky130_fd_sc_hd__xor2_1
XFILLER_165_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05832__A1 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06209_ input9/X _10432_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09104_/B sky130_fd_sc_hd__nand3_1
X_07189_ _07197_/A _07587_/B _07188_/C vssd1 vssd1 vccd1 vccd1 _07190_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10169__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05899__A1 _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10605_ _10822_/CLK _10605_/D vssd1 vssd1 vccd1 vccd1 _10605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _07729_/A _10522_/A _10535_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10985_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10467_ _10960_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10467_/X sky130_fd_sc_hd__or2_1
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05818__A _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__C1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10398_ _10938_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10398_/X sky130_fd_sc_hd__and2_1
XFILLER_69_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06560_ _06587_/A _06587_/B _06587_/C _07676_/A vssd1 vssd1 vccd1 vccd1 _06585_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08864__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05511_ _05346_/X _05510_/X _05506_/X _07889_/A vssd1 vssd1 vccd1 vccd1 _10561_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_06491_ _06568_/A vssd1 vssd1 vccd1 vccd1 _06527_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05442_ _05834_/A _05442_/B vssd1 vssd1 vccd1 vccd1 _05442_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08230_ input24/X _08164_/X _08165_/X _06061_/A _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08230_/X sky130_fd_sc_hd__o221a_1
XFILLER_166_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ _07979_/A _08306_/B _08159_/X _08173_/B _06011_/X vssd1 vssd1 vccd1 vccd1
+ _08161_/X sky130_fd_sc_hd__o221a_1
X_05373_ _10659_/Q _05373_/B vssd1 vssd1 vccd1 vccd1 _05374_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07112_ _07112_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07113_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06067__B2 _08082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08092_ _08092_/A vssd1 vssd1 vccd1 vccd1 _08092_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07043_ _07043_/A _07043_/B vssd1 vssd1 vccd1 vccd1 _07048_/B sky130_fd_sc_hd__nor2_1
XANTENNA__05814__A1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08104__A _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08994_ _08994_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _08994_/X sky130_fd_sc_hd__or2_1
XFILLER_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07945_ _07955_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07946_/A sky130_fd_sc_hd__or2_1
XFILLER_56_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07876_ hold7/X _07870_/X _07874_/X _07875_/Y vssd1 vssd1 vccd1 vccd1 _07877_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_141_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09615_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__xor2_1
X_06827_ _06844_/C _06856_/C vssd1 vssd1 vccd1 vccd1 _06883_/A sky130_fd_sc_hd__xor2_1
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09546_ _09546_/A _09546_/B vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__nand2_2
XFILLER_70_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06758_ _06758_/A _06758_/B _06758_/C _06786_/A vssd1 vssd1 vccd1 vccd1 _06759_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_24_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05709_ _08169_/B vssd1 vssd1 vccd1 vccd1 _05709_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09477_ _09436_/A _09477_/B vssd1 vssd1 vccd1 vccd1 _09477_/X sky130_fd_sc_hd__and2b_1
XFILLER_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06689_ _06690_/A _06690_/B vssd1 vssd1 vccd1 vccd1 _06691_/A sky130_fd_sc_hd__nand2_1
XFILLER_52_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08428_ _10770_/Q _10769_/Q _10768_/Q _10767_/Q vssd1 vssd1 vccd1 vccd1 _08547_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_24_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05502__B1 _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08359_ _05528_/A _08349_/X _08358_/Y vssd1 vssd1 vccd1 vccd1 _08359_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10321_ _07570_/A _10283_/X _10320_/X _10293_/X vssd1 vssd1 vccd1 vccd1 _10911_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10252_ _10252_/A _10252_/B vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__xnor2_1
XFILLER_133_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10183_ _07028_/A _10181_/X _10177_/X _10893_/Q vssd1 vssd1 vccd1 vccd1 _10893_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08949__A input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06230__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07853__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A io_wbs_m2s_data[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10519_ _10537_/B vssd1 vssd1 vccd1 vccd1 _10531_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05991_ _07899_/A vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__buf_2
X_07730_ _07730_/A _07730_/B vssd1 vssd1 vccd1 vccd1 _07731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07661_ _07661_/A _07661_/B vssd1 vssd1 vccd1 vccd1 _07665_/A sky130_fd_sc_hd__xnor2_1
XFILLER_65_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09400_ _09399_/B _09400_/B vssd1 vssd1 vccd1 vccd1 _09401_/B sky130_fd_sc_hd__and2b_1
XFILLER_65_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06612_ _06612_/A _06612_/B vssd1 vssd1 vccd1 vccd1 _06614_/C sky130_fd_sc_hd__nor2_1
XFILLER_92_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07592_ _07592_/A _07592_/B vssd1 vssd1 vccd1 vccd1 _07593_/B sky130_fd_sc_hd__nand2_1
XFILLER_34_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _10884_/Q _10900_/Q vssd1 vssd1 vccd1 vccd1 _09333_/A sky130_fd_sc_hd__and2b_1
X_06543_ _06544_/B _06544_/A vssd1 vssd1 vccd1 vccd1 _06624_/A sky130_fd_sc_hd__or2b_1
XFILLER_52_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _08304_/A _07907_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09262_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06474_ _06474_/A _06474_/B vssd1 vssd1 vccd1 vccd1 _06666_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08213_ input22/X _08212_/X _08124_/X _08208_/A _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08214_/B sky130_fd_sc_hd__o221a_1
X_05425_ _05460_/B _05366_/Y _05363_/X _10631_/Q _05424_/X vssd1 vssd1 vccd1 vccd1
+ _05425_/X sky130_fd_sc_hd__a221o_1
X_09193_ _09202_/A _09193_/B vssd1 vssd1 vccd1 vccd1 _10848_/D sky130_fd_sc_hd__nor2_2
XFILLER_119_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07938__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__and2_1
X_05356_ _05363_/A vssd1 vssd1 vccd1 vccd1 _05848_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_146_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05287_ _05401_/A _05406_/A vssd1 vssd1 vccd1 vccd1 _05287_/Y sky130_fd_sc_hd__nor2_1
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08075_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_135_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07026_ _07509_/A _07421_/A _07025_/Y vssd1 vssd1 vccd1 vccd1 _07042_/A sky130_fd_sc_hd__a21oi_1
XFILLER_150_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08977_ _09124_/A _09124_/B _09124_/C vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__or3_1
XFILLER_29_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_62_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10653_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07928_ _10615_/Q _07906_/A _05525_/A _07874_/A vssd1 vssd1 vccd1 vccd1 _07929_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_57_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07859_ _10878_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10870_ _10879_/CLK _10870_/D vssd1 vssd1 vccd1 vccd1 _10870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_77_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10879_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _09568_/A _09529_/B vssd1 vssd1 vccd1 vccd1 _09529_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07848__A _07848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10304_ _07028_/A _10283_/X _10303_/Y _10293_/X vssd1 vssd1 vccd1 vccd1 _10909_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10235_ _10233_/X _10235_/B vssd1 vssd1 vccd1 vccd1 _10246_/C sky130_fd_sc_hd__and2b_1
XFILLER_106_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10166_ _10881_/Q _10115_/X _10165_/Y _10043_/X vssd1 vssd1 vccd1 vccd1 _10881_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07951__A1 _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06199__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10097_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/B sky130_fd_sc_hd__and2_1
XFILLER_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06190_ _06187_/X _06183_/X _06189_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10595_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10184__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ _08897_/Y _08898_/X _08899_/X vssd1 vssd1 vccd1 vccd1 _10826_/D sky130_fd_sc_hd__o21a_1
XFILLER_171_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09880_/A vssd1 vssd1 vccd1 vccd1 _10097_/A sky130_fd_sc_hd__buf_2
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08831_ _08831_/A vssd1 vssd1 vccd1 vccd1 _08831_/X sky130_fd_sc_hd__clkbuf_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08804_/A _08804_/B _08760_/X _08761_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08762_/X sky130_fd_sc_hd__o311a_1
X_05974_ _06120_/S vssd1 vssd1 vccd1 vccd1 _05993_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_100_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07713_ _07713_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07713_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08693_ _08693_/A _08693_/B vssd1 vssd1 vccd1 vccd1 _08693_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07644_ _07662_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07645_/B sky130_fd_sc_hd__or2_2
XFILLER_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07170__A2 _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09213__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07575_ _07574_/A _07574_/B _07574_/C vssd1 vssd1 vccd1 vccd1 _07576_/B sky130_fd_sc_hd__a21oi_1
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09314_ _09314_/A _09314_/B vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__nor2_2
X_06526_ _06541_/C _06512_/B _06511_/A vssd1 vssd1 vccd1 vccd1 _06535_/B sky130_fd_sc_hd__o21a_1
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09245_ _08278_/A _07896_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09245_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06457_ _06457_/A _06465_/A vssd1 vssd1 vccd1 vccd1 _06458_/B sky130_fd_sc_hd__nor2_1
X_05408_ _10648_/Q vssd1 vssd1 vccd1 vccd1 _05408_/Y sky130_fd_sc_hd__clkinv_4
X_09176_ _10944_/Q _09143_/Y _09175_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09176_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06388_ _06388_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06389_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08127_ _08122_/X _08127_/B vssd1 vssd1 vccd1 vccd1 _08128_/A sky130_fd_sc_hd__and2b_1
X_05339_ _10670_/Q _05854_/A _10671_/Q vssd1 vssd1 vccd1 vccd1 _05340_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10094__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08058_ _08058_/A vssd1 vssd1 vccd1 vccd1 _08058_/X sky130_fd_sc_hd__buf_2
XFILLER_123_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07009_ _07030_/C vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xoutput58 _10845_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[11] sky130_fd_sc_hd__buf_2
Xoutput69 _10855_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[21] sky130_fd_sc_hd__buf_2
XFILLER_131_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10020_ _10021_/A _10021_/B vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08011__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10922_ _10930_/CLK _10922_/D vssd1 vssd1 vccd1 vccd1 _10922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09123__A _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10853_ _10853_/CLK _10853_/D vssd1 vssd1 vccd1 vccd1 _10853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10784_ _10784_/CLK _10784_/D vssd1 vssd1 vccd1 vccd1 _10784_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08110__A1 _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08110__B2 _05728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10218_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10329_/S sky130_fd_sc_hd__buf_2
XFILLER_121_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10149_ _10023_/A _10023_/B _10095_/A _10098_/A vssd1 vssd1 vccd1 vccd1 _10151_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_121_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05690_ _05528_/X _05564_/Y _05689_/X vssd1 vssd1 vccd1 vccd1 _10728_/D sky130_fd_sc_hd__o21ai_1
XANTENNA__08885__C1 _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07360_ _07360_/A _07407_/A vssd1 vssd1 vccd1 vccd1 _07361_/B sky130_fd_sc_hd__xnor2_1
X_06311_ _10926_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _06313_/A sky130_fd_sc_hd__nand2_1
X_07291_ _07366_/B _07291_/B _07291_/C vssd1 vssd1 vccd1 vccd1 _07369_/B sky130_fd_sc_hd__and3_1
XFILLER_164_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09030_ _10949_/Q _10432_/C _09008_/A _10933_/Q vssd1 vssd1 vccd1 vccd1 _09030_/X
+ sky130_fd_sc_hd__a22o_1
X_06242_ _10610_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06242_/X sky130_fd_sc_hd__or2_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06392__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06173_ _10592_/Q vssd1 vssd1 vccd1 vccd1 _06175_/A sky130_fd_sc_hd__inv_2
XFILLER_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09933_/B sky130_fd_sc_hd__nor2_1
XFILLER_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08168__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05736__A _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09208__A _09208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _09863_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__xnor2_1
XFILLER_140_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _08814_/A vssd1 vssd1 vccd1 vccd1 _08814_/X sky130_fd_sc_hd__clkbuf_2
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _09731_/A _09731_/B _09793_/X vssd1 vssd1 vccd1 vccd1 _09795_/B sky130_fd_sc_hd__a21o_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08745_ _08740_/X _08741_/X _08743_/Y _08744_/X vssd1 vssd1 vccd1 vccd1 _08759_/A
+ sky130_fd_sc_hd__o211a_1
X_05957_ input42/X vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__buf_6
XFILLER_39_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08676_ _08992_/A vssd1 vssd1 vccd1 vccd1 _08676_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05888_ _08180_/A _05888_/B vssd1 vssd1 vccd1 vccd1 _05888_/X sky130_fd_sc_hd__or2_1
XFILLER_42_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_39_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05471__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07715_/D _07627_/B vssd1 vssd1 vccd1 vccd1 _07628_/B sky130_fd_sc_hd__nand2_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07558_ _07557_/B _07558_/B vssd1 vssd1 vccd1 vccd1 _07559_/B sky130_fd_sc_hd__and2b_1
XFILLER_107_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06509_ _06510_/A _06510_/B vssd1 vssd1 vccd1 vccd1 _06511_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10435__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07489_ _07489_/A _07489_/B vssd1 vssd1 vccd1 vccd1 _07490_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07398__A _07728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09228_ _09228_/A _09228_/B vssd1 vssd1 vccd1 vccd1 _09229_/A sky130_fd_sc_hd__and2_1
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09159_ _05461_/A _09136_/X _09148_/X _05692_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09159_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10003_ _09930_/B _10123_/B _10139_/S _09716_/A vssd1 vssd1 vccd1 vccd1 _10003_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input21_A io_wbs_m2s_data[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08331__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10905_ _10926_/CLK _10905_/D vssd1 vssd1 vccd1 vccd1 _10905_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10836_ _10836_/CLK _10836_/D vssd1 vssd1 vccd1 vccd1 _10836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10767_ _10833_/CLK _10767_/D vssd1 vssd1 vccd1 vccd1 _10767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _10851_/CLK _10698_/D vssd1 vssd1 vccd1 vccd1 _10698_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_145_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06860_ _06860_/A _06860_/B vssd1 vssd1 vccd1 vccd1 _06862_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05811_ _05818_/A _05818_/B vssd1 vssd1 vccd1 vccd1 _05907_/A sky130_fd_sc_hd__nand2_1
X_06791_ _06792_/A _06792_/B vssd1 vssd1 vccd1 vccd1 _06833_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08530_ _10766_/Q _08419_/B _08529_/X vssd1 vssd1 vccd1 vccd1 _10766_/D sky130_fd_sc_hd__a21o_1
X_05742_ _05742_/A _05742_/B _05742_/C _05741_/Y vssd1 vssd1 vccd1 vccd1 _05788_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05291__A _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08461_ _08461_/A vssd1 vssd1 vccd1 vccd1 _10737_/D sky130_fd_sc_hd__clkbuf_1
X_05673_ _08251_/B _05602_/X _05599_/X _08251_/A _05672_/X vssd1 vssd1 vccd1 vccd1
+ _05673_/X sky130_fd_sc_hd__o221a_1
XFILLER_24_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07412_ _07412_/A _07412_/B _07412_/C vssd1 vssd1 vccd1 vccd1 _07413_/B sky130_fd_sc_hd__or3_1
XFILLER_51_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08395_/A _10754_/Q vssd1 vssd1 vccd1 vccd1 _08392_/X sky130_fd_sc_hd__or2_1
XFILLER_51_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07343_ _07528_/B _07528_/C _07528_/A vssd1 vssd1 vccd1 vccd1 _07529_/A sky130_fd_sc_hd__a21oi_2
XFILLER_10_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07274_ _07323_/B _07331_/A _07323_/A vssd1 vssd1 vccd1 vccd1 _07324_/A sky130_fd_sc_hd__a21o_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09013_ _09013_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _10341_/C sky130_fd_sc_hd__or2_1
X_06225_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06225_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06156_ _06156_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06156_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06087_ _08315_/A _08023_/A _05813_/A _05721_/Y vssd1 vssd1 vccd1 vccd1 _06087_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09915_ _09915_/A _09915_/B _09915_/C vssd1 vssd1 vccd1 vccd1 _09916_/B sky130_fd_sc_hd__nor3_1
XFILLER_58_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09846_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09848_/A sky130_fd_sc_hd__or2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09778_/B sky130_fd_sc_hd__and2_1
XFILLER_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _10979_/Q vssd1 vssd1 vccd1 vccd1 _07248_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08728_ _08830_/A vssd1 vssd1 vccd1 vccd1 _08728_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08659_/A vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__buf_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ _10653_/CLK _10621_/D vssd1 vssd1 vccd1 vccd1 _10621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _10554_/CLK _10552_/D vssd1 vssd1 vccd1 vccd1 _10552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10483_ _06143_/X _10475_/X _10482_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10965_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10187__A1 _09379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06000__A _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10819_ _10821_/CLK _10819_/D vssd1 vssd1 vccd1 vccd1 _10819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08068__B1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10457__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06010_ _08236_/A vssd1 vssd1 vccd1 vccd1 _06011_/A sky130_fd_sc_hd__inv_2
XFILLER_145_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07766__A _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10192__A _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07961_ _10537_/A _06050_/X _07983_/A vssd1 vssd1 vccd1 vccd1 _07962_/B sky130_fd_sc_hd__mux2_1
XFILLER_87_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09700_ _09769_/A _09810_/B _09769_/B _09764_/A vssd1 vssd1 vccd1 vccd1 _09701_/B
+ sky130_fd_sc_hd__a22o_1
X_06912_ _06916_/A _06912_/B vssd1 vssd1 vccd1 vccd1 _06923_/B sky130_fd_sc_hd__xor2_4
X_07892_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07892_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08597__A _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ _09631_/A _09631_/B _09631_/C vssd1 vssd1 vccd1 vccd1 _09631_/X sky130_fd_sc_hd__or3_1
XFILLER_95_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06843_ _10513_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _06848_/A sky130_fd_sc_hd__nand2_1
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10350__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09562_ _09562_/A _09562_/B _09562_/C vssd1 vssd1 vccd1 vccd1 _09563_/A sky130_fd_sc_hd__nand3_1
X_06774_ _06785_/A _06774_/B vssd1 vssd1 vccd1 vccd1 _06775_/C sky130_fd_sc_hd__and2_1
XFILLER_83_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07006__A _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08513_ _10794_/Q vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05725_ _10548_/Q vssd1 vssd1 vccd1 vccd1 _05739_/B sky130_fd_sc_hd__inv_2
X_09493_ _09454_/A _09454_/B _09390_/A vssd1 vssd1 vccd1 vccd1 _09494_/D sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08444_ _08444_/A vssd1 vssd1 vccd1 vccd1 _10732_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05656_ _06037_/A _05636_/Y _05632_/Y _10686_/Q _05655_/X vssd1 vssd1 vccd1 vccd1
+ _05656_/X sky130_fd_sc_hd__o221a_1
XFILLER_24_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08375_ _08367_/X _10731_/Q _07865_/X _08374_/X vssd1 vssd1 vccd1 vccd1 _10713_/D
+ sky130_fd_sc_hd__o211a_1
X_05587_ _10564_/Q _05593_/A _10565_/Q vssd1 vssd1 vccd1 vccd1 _05588_/B sky130_fd_sc_hd__o21ai_1
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07326_ _07326_/A vssd1 vssd1 vccd1 vccd1 _07562_/A sky130_fd_sc_hd__buf_2
XFILLER_164_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07257_ _07275_/A _07275_/B vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__nor2_1
XFILLER_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06208_ _10341_/A vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__buf_4
XFILLER_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07188_ _07188_/A _07188_/B _07188_/C vssd1 vssd1 vccd1 vccd1 _07190_/A sky130_fd_sc_hd__and3_1
XFILLER_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06139_ _10585_/Q vssd1 vssd1 vccd1 vccd1 _06140_/A sky130_fd_sc_hd__inv_2
XFILLER_155_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09829_ _09829_/A _10023_/A vssd1 vssd1 vccd1 vccd1 _09974_/A sky130_fd_sc_hd__or2_1
XFILLER_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09131__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _10822_/CLK _10604_/D vssd1 vssd1 vccd1 vccd1 _10604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10535_ _10535_/A _10537_/B _10537_/C vssd1 vssd1 vccd1 vccd1 _10535_/X sky130_fd_sc_hd__or3_1
XFILLER_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10466_ _06191_/X _10459_/X _10465_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10959_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10397_ _10389_/X _10718_/Q _10394_/X _10396_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10937_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output52_A _10581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05510_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05510_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06490_ _10974_/Q vssd1 vssd1 vccd1 vccd1 _06568_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05441_ _10673_/Q _05844_/B _08318_/A vssd1 vssd1 vccd1 vccd1 _05442_/B sky130_fd_sc_hd__o21ai_1
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08160_ _08160_/A _08160_/B vssd1 vssd1 vccd1 vccd1 _08173_/B sky130_fd_sc_hd__nor2_1
X_05372_ _10628_/Q vssd1 vssd1 vccd1 vccd1 _05460_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07111_ _07150_/A vssd1 vssd1 vccd1 vccd1 _07135_/A sky130_fd_sc_hd__inv_2
XFILLER_119_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _08091_/A vssd1 vssd1 vccd1 vccd1 _10683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07042_ _07042_/A _07042_/B vssd1 vssd1 vccd1 vccd1 _07043_/B sky130_fd_sc_hd__nor2_1
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08213__B1 _08124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08993_ _08970_/X _08983_/X _08991_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10834_/D
+ sky130_fd_sc_hd__o31a_2
XFILLER_134_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07944_ input38/X _06065_/X _07964_/A vssd1 vssd1 vccd1 vccd1 _07945_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07875_ _07875_/A vssd1 vssd1 vccd1 vccd1 _07875_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09614_ _09656_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06826_ _07682_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _06856_/C sky130_fd_sc_hd__nand2_2
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09545_ _09617_/B _09545_/B vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__xor2_1
X_06757_ _06758_/A _06758_/C _06786_/A _06769_/A vssd1 vssd1 vccd1 vccd1 _06759_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_70_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05708_ _05708_/A _05708_/B vssd1 vssd1 vccd1 vccd1 _05708_/Y sky130_fd_sc_hd__nand2_1
X_09476_ _09476_/A _09476_/B vssd1 vssd1 vccd1 vccd1 _09479_/A sky130_fd_sc_hd__nand2_1
XFILLER_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06688_ _06688_/A _06688_/B vssd1 vssd1 vccd1 vccd1 _06690_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08427_ _10782_/Q _10781_/Q _10780_/Q _10779_/Q vssd1 vssd1 vccd1 vccd1 _08432_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05639_ _10682_/Q vssd1 vssd1 vccd1 vccd1 _05719_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10097__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08358_ _05528_/A _08349_/X _08092_/A vssd1 vssd1 vccd1 vccd1 _08358_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_149_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07309_ _07309_/A _07309_/B _07309_/C vssd1 vssd1 vccd1 vccd1 _07310_/B sky130_fd_sc_hd__and3_1
XFILLER_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08289_ _08289_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08289_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10320_ _10320_/A _10320_/B vssd1 vssd1 vccd1 vccd1 _10320_/X sky130_fd_sc_hd__xor2_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10251_ _10249_/Y _10250_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _10252_/B sky130_fd_sc_hd__mux2_1
XFILLER_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06215__C1 _06200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10182_ _07008_/A _10181_/X _10177_/X _10892_/Q vssd1 vssd1 vccd1 vccd1 _10892_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08030__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09180__B2 _08191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06297__A2 _09356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10518_ _10537_/B _10518_/B vssd1 vssd1 vccd1 vccd1 _10522_/A sky130_fd_sc_hd__nor2_1
XFILLER_156_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10449_ _05982_/A _10446_/X _10448_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10952_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10470__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05990_ _08462_/A vssd1 vssd1 vccd1 vccd1 _07899_/A sky130_fd_sc_hd__buf_2
XFILLER_85_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09171__A1 _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07660_ _07668_/A _07667_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07661_/B sky130_fd_sc_hd__o21ai_1
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06611_ _06856_/A _06522_/B _06513_/D _06769_/A vssd1 vssd1 vccd1 vccd1 _06612_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_80_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07591_ _09420_/A _07475_/B _07475_/C vssd1 vssd1 vccd1 vccd1 _07592_/B sky130_fd_sc_hd__o21ai_1
XFILLER_53_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _10965_/Q _09536_/B vssd1 vssd1 vccd1 vccd1 _09451_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06542_ _06542_/A _06542_/B vssd1 vssd1 vccd1 vccd1 _06544_/A sky130_fd_sc_hd__xnor2_1
X_09261_ _10441_/A vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__clkbuf_1
X_06473_ _06670_/A _06670_/B vssd1 vssd1 vccd1 vccd1 _06671_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08212_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08212_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05424_ _05460_/C _05369_/Y _05366_/Y _10630_/Q _05423_/X vssd1 vssd1 vccd1 vccd1
+ _05424_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09192_ _09112_/A _09188_/Y _09191_/X vssd1 vssd1 vccd1 vccd1 _09193_/B sky130_fd_sc_hd__a21oi_1
XFILLER_147_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08143_ input46/X _08086_/X _08109_/X _06035_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08144_/B sky130_fd_sc_hd__o221a_1
X_05355_ _10664_/Q vssd1 vssd1 vccd1 vccd1 _06052_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08074_ _08074_/A vssd1 vssd1 vccd1 vccd1 _08074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05286_ _10649_/Q _05286_/B vssd1 vssd1 vccd1 vccd1 _05406_/A sky130_fd_sc_hd__nor2_1
XFILLER_161_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07025_ _07044_/A _07039_/C vssd1 vssd1 vccd1 vccd1 _07025_/Y sky130_fd_sc_hd__nand2_1
XFILLER_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08976_ _08976_/A vssd1 vssd1 vccd1 vccd1 _08976_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05474__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07927_ _08284_/A _07927_/B vssd1 vssd1 vccd1 vccd1 _10646_/D sky130_fd_sc_hd__nor2_1
XFILLER_130_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06289__B _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07858_ _07848_/X _05461_/A _07844_/X _07857_/Y vssd1 vssd1 vccd1 vccd1 _10627_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_84_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06809_ _10911_/Q vssd1 vssd1 vccd1 vccd1 _07570_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__05723__A1 _05721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07789_ _07789_/A _07789_/B vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__nand2_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05723__B2 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _09479_/A _09479_/B _09476_/A vssd1 vssd1 vccd1 vccd1 _09529_/B sky130_fd_sc_hd__o21ai_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08122__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _09458_/B _09458_/C _09458_/A vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__a21o_1
XFILLER_52_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10303_ _10303_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10303_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_153_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input51_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _10936_/Q _10952_/Q vssd1 vssd1 vccd1 vccd1 _10235_/B sky130_fd_sc_hd__or2b_1
XFILLER_152_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10165_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10165_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_67_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10096_ _10097_/A _10097_/B vssd1 vssd1 vccd1 vccd1 _10098_/A sky130_fd_sc_hd__nor2_1
XFILLER_102_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08830_ _08830_/A vssd1 vssd1 vccd1 vccd1 _08830_/X sky130_fd_sc_hd__clkbuf_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05294__A _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08804_/B _08760_/X _08804_/A vssd1 vssd1 vccd1 vccd1 _08761_/Y sky130_fd_sc_hd__o21ai_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05973_ _10432_/B _08981_/A vssd1 vssd1 vccd1 vccd1 _06120_/S sky130_fd_sc_hd__nand2_2
XFILLER_100_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07712_ _07601_/A _07601_/B _07711_/X vssd1 vssd1 vccd1 vccd1 _07757_/A sky130_fd_sc_hd__o21ba_2
XFILLER_39_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08692_ _08679_/X _08692_/B vssd1 vssd1 vccd1 vccd1 _08693_/B sky130_fd_sc_hd__and2b_1
XFILLER_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07643_ _07643_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07647_/A sky130_fd_sc_hd__xnor2_4
XFILLER_38_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07574_ _07574_/A _07574_/B _07574_/C vssd1 vssd1 vccd1 vccd1 _07576_/A sky130_fd_sc_hd__and3_1
XFILLER_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09313_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09314_/B sky130_fd_sc_hd__nor2_1
X_06525_ _06620_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _06621_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09244_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09244_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06456_ _06456_/A _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06465_/A sky130_fd_sc_hd__and3_1
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05407_ _10617_/Q _05480_/A vssd1 vssd1 vccd1 vccd1 _05407_/X sky130_fd_sc_hd__or2_1
X_09175_ _10960_/Q _09194_/B vssd1 vssd1 vccd1 vccd1 _09175_/Y sky130_fd_sc_hd__nor2_1
X_06387_ _06387_/A _06387_/B vssd1 vssd1 vccd1 vccd1 _06412_/B sky130_fd_sc_hd__or2_1
XANTENNA__10375__A _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08126_ _10535_/A _08123_/X _08124_/X _08117_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08127_/B sky130_fd_sc_hd__o221a_1
X_05338_ _10639_/Q vssd1 vssd1 vccd1 vccd1 _07900_/A sky130_fd_sc_hd__clkbuf_2
X_08057_ _08352_/B vssd1 vssd1 vccd1 vccd1 _08058_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_35_clock_A _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05269_ _10679_/Q vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__clkinv_4
XFILLER_162_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07008_ _07008_/A _07008_/B vssd1 vssd1 vccd1 vccd1 _07030_/C sky130_fd_sc_hd__xnor2_2
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput59 _10846_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[12] sky130_fd_sc_hd__buf_2
XFILLER_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08959_ _09736_/B vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08343__C1 _08062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10921_ _10930_/CLK _10921_/D vssd1 vssd1 vccd1 vccd1 _10921_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10852_ _10857_/CLK _10852_/D vssd1 vssd1 vccd1 vccd1 _10852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10783_ _10790_/CLK _10783_/D vssd1 vssd1 vccd1 vccd1 _10783_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08110__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10217_ _10202_/X _10206_/Y _10203_/X vssd1 vssd1 vccd1 vccd1 _10217_/X sky130_fd_sc_hd__a21bo_1
XFILLER_122_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10148_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10152_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10079_ _10079_/A _10079_/B vssd1 vssd1 vccd1 vccd1 _10081_/C sky130_fd_sc_hd__xnor2_1
XFILLER_47_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08334__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06310_ _06730_/A _06730_/B _06730_/C _06731_/B vssd1 vssd1 vccd1 vccd1 _06734_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__10444__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07290_ _07287_/A _07287_/B _07289_/X vssd1 vssd1 vccd1 vccd1 _07291_/C sky130_fd_sc_hd__a21bo_1
X_06241_ input33/X _06238_/X _06240_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10609_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_61_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10655_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06172_ input46/X vssd1 vssd1 vccd1 vccd1 _06172_/X sky130_fd_sc_hd__buf_4
XFILLER_8_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09062__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10985_/CLK sky130_fd_sc_hd__clkbuf_16
X_09931_ _09931_/A _10139_/S vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _09346_/B _09797_/B _09861_/X vssd1 vssd1 vccd1 vccd1 _09863_/B sky130_fd_sc_hd__o21a_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08813_ _08810_/X _08812_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10815_/D sky130_fd_sc_hd__a21oi_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09793_ _09730_/B _09793_/B vssd1 vssd1 vccd1 vccd1 _09793_/X sky130_fd_sc_hd__and2b_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05926__B2 _05692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05956_ _05956_/A vssd1 vssd1 vccd1 vccd1 _05956_/X sky130_fd_sc_hd__clkbuf_1
X_08744_ _10807_/Q _08744_/B vssd1 vssd1 vccd1 vccd1 _08744_/X sky130_fd_sc_hd__or2_1
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _06008_/A _08672_/X _08674_/X _10800_/Q vssd1 vssd1 vccd1 vccd1 _08675_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05887_ _07985_/A _05886_/Y _05883_/X vssd1 vssd1 vccd1 vccd1 _05888_/B sky130_fd_sc_hd__o21a_1
XFILLER_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07626_ _07700_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__xor2_2
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_clock clkbuf_opt_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _10850_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07557_ _07558_/B _07557_/B vssd1 vssd1 vccd1 vccd1 _07724_/A sky130_fd_sc_hd__and2b_1
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06508_ _06519_/A _06508_/B vssd1 vssd1 vccd1 vccd1 _06510_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07488_ _07488_/A _07488_/B _07529_/A vssd1 vssd1 vccd1 vccd1 _07489_/B sky130_fd_sc_hd__or3_1
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10945_/CLK sky130_fd_sc_hd__clkbuf_16
X_09227_ _10818_/Q _09210_/X _09212_/X _09226_/X _09203_/X vssd1 vssd1 vccd1 vccd1
+ _09228_/B sky130_fd_sc_hd__a32o_1
X_06439_ _10975_/Q _06561_/C _06440_/A _06461_/B vssd1 vssd1 vccd1 vccd1 _06442_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09158_ _09113_/X _09157_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09158_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_147_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08109_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08109_/X sky130_fd_sc_hd__clkbuf_2
X_09089_ _09081_/X _09088_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10840_/D sky130_fd_sc_hd__o21a_2
XFILLER_163_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ _10484_/A _10139_/S vssd1 vssd1 vccd1 vccd1 _10078_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08564__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09108__B2 _10719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input14_A io_wbs_m2s_addr[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10904_ _10929_/CLK _10904_/D vssd1 vssd1 vccd1 vccd1 _10904_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10835_ _10835_/CLK _10835_/D vssd1 vssd1 vccd1 vccd1 _10835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09292__A0 _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10766_ _10804_/CLK _10766_/D vssd1 vssd1 vccd1 vccd1 _10766_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ _10851_/CLK _10697_/D vssd1 vssd1 vccd1 vccd1 _10697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05810_ _10652_/Q vssd1 vssd1 vccd1 vccd1 _05905_/A sky130_fd_sc_hd__buf_2
XFILLER_83_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06790_ _06772_/A _06762_/A _07773_/B _06856_/A vssd1 vssd1 vccd1 vccd1 _06792_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08307__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05741_ _08059_/A _05741_/B vssd1 vssd1 vccd1 vccd1 _05741_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08322__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08460_ _08460_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__or2_1
X_05672_ _10699_/Q _05602_/X _05605_/X _05671_/X vssd1 vssd1 vccd1 vccd1 _05672_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07411_ _07412_/B _07412_/C _07412_/A vssd1 vssd1 vccd1 vccd1 _07549_/A sky130_fd_sc_hd__o21ai_1
XFILLER_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08391_ _08383_/X _10737_/Q _08380_/X _08390_/X vssd1 vssd1 vccd1 vccd1 _10719_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07342_ _07488_/B _07342_/B vssd1 vssd1 vccd1 vccd1 _07528_/A sky130_fd_sc_hd__or2_1
X_07273_ _07273_/A _07273_/B vssd1 vssd1 vccd1 vccd1 _07323_/A sky130_fd_sc_hd__xnor2_1
XFILLER_136_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09012_ _10480_/A _09009_/X _09086_/S vssd1 vssd1 vccd1 vccd1 _09012_/X sky130_fd_sc_hd__mux2_1
X_06224_ input26/X _06207_/X _06223_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10603_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06155_ _10588_/Q vssd1 vssd1 vccd1 vccd1 _06156_/A sky130_fd_sc_hd__inv_2
XFILLER_132_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09219__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06086_ _08093_/A _05291_/A _06065_/X _06066_/Y _06085_/X vssd1 vssd1 vccd1 vccd1
+ _06089_/C sky130_fd_sc_hd__a221o_1
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09914_ _09915_/A _09915_/B _09915_/C vssd1 vssd1 vccd1 vccd1 _09916_/A sky130_fd_sc_hd__o21a_1
XFILLER_59_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08010__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07962__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09901_/A sky130_fd_sc_hd__xnor2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input6_A io_wbs_m2s_addr[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09851_/A sky130_fd_sc_hd__nor2_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06988_ _07563_/A _07433_/A vssd1 vssd1 vccd1 vccd1 _07562_/C sky130_fd_sc_hd__nand2_2
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08727_ _08740_/A _08724_/X _08740_/B _08726_/Y _08658_/X vssd1 vssd1 vccd1 vccd1
+ _08727_/X sky130_fd_sc_hd__o311a_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05939_ _05771_/A _05841_/X _05940_/B _08315_/B _05938_/X vssd1 vssd1 vccd1 vccd1
+ _05939_/X sky130_fd_sc_hd__a221o_1
XANTENNA__08849__B1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _08778_/A vssd1 vssd1 vccd1 vccd1 _08658_/X sky130_fd_sc_hd__buf_2
XFILLER_26_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07609_ _07609_/A _07609_/B vssd1 vssd1 vccd1 vccd1 _07706_/B sky130_fd_sc_hd__xnor2_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08589_ _10782_/Q _08586_/B _08588_/Y vssd1 vssd1 vccd1 vccd1 _10782_/D sky130_fd_sc_hd__o21a_1
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10620_ _10652_/CLK _10620_/D vssd1 vssd1 vccd1 vccd1 _10620_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08077__A1 _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10551_ _10654_/CLK _10551_/D vssd1 vssd1 vccd1 vccd1 _10551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10482_ _10482_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10482_/X sky130_fd_sc_hd__or2_1
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08001__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06012__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10818_ _10822_/CLK _10818_/D vssd1 vssd1 vccd1 vccd1 _10818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08208__A _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06079__B1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10354__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10749_ _10776_/CLK _10749_/D vssd1 vssd1 vccd1 vccd1 _10749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07960_ _07960_/A vssd1 vssd1 vccd1 vccd1 _10654_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06911_ _06748_/X _06771_/B _06910_/X vssd1 vssd1 vccd1 vccd1 _06913_/A sky130_fd_sc_hd__a21bo_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07891_ _07898_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _10636_/D sky130_fd_sc_hd__nor2_1
XFILLER_96_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09630_ _09686_/A _09630_/B vssd1 vssd1 vccd1 vccd1 _09631_/C sky130_fd_sc_hd__nor2_1
X_06842_ _06842_/A vssd1 vssd1 vccd1 vccd1 _07776_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_110_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09561_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06773_ _06900_/A _06842_/A _06773_/C vssd1 vssd1 vccd1 vccd1 _06902_/A sky130_fd_sc_hd__and3_2
XFILLER_64_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05724_ _10687_/Q vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__clkbuf_2
X_08512_ _10793_/Q _08506_/X _08509_/X _10756_/Q vssd1 vssd1 vccd1 vccd1 _10756_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09492_ _09492_/A vssd1 vssd1 vccd1 vccd1 _09696_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05655_ _10685_/Q _05636_/Y _05637_/Y _08095_/A _05654_/X vssd1 vssd1 vccd1 vccd1
+ _05655_/X sky130_fd_sc_hd__a221o_1
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__or2_1
XFILLER_51_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09256__A0 _08297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _08381_/A _10747_/Q vssd1 vssd1 vccd1 vccd1 _08374_/X sky130_fd_sc_hd__or2_1
X_05586_ _10704_/Q vssd1 vssd1 vccd1 vccd1 _05771_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07325_ _07338_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07528_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07256_ _07230_/X _07256_/B vssd1 vssd1 vccd1 vccd1 _07275_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07957__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06207_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06207_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07187_ _07201_/A _07187_/B vssd1 vssd1 vccd1 vccd1 _07188_/C sky130_fd_sc_hd__xnor2_1
XFILLER_118_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06138_ _06124_/X _06131_/X _06134_/Y _06137_/X vssd1 vssd1 vccd1 vccd1 _10584_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06069_ _06062_/X _06063_/X _06069_/C _06069_/D vssd1 vssd1 vccd1 vccd1 _06070_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09828_ _09977_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _10023_/A sky130_fd_sc_hd__nand2_1
XFILLER_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09819_/A sky130_fd_sc_hd__xor2_2
XFILLER_62_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10603_ _10666_/CLK _10603_/D vssd1 vssd1 vccd1 vccd1 _10603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05808__B1 _05528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10534_ _07727_/A _10522_/X _10533_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10984_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_127_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10465_ _10959_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10465_/X sky130_fd_sc_hd__or2_1
XANTENNA__10293__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08222__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10396_ _10937_/Q _10379_/B _10395_/X vssd1 vssd1 vccd1 vccd1 _10396_/X sky130_fd_sc_hd__a21bo_1
XFILLER_124_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_83_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09322__A _09323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05440_ _10674_/Q vssd1 vssd1 vccd1 vccd1 _08318_/A sky130_fd_sc_hd__buf_2
XANTENNA__09238__A0 _08268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05371_ _07985_/A _05374_/A vssd1 vssd1 vccd1 vccd1 _05371_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_158_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07110_ _10983_/Q _07125_/A vssd1 vssd1 vccd1 vccd1 _07150_/A sky130_fd_sc_hd__nand2_1
XFILLER_119_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08090_ _08090_/A _08090_/B vssd1 vssd1 vccd1 vccd1 _08091_/A sky130_fd_sc_hd__and2_1
XFILLER_147_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07041_ _07424_/A _07041_/B vssd1 vssd1 vccd1 vccd1 _07048_/A sky130_fd_sc_hd__nor2_1
XFILLER_161_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09992__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08213__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08213__B2 _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _08992_/A vssd1 vssd1 vccd1 vccd1 _08992_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_115_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07943_ _07943_/A vssd1 vssd1 vccd1 vccd1 _10649_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07874_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07874_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09613_ _09613_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09614_/B sky130_fd_sc_hd__or3_1
X_06825_ _06845_/A _06842_/A vssd1 vssd1 vccd1 vccd1 _06844_/C sky130_fd_sc_hd__nand2_1
XFILLER_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _09501_/A _09501_/C _09501_/B vssd1 vssd1 vccd1 vccd1 _09545_/B sky130_fd_sc_hd__a21boi_1
XFILLER_37_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06756_ _06756_/A _06806_/B vssd1 vssd1 vccd1 vccd1 _06786_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09232__A _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05707_ _05702_/A _10556_/Q _10555_/Q _08196_/A vssd1 vssd1 vccd1 vccd1 _05708_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_169_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09475_ _09475_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09476_/B sky130_fd_sc_hd__nand2_1
X_06687_ _06941_/B _06944_/A _06941_/A vssd1 vssd1 vccd1 vccd1 _06942_/A sky130_fd_sc_hd__a21oi_2
XFILLER_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08426_ _10778_/Q _10777_/Q _10776_/Q _10775_/Q vssd1 vssd1 vccd1 vccd1 _08432_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05638_ _10684_/Q vssd1 vssd1 vccd1 vccd1 _08095_/A sky130_fd_sc_hd__clkbuf_2
X_05569_ _10709_/Q vssd1 vssd1 vccd1 vccd1 _08339_/A sky130_fd_sc_hd__clkbuf_2
X_08357_ _08881_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _10710_/D sky130_fd_sc_hd__nor2_1
XFILLER_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07308_ _07308_/A _07319_/A _07308_/C vssd1 vssd1 vccd1 vccd1 _07344_/B sky130_fd_sc_hd__or3_1
XFILLER_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08288_ _08278_/A _08278_/B _08287_/A vssd1 vssd1 vccd1 vccd1 _08288_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_109_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07239_ _07235_/C _07382_/A _07224_/X vssd1 vssd1 vccd1 vccd1 _07239_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_165_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10250_ _10235_/B _10237_/Y _10233_/X vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__a21o_1
XFILLER_106_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10181_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10181_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_161_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_3_0_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10517_ _10517_/A vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10448_ _10952_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10448_/X sky130_fd_sc_hd__or2_1
XFILLER_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07954__A0 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10379_ _10933_/Q _10379_/B vssd1 vssd1 vccd1 vccd1 _10379_/X sky130_fd_sc_hd__and2_1
XANTENNA__06757__B2 _06769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09317__A _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06610_ _06758_/B vssd1 vssd1 vccd1 vccd1 _06769_/A sky130_fd_sc_hd__buf_2
X_07590_ _10901_/Q vssd1 vssd1 vccd1 vccd1 _09420_/A sky130_fd_sc_hd__clkinv_2
XFILLER_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06541_ _06785_/A _06719_/C _06541_/C vssd1 vssd1 vccd1 vccd1 _06542_/B sky130_fd_sc_hd__and3_1
XFILLER_52_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10198__A _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06472_ _06472_/A _06472_/B vssd1 vssd1 vccd1 vccd1 _06670_/B sky130_fd_sc_hd__xnor2_1
X_09260_ _09260_/A vssd1 vssd1 vccd1 vccd1 _10858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05423_ _10629_/Q _05369_/Y _05371_/Y _05460_/D _05422_/X vssd1 vssd1 vccd1 vccd1
+ _05423_/X sky130_fd_sc_hd__a221o_1
X_08211_ _08114_/X _08224_/C _08207_/Y _08210_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08211_/X sky130_fd_sc_hd__o311a_1
X_09191_ _10813_/Q _09168_/X _09079_/X _10726_/Q _09190_/X vssd1 vssd1 vccd1 vccd1
+ _09191_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ _07974_/A _08044_/A _08141_/X vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__a21o_1
X_05354_ _10633_/Q vssd1 vssd1 vccd1 vccd1 _07878_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08073_ _08038_/X _08065_/B _08072_/Y _06033_/X vssd1 vssd1 vccd1 vccd1 _08073_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_147_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05285_ _10573_/Q vssd1 vssd1 vccd1 vccd1 _05286_/B sky130_fd_sc_hd__inv_2
XFILLER_174_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07024_ _07169_/A vssd1 vssd1 vccd1 vccd1 _07044_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08975_ _08995_/A vssd1 vssd1 vccd1 vccd1 _08976_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07926_ _10614_/Q _07906_/A _07910_/X _07925_/Y vssd1 vssd1 vccd1 vccd1 _07927_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_29_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07857_ _06189_/A _07849_/X _07850_/X _07856_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ _07857_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_110_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06808_ _07670_/A _06853_/A vssd1 vssd1 vccd1 vccd1 _06814_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07788_ _06741_/A _06833_/A _06833_/B _06834_/B vssd1 vssd1 vccd1 vccd1 _07789_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05490__A _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09527_ _09527_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06739_ _06758_/C vssd1 vssd1 vccd1 vccd1 _07784_/B sky130_fd_sc_hd__clkbuf_2
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09458_ _09458_/A _09458_/B _09458_/C vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__nand3_1
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08409_ _08397_/X _10744_/Q _08992_/A _08408_/X vssd1 vssd1 vccd1 vccd1 _10726_/D
+ sky130_fd_sc_hd__o211a_1
X_09389_ _10964_/Q _09396_/A _09411_/A vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__and3_1
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10232__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08025__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _10299_/X _10301_/Y _10329_/S vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__mux2_1
XFILLER_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10233_ _10952_/Q _10936_/Q vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__and2b_1
XFILLER_161_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10164_ _10164_/A _10164_/B vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_input44_A io_wbs_m2s_data[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10095_ _10095_/A _10095_/B vssd1 vssd1 vccd1 vccd1 _10097_/B sky130_fd_sc_hd__xor2_1
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07880__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08760_ _10808_/Q _08748_/X _08928_/B vssd1 vssd1 vccd1 vccd1 _08760_/X sky130_fd_sc_hd__o21a_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05972_ _09107_/B vssd1 vssd1 vccd1 vccd1 _08981_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07711_ _07603_/A _07711_/B vssd1 vssd1 vccd1 vccd1 _07711_/X sky130_fd_sc_hd__and2b_1
XFILLER_66_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08691_ _08689_/Y _08691_/B vssd1 vssd1 vccd1 vccd1 _08693_/A sky130_fd_sc_hd__and2b_1
XFILLER_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07642_ _07527_/B _07648_/B _07655_/A vssd1 vssd1 vccd1 vccd1 _07643_/B sky130_fd_sc_hd__o21ai_2
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07573_ _07573_/A _07726_/B _07573_/C vssd1 vssd1 vccd1 vccd1 _07574_/C sky130_fd_sc_hd__and3_1
XFILLER_81_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09312_ _10351_/A vssd1 vssd1 vccd1 vccd1 _09312_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06524_ _06520_/X _06602_/A _06545_/A vssd1 vssd1 vccd1 vccd1 _06620_/B sky130_fd_sc_hd__a21oi_1
XFILLER_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09243_ _09274_/A vssd1 vssd1 vccd1 vccd1 _09243_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10462__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06455_ _06468_/A _06450_/B _06478_/A vssd1 vssd1 vccd1 vccd1 _06458_/A sky130_fd_sc_hd__a21o_1
XFILLER_167_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05406_ _05406_/A _05406_/B vssd1 vssd1 vccd1 vccd1 _05480_/A sky130_fd_sc_hd__nor2_1
X_06386_ _06386_/A _06386_/B vssd1 vssd1 vccd1 vccd1 _06412_/A sky130_fd_sc_hd__xor2_4
X_09174_ _09202_/A _09174_/B vssd1 vssd1 vccd1 vccd1 _10846_/D sky130_fd_sc_hd__nor2_4
XFILLER_147_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07030__A _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05337_ _07903_/A _05337_/B vssd1 vssd1 vccd1 vccd1 _05337_/X sky130_fd_sc_hd__or2_1
X_08125_ _08201_/A vssd1 vssd1 vccd1 vccd1 _08125_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07965__A _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _08039_/X _08045_/X _08055_/X vssd1 vssd1 vccd1 vccd1 _10680_/D sky130_fd_sc_hd__o21a_1
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07007_ _07007_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07008_/B sky130_fd_sc_hd__nand2_1
XFILLER_116_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08958_ _09867_/B vssd1 vssd1 vccd1 vccd1 _09736_/B sky130_fd_sc_hd__buf_2
XFILLER_57_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07909_ _07916_/A _07909_/B vssd1 vssd1 vccd1 vccd1 _10641_/D sky130_fd_sc_hd__nor2_1
XFILLER_5_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08889_ _08889_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _08889_/X sky130_fd_sc_hd__and2_1
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10920_ _10930_/CLK _10920_/D vssd1 vssd1 vccd1 vccd1 _10920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08894__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10851_ _10851_/CLK _10851_/D vssd1 vssd1 vccd1 vccd1 _10851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10782_/CLK _10782_/D vssd1 vssd1 vccd1 vccd1 _10782_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10453__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08031__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10216_ _10203_/X _10226_/A _10202_/X vssd1 vssd1 vccd1 vccd1 _10216_/X sky130_fd_sc_hd__a21bo_1
XFILLER_122_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10147_ _10049_/C _10050_/A _09976_/Y vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__a21o_1
XFILLER_95_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10078_ _10078_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _10079_/B sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_1_0_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08885__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10444__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10476__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06240_ _10609_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06240_/X sky130_fd_sc_hd__or2_1
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06171_ _06168_/X _06158_/X _06170_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10591_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09930_ _09856_/C _09930_/B _09930_/C vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__nand3b_1
XFILLER_131_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ _10892_/Q _07008_/A vssd1 vssd1 vccd1 vccd1 _09861_/X sky130_fd_sc_hd__or2b_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08812_ input23/X _08672_/X _08674_/X hold13/A vssd1 vssd1 vccd1 vccd1 _08812_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09792_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__xor2_4
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _10807_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08743_/Y sky130_fd_sc_hd__nand2_1
X_05955_ _06019_/A _10728_/Q vssd1 vssd1 vccd1 vccd1 _05956_/A sky130_fd_sc_hd__and2_4
XFILLER_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08325__B1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _08831_/A vssd1 vssd1 vccd1 vccd1 _08674_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05886_ _05886_/A _05886_/B vssd1 vssd1 vccd1 vccd1 _05886_/Y sky130_fd_sc_hd__nor2_1
X_07625_ _07625_/A _07625_/B vssd1 vssd1 vccd1 vccd1 _07700_/B sky130_fd_sc_hd__xor2_4
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08089__C1 _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ _07556_/A _07556_/B vssd1 vssd1 vccd1 vccd1 _07557_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06507_ _06507_/A _06521_/A vssd1 vssd1 vccd1 vccd1 _06508_/B sky130_fd_sc_hd__or2_1
XFILLER_139_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07487_ _07495_/A _07495_/B vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10386__A _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09226_ _08244_/A _09225_/X _09226_/S vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__mux2_1
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06438_ _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06440_/A sky130_fd_sc_hd__and2_1
XFILLER_155_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09157_ _09114_/X _09156_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10199__B1 _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06369_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _06896_/A sky130_fd_sc_hd__and2_1
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09053__B2 _08098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08108_ _06038_/X _08043_/A _08103_/Y _08038_/A _08107_/X vssd1 vssd1 vccd1 vccd1
+ _08111_/A sky130_fd_sc_hd__a221o_1
X_09088_ _07729_/A _09087_/X _10537_/C vssd1 vssd1 vccd1 vccd1 _09088_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08039_ _08074_/A _08065_/B _05736_/A _08038_/X vssd1 vssd1 vccd1 vccd1 _08039_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10001_ _10076_/A _10001_/B vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__xnor2_1
XFILLER_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08316__B1 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10903_ _10926_/CLK _10903_/D vssd1 vssd1 vccd1 vccd1 _10903_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10834_ _10987_/CLK _10834_/D vssd1 vssd1 vccd1 vccd1 _10834_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_32_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10765_ _10807_/CLK _10765_/D vssd1 vssd1 vccd1 vccd1 _10765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_160_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ _10851_/CLK _10696_/D vssd1 vssd1 vccd1 vccd1 _10696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09296__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06014__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10362__B1 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06030__A1 _10581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05740_ _08082_/C vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05671_ _10698_/Q _05605_/B _05606_/X _08224_/A _05670_/X vssd1 vssd1 vccd1 vccd1
+ _05671_/X sky130_fd_sc_hd__a221o_1
XFILLER_36_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07410_ _07410_/A _07410_/B vssd1 vssd1 vccd1 vccd1 _07412_/A sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_78_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ _08395_/A _10753_/Q vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__or2_1
XFILLER_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07341_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07342_/B sky130_fd_sc_hd__and2_1
XFILLER_32_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07272_ _07330_/A _07335_/A vssd1 vssd1 vccd1 vccd1 _07331_/A sky130_fd_sc_hd__or2_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09011_ _09194_/B _10432_/C vssd1 vssd1 vccd1 vccd1 _09086_/S sky130_fd_sc_hd__nand2_1
X_06223_ _10603_/Q _06223_/B vssd1 vssd1 vccd1 vccd1 _06223_/X sky130_fd_sc_hd__or2_1
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06154_ _06147_/X _06131_/X _06151_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10587_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06085_ _08188_/A _07988_/A vssd1 vssd1 vccd1 vccd1 _06085_/X sky130_fd_sc_hd__xor2_1
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09913_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09915_/C sky130_fd_sc_hd__xor2_1
XFILLER_99_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09844_ _09844_/A _09844_/B _09844_/C vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__and3_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09775_ _09775_/A _09843_/A vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__xor2_1
XFILLER_85_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06987_ _07020_/B vssd1 vssd1 vccd1 vccd1 _07433_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08726_ _08724_/X _08740_/B _08740_/A vssd1 vssd1 vccd1 vccd1 _08726_/Y sky130_fd_sc_hd__o21ai_1
X_05938_ _08285_/A _05853_/X _05841_/X _05771_/A _05937_/X vssd1 vssd1 vccd1 vccd1
+ _05938_/X sky130_fd_sc_hd__o221a_1
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ _08686_/A _08659_/A vssd1 vssd1 vccd1 vccd1 _08778_/A sky130_fd_sc_hd__and2_2
X_05869_ _08000_/A _05872_/A vssd1 vssd1 vccd1 vccd1 _05869_/Y sky130_fd_sc_hd__nand2_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07608_ _07615_/A _06962_/X _07624_/A vssd1 vssd1 vccd1 vccd1 _07609_/B sky130_fd_sc_hd__a21oi_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _10782_/Q _08586_/B _08583_/A vssd1 vssd1 vccd1 vccd1 _08588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ _07539_/A _07607_/A vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__and2_1
XFILLER_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06088__A1 _05778_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06088__B2 _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _10554_/CLK _10550_/D vssd1 vssd1 vccd1 vccd1 _10550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09209_ _09037_/A _09209_/B vssd1 vssd1 vccd1 vccd1 _09274_/A sky130_fd_sc_hd__and2b_2
X_10481_ _06008_/X _10475_/X _10480_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10964_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08314__A input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08537__B1 _08462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06769__A _06769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06012__A1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10657_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05523__B1 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10847_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10817_ _10821_/CLK _10817_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06079__A1 _06113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06079__B2 _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07112__B _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10748_ _10784_/CLK _10748_/D vssd1 vssd1 vccd1 vccd1 _10748_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06009__A _10579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05826__A1 _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10679_ _10703_/CLK _10679_/D vssd1 vssd1 vccd1 vccd1 _10679_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_13_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10790_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06910_ _10502_/A _07776_/B _07783_/B _07780_/C vssd1 vssd1 vccd1 vccd1 _06910_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07890_ _10604_/Q _07888_/X _07874_/X _07889_/Y vssd1 vssd1 vccd1 vccd1 _07891_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_96_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06841_ _06841_/A vssd1 vssd1 vccd1 vccd1 _10513_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_96_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_28_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10958_/CLK sky130_fd_sc_hd__clkbuf_16
X_09560_ _09560_/A _09560_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__xnor2_1
X_06772_ _06772_/A _06772_/B vssd1 vssd1 vccd1 vccd1 _06773_/C sky130_fd_sc_hd__xnor2_1
XFILLER_167_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08511_ _10792_/Q _08506_/X _08509_/X _10755_/Q vssd1 vssd1 vccd1 vccd1 _10755_/D
+ sky130_fd_sc_hd__a22o_1
X_05723_ _05721_/Y _10542_/Q _10541_/Q _05736_/A vssd1 vssd1 vccd1 vccd1 _05732_/B
+ sky130_fd_sc_hd__a22o_1
X_09491_ _09618_/A _09491_/B vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08442_ _10769_/Q _10732_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08443_/B sky130_fd_sc_hd__mux2_1
XFILLER_169_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05654_ _10684_/Q _05637_/Y _05649_/X _05718_/A _05653_/X vssd1 vssd1 vccd1 vccd1
+ _05654_/X sky130_fd_sc_hd__o221a_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08373_ _08367_/X _10730_/Q _07865_/X _08372_/X vssd1 vssd1 vccd1 vccd1 _10712_/D
+ sky130_fd_sc_hd__o211a_1
X_05585_ _08315_/A vssd1 vssd1 vccd1 vccd1 _05803_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07324_ _07324_/A _07324_/B vssd1 vssd1 vccd1 vccd1 _07338_/B sky130_fd_sc_hd__and2_1
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07255_ _07258_/A _07258_/B _07214_/A vssd1 vssd1 vccd1 vccd1 _07256_/B sky130_fd_sc_hd__o21a_1
X_06206_ input22/X vssd1 vssd1 vccd1 vccd1 _06206_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_164_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07186_ _07186_/A _07186_/B _07186_/C vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__and3_1
XFILLER_117_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08767__B1 _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06137_ _10529_/A vssd1 vssd1 vccd1 vccd1 _06137_/X sky130_fd_sc_hd__buf_2
XFILLER_145_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07973__A _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06068_ _05693_/A _07981_/A _06065_/X _06066_/Y _06067_/X vssd1 vssd1 vccd1 vccd1
+ _06069_/D sky130_fd_sc_hd__o221a_1
XFILLER_160_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08519__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09827_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__and2_1
XFILLER_19_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09758_ _09755_/X _09757_/X _10875_/Q _09406_/X vssd1 vssd1 vccd1 vccd1 _10875_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08709_ _08709_/A _08725_/A vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__nor2_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09689_ _09689_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09755_/A sky130_fd_sc_hd__or2b_1
XFILLER_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10602_ _10814_/CLK _10602_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10533_ _10533_/A _10537_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10533_/X sky130_fd_sc_hd__or3_1
XFILLER_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10464_ _06187_/X _10459_/X _10463_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10958_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10395_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_leaf_26_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05370_ _10660_/Q vssd1 vssd1 vccd1 vccd1 _07985_/A sky130_fd_sc_hd__clkinv_2
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10484__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07040_ _07416_/A _07433_/A _07434_/A _07567_/A vssd1 vssd1 vccd1 vccd1 _07041_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_146_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06224__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08991_ _10799_/Q _08985_/X _08988_/X _10712_/Q _08990_/X vssd1 vssd1 vccd1 vccd1
+ _08991_/X sky130_fd_sc_hd__a221o_1
XFILLER_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07942_ _07955_/A _07942_/B vssd1 vssd1 vccd1 vccd1 _07943_/A sky130_fd_sc_hd__or2_1
XFILLER_69_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07873_ _07880_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _10631_/D sky130_fd_sc_hd__nor2_1
XANTENNA__06202__A input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09612_ _09613_/A _09613_/B _09613_/C vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__o21ai_2
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06824_ _06824_/A _06824_/B vssd1 vssd1 vccd1 vccd1 _06875_/A sky130_fd_sc_hd__or2_1
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09543_ _09618_/B _09543_/B vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06755_ _06755_/A _06755_/B vssd1 vssd1 vccd1 vccd1 _06806_/B sky130_fd_sc_hd__xnor2_4
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05706_ _05877_/A vssd1 vssd1 vccd1 vccd1 _08196_/A sky130_fd_sc_hd__inv_2
X_09474_ _09475_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__or2_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06686_ _06686_/A _06686_/B vssd1 vssd1 vccd1 vccd1 _06941_/A sky130_fd_sc_hd__xnor2_1
XFILLER_169_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08425_ _08624_/B vssd1 vssd1 vccd1 vccd1 _08661_/A sky130_fd_sc_hd__buf_2
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05637_ _10545_/Q _05637_/B vssd1 vssd1 vccd1 vccd1 _05637_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08356_ _08348_/Y _08086_/X _08157_/A _08354_/X _08355_/X vssd1 vssd1 vccd1 vccd1
+ _08357_/B sky130_fd_sc_hd__o221a_1
X_05568_ _08351_/A vssd1 vssd1 vccd1 vccd1 _08350_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07307_ _07307_/A _07307_/B vssd1 vssd1 vccd1 vccd1 _07347_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08287_ _08287_/A _08295_/C vssd1 vssd1 vccd1 vccd1 _08287_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10394__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05499_ _05374_/X _05497_/X _05490_/A _05461_/A vssd1 vssd1 vccd1 vccd1 _10552_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07238_ _07211_/A _07125_/A _07244_/B _07237_/X vssd1 vssd1 vccd1 vccd1 _07264_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_153_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07169_ _07169_/A _07169_/B vssd1 vssd1 vccd1 vccd1 _07184_/B sky130_fd_sc_hd__nand2_1
XFILLER_161_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06215__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10180_ _07013_/A _10174_/X _10177_/X _10891_/Q vssd1 vssd1 vccd1 vccd1 _10891_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09142__B _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10516_ _06168_/X _10497_/B _10515_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10978_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10447_ _10472_/B vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10378_ _10365_/X _10713_/Q _10375_/X _10377_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10932_/D sky130_fd_sc_hd__o221a_1
XANTENNA__08502__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07954__A1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06540_ _06540_/A vssd1 vssd1 vccd1 vccd1 _06719_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06471_ _06474_/A _06474_/B vssd1 vssd1 vccd1 vccd1 _06666_/B sky130_fd_sc_hd__or2_1
X_08210_ _08218_/B _08061_/A _08208_/Y _08209_/Y _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08210_/X sky130_fd_sc_hd__a311o_1
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05422_ _10628_/Q _05371_/Y _05374_/X _05461_/A _05421_/X vssd1 vssd1 vccd1 vccd1
+ _05422_/X sky130_fd_sc_hd__o221a_1
X_09190_ _08198_/A _09226_/S _09203_/A _09189_/X vssd1 vssd1 vccd1 vccd1 _09190_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_140_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08141_ _08058_/A _08137_/Y _08140_/Y _08113_/A _08096_/A vssd1 vssd1 vccd1 vccd1
+ _08141_/X sky130_fd_sc_hd__a221o_1
X_05353_ _05353_/A _05353_/B vssd1 vssd1 vccd1 vccd1 _05353_/X sky130_fd_sc_hd__and2_1
XFILLER_174_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08072_ _08075_/A _08072_/B vssd1 vssd1 vccd1 vccd1 _08072_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_135_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05284_ _10650_/Q _10574_/Q vssd1 vssd1 vccd1 vccd1 _05401_/A sky130_fd_sc_hd__xor2_1
XFILLER_162_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07023_ _07222_/A vssd1 vssd1 vccd1 vccd1 _07169_/A sky130_fd_sc_hd__buf_2
XFILLER_128_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08974_ _08974_/A vssd1 vssd1 vccd1 vccd1 _08974_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07925_ _07925_/A vssd1 vssd1 vccd1 vccd1 _07925_/Y sky130_fd_sc_hd__inv_2
XFILLER_60_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07856_ _10877_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09243__A _09274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06807_ _06818_/A _06817_/B vssd1 vssd1 vccd1 vccd1 _06853_/A sky130_fd_sc_hd__or2_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07787_ _07787_/A _07787_/B vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09526_ _09625_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__xnor2_1
X_06738_ _06752_/A _06738_/B vssd1 vssd1 vccd1 vccd1 _06758_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__08122__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _09456_/B _09456_/C _09456_/A vssd1 vssd1 vccd1 vccd1 _09458_/C sky130_fd_sc_hd__a21o_1
XFILLER_52_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06669_ _06686_/A _06686_/B vssd1 vssd1 vccd1 vccd1 _06915_/B sky130_fd_sc_hd__and2_1
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08408_ _08408_/A _10760_/Q vssd1 vssd1 vccd1 vccd1 _08408_/X sky130_fd_sc_hd__or2_1
X_09388_ _09388_/A _09388_/B vssd1 vssd1 vccd1 vccd1 _09411_/A sky130_fd_sc_hd__xnor2_2
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08339_ _08339_/A _08339_/B _08339_/C vssd1 vssd1 vccd1 vccd1 _08350_/B sky130_fd_sc_hd__and3_1
XANTENNA__08306__B _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10301_ _10301_/A _10301_/B vssd1 vssd1 vccd1 vccd1 _10301_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10232_ _07056_/A _10115_/X _10231_/X _10043_/X vssd1 vssd1 vccd1 vccd1 _10902_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10163_ _10112_/A _10112_/B _10162_/X vssd1 vssd1 vccd1 vccd1 _10164_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09138__B1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input37_A io_wbs_m2s_data[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _10097_/A _10025_/B vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__or2b_1
XFILLER_121_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08361__A1 _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09153__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08992__A _08992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10189__A_N _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07872__B1 _07848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08821__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05971_ _08965_/A _09124_/B vssd1 vssd1 vccd1 vccd1 _09107_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07710_ _07607_/A _07604_/B _07539_/A vssd1 vssd1 vccd1 vccd1 _07758_/A sky130_fd_sc_hd__o21ai_2
X_08690_ _10802_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08691_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07641_ _07641_/A _07641_/B vssd1 vssd1 vccd1 vccd1 _07693_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07572_ _09379_/B _07572_/B vssd1 vssd1 vccd1 vccd1 _07574_/B sky130_fd_sc_hd__xnor2_1
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10002__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09311_ _10043_/A _09309_/Y _09326_/A _10192_/A _10866_/Q vssd1 vssd1 vccd1 vccd1
+ _10866_/D sky130_fd_sc_hd__a32o_1
X_06523_ _06532_/A _06523_/B _06523_/C vssd1 vssd1 vccd1 vccd1 _06545_/A sky130_fd_sc_hd__and3_1
XFILLER_22_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09242_ _09242_/A vssd1 vssd1 vccd1 vccd1 _10855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06454_ _06477_/A _06477_/B vssd1 vssd1 vccd1 vccd1 _06478_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08407__A _09090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05405_ _05405_/A _05643_/A vssd1 vssd1 vccd1 vccd1 _05406_/B sky130_fd_sc_hd__nor2_1
X_09173_ _09112_/X _09167_/Y _09172_/X vssd1 vssd1 vccd1 vccd1 _09174_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06385_ _06305_/A _06274_/B _06374_/B _06303_/A vssd1 vssd1 vccd1 vccd1 _06386_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_159_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08124_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08124_/X sky130_fd_sc_hd__clkbuf_2
X_05336_ _05336_/A _05336_/B vssd1 vssd1 vccd1 vccd1 _05337_/B sky130_fd_sc_hd__and2_1
XANTENNA__07030__B _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ _06124_/A _08047_/X _08052_/X _08082_/D _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08055_/X sky130_fd_sc_hd__o221a_1
XFILLER_119_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07006_ _07197_/A vssd1 vssd1 vccd1 vccd1 _07567_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07981__A _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08957_ _09610_/B vssd1 vssd1 vccd1 vccd1 _09867_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_76_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07908_ _10609_/Q _07906_/X _07892_/X _07907_/Y vssd1 vssd1 vccd1 vccd1 _07909_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08888_ _10825_/Q _08888_/B vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__or2_1
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07839_ _06170_/A _07828_/X _07829_/X _07838_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07839_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10150__A1 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _10850_/CLK _10850_/D vssd1 vssd1 vccd1 vccd1 _10850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09509_ _09867_/A _09610_/B _09555_/B _09599_/B vssd1 vssd1 vccd1 vccd1 _09613_/A
+ sky130_fd_sc_hd__and4_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ _10782_/CLK _10781_/D vssd1 vssd1 vccd1 vccd1 _10781_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08317__A _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07082__A1 _09356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08052__A _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10215_ _10226_/B _10226_/C vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__nand2_1
XFILLER_122_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10146_ _10146_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10429__C1 _06257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10979_ _10984_/CLK _10979_/D vssd1 vssd1 vccd1 vccd1 _10979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06170_ _06170_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06170_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06970__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_74_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09860_ _09735_/A _09735_/B _09859_/Y _09432_/A vssd1 vssd1 vccd1 vccd1 _09864_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _10815_/Q vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__clkbuf_2
X_09791_ _09711_/B _09727_/B _09711_/A vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__o21bai_4
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10380__A1 _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08742_ _08744_/B vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__buf_2
X_05954_ _05954_/A vssd1 vssd1 vccd1 vccd1 _05954_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_66_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08673_ _08686_/A _08830_/A vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10132__A1 _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05885_ _05885_/A vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__buf_2
XFILLER_93_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07624_ _07624_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _07625_/B sky130_fd_sc_hd__nor2_2
XFILLER_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07555_ _07732_/A _07555_/B _07713_/B vssd1 vssd1 vccd1 vccd1 _07556_/B sky130_fd_sc_hd__and3_1
XANTENNA__08089__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06506_ _06517_/A _06506_/B vssd1 vssd1 vccd1 vccd1 _06507_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07486_ _07485_/A _07485_/B _07493_/B _07493_/A vssd1 vssd1 vccd1 vccd1 _07495_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_139_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09225_ _08242_/A _07885_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09225_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06437_ _10975_/Q _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06472_/A sky130_fd_sc_hd__and3_1
XFILLER_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09156_ _10942_/Q _09143_/Y _09155_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09156_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07976__A _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06368_ _06451_/C _06368_/B vssd1 vssd1 vccd1 vccd1 _06895_/B sky130_fd_sc_hd__nor2_2
XFILLER_108_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08107_ _08113_/A _08104_/Y _08115_/B _06024_/A vssd1 vssd1 vccd1 vccd1 _08107_/X
+ sky130_fd_sc_hd__a31o_1
X_05319_ _10646_/Q vssd1 vssd1 vccd1 vccd1 _07925_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09087_ _10513_/A _09086_/X _09087_/S vssd1 vssd1 vccd1 vccd1 _09087_/X sky130_fd_sc_hd__mux2_1
X_06299_ _10920_/Q _10903_/Q vssd1 vssd1 vccd1 vccd1 _06304_/B sky130_fd_sc_hd__or2_1
X_08038_ _08038_/A vssd1 vssd1 vccd1 vccd1 _08038_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10000_ _09801_/A _09933_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _10001_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09989_ _09989_/A _09989_/B vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__xnor2_1
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10902_ _10926_/CLK _10902_/D vssd1 vssd1 vccd1 vccd1 _10902_/Q sky130_fd_sc_hd__dfxtp_2
X_10833_ _10833_/CLK _10833_/D vssd1 vssd1 vccd1 vccd1 _10833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10426__A2 _10726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10764_ _10833_/CLK _10764_/D vssd1 vssd1 vccd1 vccd1 _10764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08047__A _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10695_ _10851_/CLK _10695_/D vssd1 vssd1 vccd1 vccd1 _10695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08252__B1 _05598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06014__B input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10362__A1 _08491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10129_ _10129_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10251__S _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06030__A2 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07126__A _10985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10114__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05670_ _08224_/B _05610_/X _05606_/X _10697_/Q _05669_/X vssd1 vssd1 vccd1 vccd1
+ _05670_/X sky130_fd_sc_hd__o221a_1
XFILLER_91_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10487__A _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07340_ _07525_/A _07525_/B _07526_/A vssd1 vssd1 vccd1 vccd1 _07528_/C sky130_fd_sc_hd__a21o_1
XFILLER_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07271_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07335_/A sky130_fd_sc_hd__or2_1
X_09010_ _09124_/A vssd1 vssd1 vccd1 vccd1 _09194_/B sky130_fd_sc_hd__clkbuf_2
X_06222_ input25/X _06207_/X _06220_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10602_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06153_ _10343_/A vssd1 vssd1 vccd1 vccd1 _06153_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__06254__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08794__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06084_ _05291_/A _08093_/A _05766_/Y _05830_/A vssd1 vssd1 vccd1 vccd1 _06089_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09912_ _09842_/A _09842_/B _09841_/A vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__a21oi_2
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09843_ _09843_/A _09775_/A vssd1 vssd1 vccd1 vccd1 _09844_/C sky130_fd_sc_hd__or2b_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09771_/B _09773_/X _09705_/B _09708_/A vssd1 vssd1 vccd1 vccd1 _09843_/A
+ sky130_fd_sc_hd__o31a_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _06997_/B _06986_/B vssd1 vssd1 vccd1 vccd1 _07020_/B sky130_fd_sc_hd__xnor2_1
XFILLER_74_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05937_ _08277_/A _05935_/B _05853_/X _08285_/A _05936_/X vssd1 vssd1 vccd1 vccd1
+ _05937_/X sky130_fd_sc_hd__a221o_1
X_08725_ _08725_/A _08725_/B vssd1 vssd1 vccd1 vccd1 _08740_/B sky130_fd_sc_hd__and2_1
XFILLER_73_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _10369_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _08659_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05868_ _10665_/Q vssd1 vssd1 vccd1 vccd1 _08000_/A sky130_fd_sc_hd__buf_2
XFILLER_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07607_ _07607_/A _07607_/B vssd1 vssd1 vccd1 vccd1 _07610_/A sky130_fd_sc_hd__nand2_2
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _10781_/Q _08583_/B _08586_/Y vssd1 vssd1 vccd1 vccd1 _10781_/D sky130_fd_sc_hd__o21a_1
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05799_ _05717_/B _05798_/Y _05708_/A vssd1 vssd1 vccd1 vccd1 _05799_/X sky130_fd_sc_hd__o21a_1
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07538_ _07606_/A _07606_/B vssd1 vssd1 vccd1 vccd1 _07607_/A sky130_fd_sc_hd__or2_1
XFILLER_41_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06088__A2 _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07469_ _07746_/A _07469_/B vssd1 vssd1 vccd1 vccd1 _07497_/A sky130_fd_sc_hd__xor2_1
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09208_ _09208_/A vssd1 vssd1 vccd1 vccd1 _10850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10480_ _10480_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10480_/X sky130_fd_sc_hd__or2_1
XFILLER_148_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09139_ _10808_/Q _08985_/X _08988_/X _10721_/Q _09138_/X vssd1 vssd1 vccd1 vccd1
+ _09139_/X sky130_fd_sc_hd__a221o_1
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06115__A _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05954__A _05954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_9_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10798_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10816_ _10822_/CLK _10816_/D vssd1 vssd1 vccd1 vccd1 _10816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08068__A3 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06079__A2 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10747_ _10784_/CLK _10747_/D vssd1 vssd1 vccd1 vccd1 _10747_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10678_ _10859_/CLK _10678_/D vssd1 vssd1 vccd1 vccd1 _10678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06840_ _07789_/A _06840_/B vssd1 vssd1 vccd1 vccd1 _06864_/A sky130_fd_sc_hd__and2_1
XFILLER_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06771_ _06940_/A _06771_/B vssd1 vssd1 vccd1 vccd1 _06772_/B sky130_fd_sc_hd__nand2_1
X_08510_ _10791_/Q _08506_/X _08509_/X _10754_/Q vssd1 vssd1 vccd1 vccd1 _10754_/D
+ sky130_fd_sc_hd__a22o_1
X_05722_ _05913_/A vssd1 vssd1 vccd1 vccd1 _05736_/A sky130_fd_sc_hd__buf_4
X_09490_ _09489_/A _09642_/A _09492_/A _09555_/A vssd1 vssd1 vccd1 vccd1 _09491_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__08161__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08441_ _08476_/S vssd1 vssd1 vccd1 vccd1 _08455_/S sky130_fd_sc_hd__clkbuf_2
X_05653_ _05651_/Y _05652_/X _05649_/X _05718_/A vssd1 vssd1 vccd1 vccd1 _05653_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08372_ _08381_/A _10746_/Q vssd1 vssd1 vccd1 vccd1 _08372_/X sky130_fd_sc_hd__or2_1
X_05584_ _10706_/Q vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__buf_2
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07323_ _07323_/A _07323_/B _07331_/A vssd1 vssd1 vccd1 vccd1 _07324_/B sky130_fd_sc_hd__nand3_1
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07254_ _07254_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07258_/B sky130_fd_sc_hd__and2_1
XANTENNA__05817__A2 _09078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08415__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06205_ _06202_/X _06183_/X _06204_/Y _06200_/X vssd1 vssd1 vccd1 vccd1 _10598_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07185_ _07185_/A _07185_/B vssd1 vssd1 vccd1 vccd1 _07201_/A sky130_fd_sc_hd__xnor2_1
XFILLER_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06136_ _08166_/A vssd1 vssd1 vccd1 vccd1 _10529_/A sky130_fd_sc_hd__buf_4
XFILLER_132_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07975__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06067_ _05756_/A _08235_/A _05818_/A _08082_/A vssd1 vssd1 vccd1 vccd1 _06067_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_59_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08150__A _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09826_ _09815_/A _09815_/B _09825_/X vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__a21o_1
XFILLER_87_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09757_ _09757_/A _09757_/B vssd1 vssd1 vccd1 vccd1 _09757_/X sky130_fd_sc_hd__or2_1
X_06969_ _07007_/A vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__buf_2
XFILLER_73_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _10804_/Q _08732_/B vssd1 vssd1 vccd1 vccd1 _08725_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _10043_/A _09686_/X _09755_/B _10192_/A _10874_/Q vssd1 vssd1 vccd1 vccd1
+ _10874_/D sky130_fd_sc_hd__a32o_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _08638_/B _10793_/Q _08600_/A _08642_/D _10795_/Q vssd1 vssd1 vccd1 vccd1
+ _08640_/B sky130_fd_sc_hd__a41o_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10601_ _10814_/CLK _10601_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10532_ _07713_/A _10522_/X _10531_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10983_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_128_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10463_ _10958_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10463_/X sky130_fd_sc_hd__or2_1
XFILLER_10_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10394_ _10535_/A _10394_/B _10394_/C vssd1 vssd1 vccd1 vccd1 _10394_/X sky130_fd_sc_hd__and3_1
XFILLER_136_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05441__B1 _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08060__A _08352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09603__B _09610_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08997__A1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08235__A _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08749__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ _10765_/Q _09037_/A _08990_/C vssd1 vssd1 vccd1 vccd1 _08990_/X sky130_fd_sc_hd__and3_1
XFILLER_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07941_ input27/X _05813_/A _07964_/A vssd1 vssd1 vccd1 vccd1 _07942_/B sky130_fd_sc_hd__mux2_1
XFILLER_69_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07872_ _10599_/Q _07870_/X _07848_/A _07871_/Y vssd1 vssd1 vccd1 vccd1 _07873_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09611_ _09611_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09613_/C sky130_fd_sc_hd__nor2_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06823_ _06823_/A _06823_/B vssd1 vssd1 vccd1 vccd1 _06824_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05735__B2 _05733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09542_ _09542_/A _09542_/B _09542_/C vssd1 vssd1 vccd1 vccd1 _09543_/B sky130_fd_sc_hd__and3_1
X_06754_ _06317_/B _06729_/B _06317_/A vssd1 vssd1 vccd1 vccd1 _06755_/B sky130_fd_sc_hd__a21bo_1
XFILLER_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05705_ _05704_/Y _05663_/A _10553_/Q _08181_/A vssd1 vssd1 vccd1 vccd1 _05708_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09473_ _09524_/A _09473_/B vssd1 vssd1 vccd1 vccd1 _09475_/B sky130_fd_sc_hd__xnor2_1
X_06685_ _06943_/B _06943_/C _06943_/A vssd1 vssd1 vccd1 vccd1 _06944_/A sky130_fd_sc_hd__a21o_1
XANTENNA__05499__B1 _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08424_ _08424_/A _08424_/B vssd1 vssd1 vccd1 vccd1 _08624_/B sky130_fd_sc_hd__xnor2_4
X_05636_ _05636_/A _05636_/B vssd1 vssd1 vccd1 vccd1 _05636_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08355_/X sky130_fd_sc_hd__or2_1
XFILLER_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05567_ _10710_/Q vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__buf_2
X_07306_ _07349_/B _07349_/C _07349_/A vssd1 vssd1 vccd1 vccd1 _07461_/B sky130_fd_sc_hd__o21a_1
XFILLER_165_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08286_ _08287_/A _08295_/C vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__and2_1
X_05498_ _05378_/Y _05497_/X _05490_/X _05461_/B vssd1 vssd1 vccd1 vccd1 _10551_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_137_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07237_ _07236_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07237_/X sky130_fd_sc_hd__and2b_1
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07984__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07168_ _07196_/A _07334_/A _07195_/A vssd1 vssd1 vccd1 vccd1 _07192_/B sky130_fd_sc_hd__a21o_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06119_ _07880_/A _06119_/B vssd1 vssd1 vccd1 vccd1 _10582_/D sky130_fd_sc_hd__nor2_1
X_07099_ _07219_/B vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_74_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10857_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09809_ _09883_/A _09809_/B vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__xor2_2
XFILLER_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10788_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_27_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10940_/CLK sky130_fd_sc_hd__clkbuf_16
X_10515_ _10515_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10515_/X sky130_fd_sc_hd__or2_1
XFILLER_156_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10446_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10446_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10538__A1 _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10377_ _06008_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10377_/X sky130_fd_sc_hd__a21bo_1
XFILLER_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06470_ _06470_/A _06470_/B vssd1 vssd1 vccd1 vccd1 _06474_/B sky130_fd_sc_hd__nor2_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05421_ _05461_/B _05378_/Y _05374_/X _10627_/Q _05420_/X vssd1 vssd1 vccd1 vccd1
+ _05421_/X sky130_fd_sc_hd__a221o_1
XFILLER_53_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10495__A _10495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08140_ _08148_/B _08140_/B vssd1 vssd1 vccd1 vccd1 _08140_/Y sky130_fd_sc_hd__nor2_1
X_05352_ _10666_/Q _05358_/A vssd1 vssd1 vccd1 vccd1 _05353_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08071_ _08082_/B vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05283_ _10574_/Q vssd1 vssd1 vccd1 vccd1 _05283_/Y sky130_fd_sc_hd__inv_2
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ _10980_/Q vssd1 vssd1 vccd1 vccd1 _07222_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08973_ _09211_/A vssd1 vssd1 vccd1 vccd1 _08974_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06213__A _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07924_ _08284_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _10645_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07855_ _07848_/X _05461_/B _07844_/X _07854_/Y vssd1 vssd1 vccd1 vccd1 _10626_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06806_ _06806_/A _06806_/B vssd1 vssd1 vccd1 vccd1 _06817_/B sky130_fd_sc_hd__or2_1
XFILLER_72_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07786_ _07786_/A _07786_/B vssd1 vssd1 vccd1 vccd1 _07787_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09525_ _09626_/A _09625_/B vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06737_ _06745_/B _06746_/A _07675_/A vssd1 vssd1 vccd1 vccd1 _06738_/B sky130_fd_sc_hd__a21o_1
XFILLER_64_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07979__A _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09456_ _09456_/A _09456_/B _09456_/C vssd1 vssd1 vccd1 vccd1 _09458_/B sky130_fd_sc_hd__nand3_1
XFILLER_25_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06668_ _06668_/A _06668_/B vssd1 vssd1 vccd1 vccd1 _06686_/B sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_69_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05619_ _05663_/B _05619_/B vssd1 vssd1 vccd1 vccd1 _05619_/X sky130_fd_sc_hd__and2_1
X_08407_ _09090_/A vssd1 vssd1 vccd1 vccd1 _08992_/A sky130_fd_sc_hd__buf_2
X_09387_ _09387_/A _09424_/A vssd1 vssd1 vccd1 vccd1 _09388_/B sky130_fd_sc_hd__nand2_1
X_06599_ _06599_/A _06599_/B vssd1 vssd1 vccd1 vccd1 _06616_/A sky130_fd_sc_hd__xnor2_1
XFILLER_8_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08338_ _06033_/X _08334_/X _08336_/Y _08337_/X vssd1 vssd1 vccd1 vccd1 _10708_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_137_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _08278_/B _08253_/X _08267_/Y _08268_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08269_/X sky130_fd_sc_hd__a311o_1
XFILLER_125_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10300_ _10300_/A _10300_/B vssd1 vssd1 vccd1 vccd1 _10301_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10231_ _10246_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__xor2_2
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10162_ _10110_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10162_/X sky130_fd_sc_hd__and2b_1
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06123__A input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09138__A1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10093_ _10121_/S _10093_/B vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__nor2_2
XFILLER_121_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05962__A input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09074__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10429_ _10408_/A _10727_/Q _10427_/X _10428_/X _06257_/X vssd1 vssd1 vccd1 vccd1
+ _10946_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06060__B1 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05970_ _06126_/D vssd1 vssd1 vccd1 vccd1 _09124_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_112_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08337__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07640_ _07645_/A _07644_/B _07662_/A vssd1 vssd1 vccd1 vccd1 _07641_/B sky130_fd_sc_hd__a21oi_1
XFILLER_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07571_ _07678_/A _07571_/B vssd1 vssd1 vccd1 vccd1 _07572_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09310_ _09313_/B _09396_/A _09310_/C vssd1 vssd1 vccd1 vccd1 _09326_/A sky130_fd_sc_hd__or3_1
X_06522_ _06600_/A _06522_/B _06522_/C vssd1 vssd1 vccd1 vccd1 _06602_/A sky130_fd_sc_hd__and3_1
XFILLER_62_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_70_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09241_ _09259_/A _09241_/B vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__and2_1
XFILLER_61_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06453_ _06453_/A _06453_/B vssd1 vssd1 vccd1 vccd1 _06477_/B sky130_fd_sc_hd__or2_1
XFILLER_166_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05404_ _10573_/Q vssd1 vssd1 vccd1 vccd1 _05643_/A sky130_fd_sc_hd__clkbuf_2
X_09172_ _08771_/A _09168_/X _09079_/X _10724_/Q _09171_/X vssd1 vssd1 vccd1 vccd1
+ _09172_/X sky130_fd_sc_hd__a221o_1
X_06384_ _06719_/A vssd1 vssd1 vccd1 vccd1 _10515_/A sky130_fd_sc_hd__buf_4
XFILLER_119_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08123_/X sky130_fd_sc_hd__clkbuf_2
X_05335_ _08298_/A _05340_/A vssd1 vssd1 vccd1 vccd1 _05336_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08054_ _08175_/A vssd1 vssd1 vccd1 vccd1 _08054_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07005_ _07188_/A vssd1 vssd1 vccd1 vccd1 _07197_/A sky130_fd_sc_hd__buf_2
XFILLER_162_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09368__B2 _09356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07039__A _07416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08040__A1 _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05929__A1 _05877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08956_ _09449_/A vssd1 vssd1 vccd1 vccd1 _09610_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07907_ _07907_/A vssd1 vssd1 vccd1 vccd1 _07907_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08887_ _10825_/Q _08902_/B vssd1 vssd1 vccd1 vccd1 _08889_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07838_ _10873_/Q _07845_/B vssd1 vssd1 vccd1 vccd1 _07838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07769_ _07769_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07771_/A sky130_fd_sc_hd__xnor2_1
XFILLER_112_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09508_ _09508_/A _09508_/B vssd1 vssd1 vccd1 vccd1 _09599_/B sky130_fd_sc_hd__xor2_4
XANTENNA__10438__B1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _10782_/CLK _10780_/D vssd1 vssd1 vccd1 vccd1 _10780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09439_ _09438_/A _09438_/B _10351_/A vssd1 vssd1 vccd1 vccd1 _09439_/X sky130_fd_sc_hd__o21a_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05957__A input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08031__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ _10214_/A vssd1 vssd1 vccd1 vccd1 _10226_/C sky130_fd_sc_hd__inv_2
XFILLER_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06042__B1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__05692__A _05692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10076_ _10076_/A _10001_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__or2b_1
XFILLER_48_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08334__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10978_ _10978_/CLK _10978_/D vssd1 vssd1 vccd1 vccd1 _10978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09339__A _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08022__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08810_ _08810_/A _08814_/A _08817_/B vssd1 vssd1 vccd1 vccd1 _08810_/X sky130_fd_sc_hd__or3b_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09790_ _09827_/A _09827_/B vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__xor2_4
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08741_ _10806_/Q _10805_/Q _10804_/Q _08701_/A _08744_/B vssd1 vssd1 vccd1 vccd1
+ _08741_/X sky130_fd_sc_hd__o41a_1
X_05953_ _06019_/A _10540_/Q vssd1 vssd1 vccd1 vccd1 _05954_/A sky130_fd_sc_hd__and2_4
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08325__A2 _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ _08830_/A vssd1 vssd1 vccd1 vccd1 _08672_/X sky130_fd_sc_hd__clkbuf_2
X_05884_ _07988_/A _05883_/X _05878_/B vssd1 vssd1 vccd1 vccd1 _05884_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_94_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07623_ _07623_/A _07623_/B vssd1 vssd1 vccd1 vccd1 _07700_/A sky130_fd_sc_hd__xor2_4
XANTENNA__09286__A0 _08339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08089__A1 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07554_ _07426_/A _07425_/B _07425_/A vssd1 vssd1 vccd1 vccd1 _07556_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__08089__B2 _05733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06505_ _06521_/A _06517_/C _06503_/Y _06517_/B _06758_/A vssd1 vssd1 vccd1 vccd1
+ _06519_/A sky130_fd_sc_hd__o2111a_1
X_07485_ _07485_/A _07485_/B vssd1 vssd1 vccd1 vccd1 _07493_/B sky130_fd_sc_hd__xnor2_1
XFILLER_139_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09224_ _09224_/A vssd1 vssd1 vccd1 vccd1 _10852_/D sky130_fd_sc_hd__buf_4
X_06436_ _06436_/A _06456_/A _07682_/B _06460_/B vssd1 vssd1 vccd1 vccd1 _06468_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_148_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06367_ _06367_/A _06917_/A vssd1 vssd1 vccd1 vccd1 _06368_/B sky130_fd_sc_hd__nand2_1
X_09155_ _10958_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05318_ _05318_/A _05318_/B vssd1 vssd1 vccd1 vccd1 _05318_/X sky130_fd_sc_hd__and2_1
X_08106_ _08116_/B vssd1 vssd1 vccd1 vccd1 _08115_/B sky130_fd_sc_hd__inv_2
XFILLER_163_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09249__A _09249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06298_ _10920_/Q _10903_/Q vssd1 vssd1 vccd1 vccd1 _06304_/A sky130_fd_sc_hd__nand2_1
X_09086_ _10491_/A _09085_/X _09086_/S vssd1 vssd1 vccd1 vccd1 _09086_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08037_ _08037_/A vssd1 vssd1 vccd1 vccd1 _08038_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07992__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _10065_/C _10065_/B vssd1 vssd1 vccd1 vccd1 _09989_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08939_ input6/X input5/X _08939_/C input15/X vssd1 vssd1 vccd1 vccd1 _09142_/D sky130_fd_sc_hd__or4b_4
XFILLER_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10901_ _10980_/CLK _10901_/D vssd1 vssd1 vccd1 vccd1 _10901_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_45_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10832_ _10833_/CLK _10832_/D vssd1 vssd1 vccd1 vccd1 _10832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ _10770_/CLK _10763_/D vssd1 vssd1 vccd1 vccd1 _10763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10694_ _10851_/CLK _10694_/D vssd1 vssd1 vccd1 vccd1 _10694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07055__A2 _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08004__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10128_ _10075_/A _10074_/A _10074_/B _10085_/A vssd1 vssd1 vccd1 vccd1 _10146_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08307__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10059_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09268__A0 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07270_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07334_/B sky130_fd_sc_hd__or2_1
X_06221_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06221_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06152_ _08166_/A vssd1 vssd1 vccd1 vccd1 _10343_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06083_ _05766_/Y _05830_/A _07976_/A _05711_/Y vssd1 vssd1 vccd1 vccd1 _06089_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09911_ _09911_/A _09911_/B vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__nand2_1
XFILLER_99_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09842_ _09842_/A _09842_/B vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__xnor2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09773_/X sky130_fd_sc_hd__and2_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _07007_/A _06997_/C vssd1 vssd1 vccd1 vccd1 _06986_/B sky130_fd_sc_hd__nand2_1
XFILLER_101_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08724_ _10804_/Q _08701_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08724_/X sky130_fd_sc_hd__o21a_1
XFILLER_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05936_ _08277_/B _05858_/Y _05860_/X _05934_/X _05935_/X vssd1 vssd1 vccd1 vccd1
+ _05936_/X sky130_fd_sc_hd__o221a_1
XFILLER_113_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08655_ _08971_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__and2_1
X_05867_ _08233_/A _05866_/X _05863_/X _10699_/Q vssd1 vssd1 vccd1 vccd1 _05867_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ _07606_/A _07606_/B vssd1 vssd1 vccd1 vccd1 _07607_/B sky130_fd_sc_hd__nand2_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08586_ _08586_/A _08586_/B vssd1 vssd1 vccd1 vccd1 _08586_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05798_ _05798_/A _05798_/B vssd1 vssd1 vccd1 vccd1 _05798_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07537_ _07505_/X _07536_/X _07622_/A vssd1 vssd1 vccd1 vccd1 _07606_/B sky130_fd_sc_hd__o21a_1
XFILLER_23_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07987__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08482__A1 _10744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07501_/A sky130_fd_sc_hd__or2b_1
XFILLER_139_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09207_ _09228_/A _09207_/B vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__and2_4
X_06419_ _06386_/A _06386_/B _06418_/Y vssd1 vssd1 vccd1 vccd1 _06420_/B sky130_fd_sc_hd__o21a_1
XFILLER_148_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07399_ _07377_/A _07587_/B _07398_/B _07560_/A vssd1 vssd1 vccd1 vccd1 _07399_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09138_ _07976_/A _09123_/X _09127_/X _09137_/X vssd1 vssd1 vccd1 vccd1 _09138_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09069_ _09639_/B vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08537__A2 _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input12_A io_wbs_m2s_addr[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08058__A _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _10821_/CLK _10815_/D vssd1 vssd1 vccd1 vccd1 _10815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10746_ _10784_/CLK _10746_/D vssd1 vssd1 vccd1 vccd1 _10746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10677_ _10859_/CLK _10677_/D vssd1 vssd1 vccd1 vccd1 _10677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output80_A _10865_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06770_ _07682_/A _06842_/A vssd1 vssd1 vccd1 vccd1 _06940_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05721_ _08082_/C vssd1 vssd1 vccd1 vccd1 _05721_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10498__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08440_ _08440_/A vssd1 vssd1 vccd1 vccd1 _10731_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05652_ _05652_/A _05652_/B _05652_/C vssd1 vssd1 vccd1 vccd1 _05652_/X sky130_fd_sc_hd__or3_1
X_05583_ _05681_/B _05583_/B vssd1 vssd1 vccd1 vccd1 _05583_/Y sky130_fd_sc_hd__nor2_1
XFILLER_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08371_ _08547_/A vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07322_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07338_/A sky130_fd_sc_hd__nor2_1
XFILLER_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07253_ _07264_/B _07514_/A _07264_/A vssd1 vssd1 vccd1 vccd1 _07254_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08415__B input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06204_ _06204_/A _06204_/B vssd1 vssd1 vccd1 vccd1 _06204_/Y sky130_fd_sc_hd__nand2_1
X_07184_ _07184_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07185_/B sky130_fd_sc_hd__nor2_1
XFILLER_129_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06135_ _09403_/A vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_172_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09527__A _09527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06066_ _08082_/B vssd1 vssd1 vccd1 vccd1 _06066_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input4_A io_wbs_m2s_addr[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _09814_/B _09825_/B vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__and2b_1
XFILLER_24_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09756_ _09755_/A _09755_/B _09755_/C vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__a21oi_1
XFILLER_100_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06968_ _09381_/A vssd1 vssd1 vccd1 vccd1 _07007_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08707_ _08705_/X _08706_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10803_/D sky130_fd_sc_hd__a21oi_1
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05919_ _08095_/A _05906_/X _05904_/Y _06037_/A _05918_/X vssd1 vssd1 vccd1 vccd1
+ _05919_/X sky130_fd_sc_hd__a221o_1
XFILLER_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09687_ _09686_/A _09686_/B _09686_/C vssd1 vssd1 vccd1 vccd1 _09755_/B sky130_fd_sc_hd__o21ai_1
XFILLER_55_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06899_ _06899_/A _06899_/B vssd1 vssd1 vccd1 vccd1 _06928_/A sky130_fd_sc_hd__xnor2_4
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _10795_/Q _08638_/B _08638_/C vssd1 vssd1 vccd1 vccd1 _08638_/X sky130_fd_sc_hd__and3_1
XFILLER_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08569_ _08572_/B _08565_/X _08583_/A vssd1 vssd1 vccd1 vccd1 _08569_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10600_ _10814_/CLK _10600_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10262__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ _10531_/A _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10531_/X sky130_fd_sc_hd__or3_1
XFILLER_155_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10462_ _06182_/X _10459_/X _10461_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10957_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06126__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10393_ _10389_/X _10717_/Q _10390_/X _10391_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10936_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05965__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10729_ _10807_/CLK _10729_/D vssd1 vssd1 vccd1 vccd1 _10729_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08235__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07940_ _08445_/A vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07871_ _07871_/A vssd1 vssd1 vccd1 vccd1 _07871_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09610_ _09610_/A _09610_/B _09610_/C _09717_/A vssd1 vssd1 vccd1 vccd1 _09611_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06822_ _06823_/A _06823_/B vssd1 vssd1 vccd1 vccd1 _06824_/A sky130_fd_sc_hd__and2_1
XFILLER_96_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09082__A _10969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ _09542_/A _09542_/B _09542_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__a21oi_1
XFILLER_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06753_ _06804_/A _06806_/A vssd1 vssd1 vccd1 vccd1 _06756_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05704_ _08188_/A vssd1 vssd1 vccd1 vccd1 _05704_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09472_ _10066_/A _09472_/B vssd1 vssd1 vccd1 vccd1 _09473_/B sky130_fd_sc_hd__nor2_1
X_06684_ _06684_/A _06684_/B vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__xnor2_1
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08423_ _10833_/Q _10832_/Q vssd1 vssd1 vccd1 vccd1 _08424_/B sky130_fd_sc_hd__xor2_2
XFILLER_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10492__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05635_ _10546_/Q _05635_/B vssd1 vssd1 vccd1 vccd1 _05636_/B sky130_fd_sc_hd__and2_1
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08354_ _08263_/A _08349_/X _08350_/Y _08353_/X _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08354_/X sky130_fd_sc_hd__o32a_1
X_05566_ _05566_/A _05566_/B vssd1 vssd1 vccd1 vccd1 _05687_/B sky130_fd_sc_hd__and2_1
X_07305_ _07305_/A _07305_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__xnor2_1
XFILLER_137_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08285_ _08285_/A vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05497_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05497_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_137_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10935_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07236_ _07236_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07244_/B sky130_fd_sc_hd__xnor2_2
XFILLER_152_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07167_ _07169_/A _07167_/B vssd1 vssd1 vccd1 vccd1 _07195_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06118_ _07848_/A _06033_/X _06117_/X vssd1 vssd1 vccd1 vccd1 _06119_/B sky130_fd_sc_hd__a21oi_1
XFILLER_161_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07098_ _07098_/A _07098_/B vssd1 vssd1 vccd1 vccd1 _07219_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_65_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06049_ _10659_/Q vssd1 vssd1 vccd1 vccd1 _07981_/A sky130_fd_sc_hd__buf_2
XFILLER_114_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08373__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _09876_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09809_/B sky130_fd_sc_hd__or2_1
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09739_ _09802_/C vssd1 vssd1 vccd1 vccd1 _09930_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10483__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10514_ _06163_/X _10497_/B _10513_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10977_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _10951_/Q _10431_/X _10444_/X vssd1 vssd1 vccd1 vccd1 _10951_/D sky130_fd_sc_hd__a21o_1
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10376_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_151_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07415__A _07415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05420_ _10626_/Q _05378_/Y _05380_/Y _05461_/C _05419_/X vssd1 vssd1 vccd1 vccd1
+ _05420_/X sky130_fd_sc_hd__o221a_1
XFILLER_33_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05351_ _10634_/Q vssd1 vssd1 vccd1 vccd1 _07882_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05282_ _10650_/Q vssd1 vssd1 vccd1 vccd1 _06065_/A sky130_fd_sc_hd__clkbuf_2
X_08070_ _08064_/X _08068_/X _08069_/X vssd1 vssd1 vccd1 vccd1 _10681_/D sky130_fd_sc_hd__o21a_1
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07021_ _07021_/A _07030_/C vssd1 vssd1 vccd1 vccd1 _07421_/A sky130_fd_sc_hd__nand2_2
XFILLER_128_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08972_ _08972_/A vssd1 vssd1 vccd1 vccd1 _08972_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_114_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07923_ _10613_/Q _07906_/X _07910_/X _07922_/Y vssd1 vssd1 vccd1 vccd1 _07924_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_68_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07854_ _06185_/A _07849_/X _07850_/X _07852_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ _07854_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_29_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06805_ _06805_/A _06805_/B vssd1 vssd1 vccd1 vccd1 _06818_/A sky130_fd_sc_hd__xor2_4
XFILLER_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07785_ _07785_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _07786_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08107__B1 _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ _09524_/A _09472_/B vssd1 vssd1 vccd1 vccd1 _09625_/B sky130_fd_sc_hd__or2b_1
XFILLER_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06736_ _06736_/A vssd1 vssd1 vccd1 vccd1 _07675_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _09454_/A _09454_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _09456_/C sky130_fd_sc_hd__a21o_1
X_06667_ _06667_/A _06671_/A vssd1 vssd1 vccd1 vccd1 _06686_/A sky130_fd_sc_hd__xnor2_1
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08406_ _08397_/X _10743_/Q _08394_/X _08405_/X vssd1 vssd1 vccd1 vccd1 _10725_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05618_ _10552_/Q _05623_/A _10553_/Q vssd1 vssd1 vccd1 vccd1 _05619_/B sky130_fd_sc_hd__o21ai_1
X_09386_ _09449_/A _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__and3_1
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06598_ _06618_/A _06618_/B vssd1 vssd1 vccd1 vccd1 _06668_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10836__D _10836_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ input36/X _08248_/X _08088_/X _05574_/X _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08337_/X sky130_fd_sc_hd__o221a_1
X_05549_ _05549_/A _05636_/A vssd1 vssd1 vccd1 vccd1 _05629_/B sky130_fd_sc_hd__nand2_1
X_08268_ _08268_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08268_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _10980_/Q _07219_/B vssd1 vssd1 vccd1 vccd1 _07249_/B sky130_fd_sc_hd__and2_1
XFILLER_118_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08199_ _08208_/B _08061_/A _08197_/Y _08198_/Y _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08199_/X sky130_fd_sc_hd__a311o_1
XFILLER_119_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _10246_/B _10228_/A _10291_/S vssd1 vssd1 vccd1 vccd1 _10231_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10161_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10164_/A sky130_fd_sc_hd__xnor2_1
XFILLER_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10092_ _10155_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10093_/B sky130_fd_sc_hd__a21oi_1
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05962__B _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07321__A1 _07560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08821__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10428_ _06206_/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10428_/X sky130_fd_sc_hd__a21bo_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10351_/X _06806_/B _10355_/X _10926_/Q vssd1 vssd1 vccd1 vccd1 _10926_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06060__A1 _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08337__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09344__B _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07570_ _07570_/A _09920_/B _07570_/C vssd1 vssd1 vccd1 vccd1 _07571_/B sky130_fd_sc_hd__or3_1
XFILLER_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06521_ _06521_/A _06521_/B vssd1 vssd1 vccd1 vccd1 _06522_/C sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_13_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09240_ _10820_/Q _09210_/X _09212_/X _09238_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09241_/B sky130_fd_sc_hd__a32o_1
XANTENNA__05323__B1 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06452_ _06626_/A _06568_/B _06451_/C vssd1 vssd1 vccd1 vccd1 _06453_/B sky130_fd_sc_hd__a21oi_1
XFILLER_167_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05403_ _10649_/Q vssd1 vssd1 vccd1 vccd1 _05405_/A sky130_fd_sc_hd__clkinv_2
X_09171_ _05883_/A _09123_/X _09203_/A _09170_/X vssd1 vssd1 vccd1 vccd1 _09171_/X
+ sky130_fd_sc_hd__o211a_1
X_06383_ _06872_/A _06872_/B _06383_/C vssd1 vssd1 vccd1 vccd1 _06874_/A sky130_fd_sc_hd__and3_1
XANTENNA__09065__A1 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08122_ _08114_/X _08130_/B _08116_/Y _08121_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08122_/X sky130_fd_sc_hd__o311a_1
X_05334_ _10672_/Q vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__buf_2
XANTENNA__08812__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ _09403_/A vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__buf_4
XFILLER_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07004_ _07211_/A vssd1 vssd1 vccd1 vccd1 _07188_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_116_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10784_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_115_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08955_ _10963_/Q vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08328__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07906_ _07906_/A vssd1 vssd1 vccd1 vccd1 _07906_/X sky130_fd_sc_hd__clkbuf_1
X_08886_ _08814_/X _08883_/Y _08884_/X _08885_/X vssd1 vssd1 vccd1 vccd1 _10824_/D
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08879__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07837_ _07827_/X _05462_/B _07823_/X _07836_/Y vssd1 vssd1 vccd1 vccd1 _10622_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10804_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07768_ _07768_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07769_/B sky130_fd_sc_hd__xnor2_1
XFILLER_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09270__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ _09507_/A _09676_/C vssd1 vssd1 vccd1 vccd1 _09508_/B sky130_fd_sc_hd__xnor2_4
XFILLER_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10438__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06719_ _06719_/A _06719_/B _06719_/C vssd1 vssd1 vccd1 vccd1 _06720_/B sky130_fd_sc_hd__and3_1
XFILLER_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _09690_/A _09690_/B _07698_/X vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__o21ai_2
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _09438_/Y sky130_fd_sc_hd__nand2_1
XFILLER_158_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09369_ _10889_/Q _10905_/Q vssd1 vssd1 vccd1 vccd1 _09369_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09056__A1 _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10213_ _10950_/Q _10934_/Q vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__and2b_1
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08031__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input42_A io_wbs_m2s_data[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06042__B2 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10144_ _10144_/A _10144_/B vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__xnor2_1
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__xnor2_1
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09531__A2 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10977_ _10977_/CLK _10977_/D vssd1 vssd1 vccd1 vccd1 _10977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05883__A _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07781__A1 _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08740_ _08740_/A _08740_/B _08740_/C vssd1 vssd1 vccd1 vccd1 _08740_/X sky130_fd_sc_hd__and3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07781__B2 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05952_ _10583_/Q vssd1 vssd1 vccd1 vccd1 _06019_/A sky130_fd_sc_hd__buf_6
XFILLER_66_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08671_ _08671_/A vssd1 vssd1 vccd1 vccd1 _08830_/A sky130_fd_sc_hd__clkbuf_2
X_05883_ _05883_/A _10659_/Q _05891_/A vssd1 vssd1 vccd1 vccd1 _05883_/X sky130_fd_sc_hd__or3_1
X_07622_ _07622_/A _07622_/B vssd1 vssd1 vccd1 vccd1 _07623_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07715__A_N _09379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__A _09090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07553_ _07430_/A _07430_/B _07429_/A vssd1 vssd1 vccd1 vccd1 _07558_/B sky130_fd_sc_hd__o21a_1
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08089__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06504_ _06517_/A vssd1 vssd1 vccd1 vccd1 _06758_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_07484_ _07509_/A _07025_/Y _07483_/X vssd1 vssd1 vccd1 vccd1 _07485_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09223_ _09228_/A _09223_/B vssd1 vssd1 vccd1 vccd1 _09224_/A sky130_fd_sc_hd__and2_1
X_06435_ _06435_/A vssd1 vssd1 vccd1 vccd1 _06486_/A sky130_fd_sc_hd__clkinv_2
XFILLER_22_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09154_ _09154_/A vssd1 vssd1 vccd1 vccd1 _09202_/A sky130_fd_sc_hd__clkbuf_4
X_06366_ _10978_/Q _06459_/B vssd1 vssd1 vccd1 vccd1 _06917_/A sky130_fd_sc_hd__nand2_2
X_08105_ _08105_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _08116_/B sky130_fd_sc_hd__nor2_1
X_05317_ _08352_/A _05827_/A vssd1 vssd1 vccd1 vccd1 _05318_/B sky130_fd_sc_hd__nand2_1
XFILLER_147_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09085_ _10937_/Q _09008_/X _08947_/A _10953_/Q vssd1 vssd1 vccd1 vccd1 _09085_/X
+ sky130_fd_sc_hd__a22o_1
X_06297_ _10921_/Q _09356_/A _06416_/A _06302_/B vssd1 vssd1 vccd1 vccd1 _06730_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_162_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08036_ _08236_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _08074_/A sky130_fd_sc_hd__nor2_2
XFILLER_163_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09987_ _09921_/B _09922_/B _09377_/X vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__o21ai_1
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07772__A1 _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08938_ _08938_/A vssd1 vssd1 vccd1 vccd1 _10833_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ _08814_/X _08866_/X _08867_/Y _08868_/X vssd1 vssd1 vccd1 vccd1 _10822_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10900_ _10926_/CLK _10900_/D vssd1 vssd1 vccd1 vccd1 _10900_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09204__S _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _10833_/CLK _10831_/D vssd1 vssd1 vccd1 vccd1 _10831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10762_ _10770_/CLK _10762_/D vssd1 vssd1 vccd1 vccd1 _10762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10693_ _10693_/CLK _10693_/D vssd1 vssd1 vccd1 vccd1 _10693_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06799__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10127_ _10087_/A _10087_/B _10090_/A vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__o21a_1
XFILLER_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10058_ _10487_/A _10123_/B _10057_/C vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__a21oi_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06220_ hold5/A _06223_/B vssd1 vssd1 vccd1 vccd1 _06220_/X sky130_fd_sc_hd__or2_1
XFILLER_145_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06151_ _06151_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_145_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06254__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06082_ _06082_/A _06082_/B _06082_/C _06081_/X vssd1 vssd1 vccd1 vccd1 _06082_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_144_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09910_ _09910_/A _10049_/C vssd1 vssd1 vccd1 vccd1 _09911_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10338__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09841_ _09841_/A _09841_/B vssd1 vssd1 vccd1 vccd1 _09842_/B sky130_fd_sc_hd__nor2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09772_ _09844_/B _09772_/B vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__and2_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ _07083_/A _07061_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _06997_/C sky130_fd_sc_hd__or3_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08919_/B vssd1 vssd1 vccd1 vccd1 _08918_/B sky130_fd_sc_hd__buf_2
X_05935_ _10702_/Q _05935_/B vssd1 vssd1 vccd1 vccd1 _05935_/X sky130_fd_sc_hd__or2_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08654_ _09016_/A _09126_/A vssd1 vssd1 vccd1 vccd1 _08971_/A sky130_fd_sc_hd__nor2_1
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05866_ _05350_/B _05854_/B _05865_/Y vssd1 vssd1 vccd1 vccd1 _05866_/X sky130_fd_sc_hd__o21a_1
XFILLER_27_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07605_ _07708_/A _07605_/B vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__xor2_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08585_ _10781_/Q _10780_/Q _08585_/C vssd1 vssd1 vccd1 vccd1 _08586_/B sky130_fd_sc_hd__and3_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05797_ _08160_/A _05694_/Y _05712_/Y _08146_/A _05713_/X vssd1 vssd1 vccd1 vccd1
+ _05798_/B sky130_fd_sc_hd__o221a_1
XFILLER_35_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07536_ _07617_/B _07618_/B vssd1 vssd1 vccd1 vccd1 _07536_/X sky130_fd_sc_hd__or2_1
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07467_ _07746_/A _07469_/B _07466_/Y vssd1 vssd1 vccd1 vccd1 _07499_/B sky130_fd_sc_hd__o21ai_1
XFILLER_50_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ hold13/A _09168_/X _09203_/X _09205_/X vssd1 vssd1 vccd1 vccd1 _09207_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_139_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06418_ _10921_/Q _07061_/A vssd1 vssd1 vccd1 vccd1 _06418_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08219__C1 _06011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ _07728_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07753_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08164__A _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__D _10844_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ _05461_/C _09136_/X _06212_/B _08150_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09137_/X sky130_fd_sc_hd__a221o_1
XFILLER_120_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06349_ _06436_/A _06568_/B vssd1 vssd1 vccd1 vccd1 _06457_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06245__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09068_ _10968_/Q vssd1 vssd1 vccd1 vccd1 _09639_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08019_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08019_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_134_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08339__A _08339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _10814_/CLK _10814_/D vssd1 vssd1 vccd1 vccd1 _10814_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10745_ _10770_/CLK _10745_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10676_ _10855_/CLK _10676_/D vssd1 vssd1 vccd1 vccd1 _10676_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08074__A _08074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10109__A _10109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08521__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07418__A _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07736__A1 _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05720_ _08082_/A _05536_/B _05737_/B _08082_/B vssd1 vssd1 vccd1 vccd1 _05794_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08161__A1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05651_ _05652_/A _05652_/B _05652_/C vssd1 vssd1 vccd1 vccd1 _05651_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08370_ _10251_/S vssd1 vssd1 vccd1 vccd1 _08547_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05582_ _05769_/A _05582_/B vssd1 vssd1 vccd1 vccd1 _05583_/B sky130_fd_sc_hd__and2_1
X_07321_ _07560_/A _07394_/A _07151_/C vssd1 vssd1 vccd1 vccd1 _07322_/B sky130_fd_sc_hd__a21oi_1
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07252_ _07513_/A _07516_/A vssd1 vssd1 vccd1 vccd1 _07514_/A sky130_fd_sc_hd__or2_1
XFILLER_104_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06203_ _10598_/Q vssd1 vssd1 vccd1 vccd1 _06204_/A sky130_fd_sc_hd__inv_2
XANTENNA__08415__C input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07183_ _07183_/A _07183_/B vssd1 vssd1 vccd1 vccd1 _07208_/A sky130_fd_sc_hd__xnor2_1
XFILLER_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06134_ _06134_/A _06145_/B vssd1 vssd1 vccd1 vccd1 _06134_/Y sky130_fd_sc_hd__nand2_1
XFILLER_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07975__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06065_ _06065_/A vssd1 vssd1 vccd1 vccd1 _06065_/X sky130_fd_sc_hd__buf_4
XFILLER_117_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09824_ _09824_/A _09824_/B vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__xnor2_2
XFILLER_101_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06967_ _07112_/A vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__clkbuf_4
X_09755_ _09755_/A _09755_/B _09755_/C vssd1 vssd1 vccd1 vccd1 _09755_/X sky130_fd_sc_hd__and3_1
XFILLER_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08706_ _10531_/A _08672_/X _08674_/X _08701_/A vssd1 vssd1 vccd1 vccd1 _08706_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_39_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05918_ _08095_/A _05906_/X _05909_/Y _05718_/A _05917_/X vssd1 vssd1 vccd1 vccd1
+ _05918_/X sky130_fd_sc_hd__o221a_1
X_09686_ _09686_/A _09686_/B _09686_/C vssd1 vssd1 vccd1 vccd1 _09686_/X sky130_fd_sc_hd__or3_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06898_ _06930_/A _06930_/B vssd1 vssd1 vccd1 vccd1 _06936_/A sky130_fd_sc_hd__xor2_4
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08152__B2 _08074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _08638_/B _08638_/C _08636_/Y vssd1 vssd1 vccd1 vccd1 _10794_/D sky130_fd_sc_hd__o21a_1
XFILLER_55_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10839__D _10839_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05849_ _10667_/Q _10666_/Q _10665_/Q _05872_/A vssd1 vssd1 vccd1 vccd1 _05863_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07998__A _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ _08568_/A vssd1 vssd1 vccd1 vccd1 _10775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07519_ _09303_/B _07519_/B vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__or2_1
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08499_ _08498_/X _08496_/X _08494_/X _10748_/Q vssd1 vssd1 vccd1 vccd1 _10748_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10530_ _07732_/A _10522_/X _10528_/X _10529_/X vssd1 vssd1 vccd1 vccd1 _10982_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_128_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10461_ _10957_/Q _10469_/B vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or2_1
XFILLER_136_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06126__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07937__S _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10392_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06142__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05981__A _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08143__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08143__B2 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10728_ _10728_/CLK _10728_/D vssd1 vssd1 vccd1 vccd1 _10728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10659_ _10665_/CLK _10659_/D vssd1 vssd1 vccd1 vccd1 _10659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09628__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07870_ _07906_/A vssd1 vssd1 vccd1 vccd1 _07870_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_122_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06821_ _06821_/A _06821_/B vssd1 vssd1 vccd1 vccd1 _06823_/B sky130_fd_sc_hd__xor2_1
XFILLER_84_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09540_ _09458_/A _09599_/A _09696_/A vssd1 vssd1 vccd1 vccd1 _09542_/C sky130_fd_sc_hd__nand3b_1
XFILLER_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06752_ _06752_/A _06752_/B _06752_/C _06746_/A vssd1 vssd1 vccd1 vccd1 _06806_/A
+ sky130_fd_sc_hd__or4b_1
XANTENNA__08134__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05703_ _10693_/Q vssd1 vssd1 vccd1 vccd1 _08188_/A sky130_fd_sc_hd__clkbuf_2
X_09471_ _09471_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09472_/B sky130_fd_sc_hd__and2_1
X_06683_ _06945_/A _06945_/B _06948_/A vssd1 vssd1 vccd1 vccd1 _06943_/C sky130_fd_sc_hd__or3_1
XFILLER_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08422_ _10763_/Q _10764_/Q _08421_/Y vssd1 vssd1 vccd1 vccd1 _08424_/A sky130_fd_sc_hd__o21ai_2
X_05634_ _10685_/Q vssd1 vssd1 vccd1 vccd1 _06037_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08353_ _08037_/A _06115_/B _08351_/Y _08352_/Y vssd1 vssd1 vccd1 vccd1 _08353_/X
+ sky130_fd_sc_hd__a31o_1
X_05565_ _10570_/Q _05576_/A _10571_/Q vssd1 vssd1 vccd1 vccd1 _05566_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07304_ _07289_/A _07304_/B vssd1 vssd1 vccd1 vccd1 _07305_/A sky130_fd_sc_hd__and2b_1
XFILLER_165_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08284_ _08284_/A _08284_/B vssd1 vssd1 vccd1 vccd1 _10702_/D sky130_fd_sc_hd__nor2_1
X_05496_ _05380_/Y _05489_/X _05495_/X _05461_/C vssd1 vssd1 vccd1 vccd1 _10550_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07235_ _07515_/A _07235_/B _07235_/C vssd1 vssd1 vccd1 vccd1 _07237_/B sky130_fd_sc_hd__and3b_1
XFILLER_165_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07166_ _07166_/A _07166_/B vssd1 vssd1 vccd1 vccd1 _07334_/A sky130_fd_sc_hd__nand2_2
XFILLER_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06117_ _08065_/B _08258_/A _06117_/C _06117_/D vssd1 vssd1 vccd1 vccd1 _06117_/X
+ sky130_fd_sc_hd__and4b_2
X_07097_ _10913_/Q _07102_/A vssd1 vssd1 vccd1 vccd1 _07098_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06048_ _10710_/Q _08032_/A _06045_/X _06047_/X vssd1 vssd1 vccd1 vccd1 _06071_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09273__A _09273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09807_ _09807_/A _09856_/C vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10180__A1 _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07999_ input23/X _07987_/X _07998_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10664_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09738_ _09919_/B vssd1 vssd1 vccd1 vccd1 _10129_/B sky130_fd_sc_hd__clkbuf_2
X_09669_ _09731_/A _09669_/B vssd1 vssd1 vccd1 vccd1 _09671_/B sky130_fd_sc_hd__or2_2
XFILLER_43_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06137__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10513_ _10513_/A _10515_/B vssd1 vssd1 vccd1 vccd1 _10513_/X sky130_fd_sc_hd__or2_1
XFILLER_155_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05976__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ _05958_/X _10440_/B _05977_/X vssd1 vssd1 vccd1 vccd1 _10444_/X sky130_fd_sc_hd__a21o_1
XFILLER_171_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08352__A _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10375_ _10932_/Q _10379_/B vssd1 vssd1 vccd1 vccd1 _10375_/X sky130_fd_sc_hd__and2_1
XFILLER_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06611__B2 _06769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10171__A1 _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10122__A _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07431__A _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05350_ _10667_/Q _05350_/B vssd1 vssd1 vccd1 vccd1 _05350_/X sky130_fd_sc_hd__xor2_2
XFILLER_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05281_ _10575_/Q vssd1 vssd1 vccd1 vccd1 _05454_/A sky130_fd_sc_hd__inv_2
XFILLER_174_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07020_ _07021_/A _07020_/B vssd1 vssd1 vccd1 vccd1 _07509_/A sky130_fd_sc_hd__nand2_2
XFILLER_134_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08971_ _08971_/A _08971_/B vssd1 vssd1 vccd1 vccd1 _08972_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07922_ _07922_/A vssd1 vssd1 vccd1 vccd1 _07922_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09093__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07853_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07853_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06804_ _06804_/A vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__buf_2
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07784_ _10510_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _07785_/B sky130_fd_sc_hd__nand2_1
XFILLER_25_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09523_ _10131_/A vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__clkbuf_2
X_06735_ _06735_/A _06735_/B vssd1 vssd1 vccd1 vccd1 _06746_/A sky130_fd_sc_hd__xor2_4
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06118__B1 _06117_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09454_ _09454_/A _09454_/B _09454_/C vssd1 vssd1 vccd1 vccd1 _09456_/B sky130_fd_sc_hd__nand3_1
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06666_ _06666_/A _06666_/B vssd1 vssd1 vccd1 vccd1 _06667_/A sky130_fd_sc_hd__nand2_1
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08405_ _08408_/A _10759_/Q vssd1 vssd1 vccd1 vccd1 _08405_/X sky130_fd_sc_hd__or2_1
X_05617_ _10552_/Q _05623_/A vssd1 vssd1 vccd1 vccd1 _05617_/X sky130_fd_sc_hd__xor2_1
X_09385_ _09810_/A _09383_/A _09417_/A vssd1 vssd1 vccd1 vccd1 _09533_/C sky130_fd_sc_hd__a21o_1
XFILLER_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06597_ _06549_/A _06597_/B _06597_/C vssd1 vssd1 vccd1 vccd1 _06618_/B sky130_fd_sc_hd__nand3b_1
XFILLER_51_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08336_ _05574_/X _08339_/C _08335_/Y vssd1 vssd1 vccd1 vccd1 _08336_/Y sky130_fd_sc_hd__a21oi_1
X_05548_ _10546_/Q _05635_/B vssd1 vssd1 vccd1 vccd1 _05636_/A sky130_fd_sc_hd__nor2_1
X_08267_ _08267_/A _08267_/B vssd1 vssd1 vccd1 vccd1 _08267_/Y sky130_fd_sc_hd__nand2_1
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05479_ _05479_/A vssd1 vssd1 vccd1 vccd1 _05489_/A sky130_fd_sc_hd__clkbuf_2
X_07218_ _07222_/A _07215_/B _07216_/B _10979_/Q vssd1 vssd1 vccd1 vccd1 _07218_/X
+ sky130_fd_sc_hd__a22o_1
X_08198_ _08198_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07149_ _07511_/A _07327_/A _07149_/C vssd1 vssd1 vccd1 vccd1 _07150_/B sky130_fd_sc_hd__and3b_1
XANTENNA__10852__D _10852_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10207__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10091_ _10155_/A _10091_/B _10091_/C vssd1 vssd1 vccd1 vccd1 _10121_/S sky130_fd_sc_hd__and3_1
XFILLER_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08082__A _08082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10427_ _10946_/Q _10427_/B vssd1 vssd1 vccd1 vccd1 _10427_/X sky130_fd_sc_hd__and2_1
XFILLER_171_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10117__A _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10358_ _10351_/X _06752_/A _10355_/X _10925_/Q vssd1 vssd1 vccd1 vccd1 _10925_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06060__A2 _08023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10289_ _10289_/A _10289_/B vssd1 vssd1 vccd1 vccd1 _10289_/X sky130_fd_sc_hd__or2_1
XANTENNA__08337__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10954_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06984__B _07061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06520_ _06532_/A _06523_/B _06523_/C vssd1 vssd1 vccd1 vccd1 _06520_/X sky130_fd_sc_hd__a21o_1
XFILLER_46_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07161__A _10982_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06451_ _06456_/A _06568_/B _06451_/C vssd1 vssd1 vccd1 vccd1 _06453_/A sky130_fd_sc_hd__and3_1
XANTENNA__05323__A1 _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05402_ _10618_/Q _05483_/A vssd1 vssd1 vccd1 vccd1 _05402_/X sky130_fd_sc_hd__or2_1
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09170_ _05460_/D _09136_/X _09148_/X _08180_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09170_/X sky130_fd_sc_hd__a221o_1
X_06382_ _06394_/A _06382_/B vssd1 vssd1 vccd1 vccd1 _06383_/C sky130_fd_sc_hd__or2_1
XFILLER_159_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08121_ _08132_/B _08061_/A _08117_/Y _08119_/Y _08120_/X vssd1 vssd1 vccd1 vccd1
+ _08121_/X sky130_fd_sc_hd__a311o_1
X_05333_ _10640_/Q vssd1 vssd1 vccd1 vccd1 _07903_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08052_ _08052_/A vssd1 vssd1 vccd1 vccd1 _08052_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07003_ _10981_/Q vssd1 vssd1 vccd1 vccd1 _07211_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_116_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08954_ _09098_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _10474_/B sky130_fd_sc_hd__nor2_2
XANTENNA__08328__A1 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ _07916_/A _07905_/B vssd1 vssd1 vccd1 vccd1 _10640_/D sky130_fd_sc_hd__nor2_1
XFILLER_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08885_ input33/X _08819_/X _08820_/X _10824_/Q _10412_/A vssd1 vssd1 vccd1 vccd1
+ _08885_/X sky130_fd_sc_hd__o221a_1
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10135__B2 _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07836_ _06165_/A _07828_/X _07829_/X _07835_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07836_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_99_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07767_ _10506_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _07768_/B sky130_fd_sc_hd__nand2_1
X_09506_ _09506_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09676_/C sky130_fd_sc_hd__nor2_2
X_06718_ _06718_/A _06718_/B vssd1 vssd1 vccd1 vccd1 _06720_/A sky130_fd_sc_hd__nand2_1
X_07698_ _07698_/A _07698_/B vssd1 vssd1 vccd1 vccd1 _07698_/X sky130_fd_sc_hd__or2_1
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10847__D _10847_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09437_ _09437_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__or2_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06649_ _06663_/A _06692_/A _06692_/B _06622_/B vssd1 vssd1 vccd1 vccd1 _06650_/C
+ sky130_fd_sc_hd__a31o_1
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09368_ _09676_/A _09546_/A _09546_/B _09367_/Y _09356_/A vssd1 vssd1 vccd1 vccd1
+ _09607_/A sky130_fd_sc_hd__a32o_2
XFILLER_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08319_ _08324_/B _08253_/X _08317_/Y _08318_/Y vssd1 vssd1 vccd1 vccd1 _08319_/X
+ sky130_fd_sc_hd__a31o_1
X_09299_ _10343_/A _09299_/B vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__and2_1
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06134__B _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10212_ _10934_/Q _10950_/Q vssd1 vssd1 vccd1 vccd1 _10226_/B sky130_fd_sc_hd__or2b_1
XFILLER_107_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10143_ _10143_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10144_/B sky130_fd_sc_hd__xnor2_1
XFILLER_122_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input35_A io_wbs_m2s_data[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10074_ _10074_/A _10074_/B vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06150__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10429__A2 _10727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ _10976_/CLK _10976_/D vssd1 vssd1 vccd1 vccd1 _10976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05951_ _05717_/X _05788_/X _05809_/X _05950_/Y vssd1 vssd1 vccd1 vccd1 _10540_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08670_ _08670_/A _08670_/B _08670_/C vssd1 vssd1 vccd1 vccd1 _08670_/X sky130_fd_sc_hd__and3_1
X_05882_ _10658_/Q _05895_/A vssd1 vssd1 vccd1 vccd1 _05891_/A sky130_fd_sc_hd__or2_1
XFILLER_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06995__A _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08730__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07621_ _07621_/A _07702_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__xnor2_2
XFILLER_66_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07552_ _07448_/A _07448_/B _07447_/A vssd1 vssd1 vccd1 vccd1 _07583_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__10838__CLK _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06503_ _06503_/A _06503_/B vssd1 vssd1 vccd1 vccd1 _06503_/Y sky130_fd_sc_hd__nor2_1
X_07483_ _07442_/X _07728_/B _07729_/B _07715_/C vssd1 vssd1 vccd1 vccd1 _07483_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09222_ hold3/A _09210_/X _09212_/X _09221_/X _09203_/X vssd1 vssd1 vccd1 vccd1 _09223_/B
+ sky130_fd_sc_hd__a32o_1
X_06434_ _06434_/A _06434_/B vssd1 vssd1 vccd1 vccd1 _06435_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _10844_/D sky130_fd_sc_hd__nor2_4
XANTENNA__08246__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06365_ _07682_/B _06365_/B _06451_/C _06367_/A vssd1 vssd1 vccd1 vccd1 _06872_/B
+ sky130_fd_sc_hd__or4b_2
X_08104_ _08105_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _08104_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05316_ _08034_/A _05318_/A vssd1 vssd1 vccd1 vccd1 _05525_/B sky130_fd_sc_hd__xnor2_4
X_09084_ _09908_/A vssd1 vssd1 vccd1 vccd1 _10491_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06296_ _10922_/Q _10905_/Q vssd1 vssd1 vccd1 vccd1 _06302_/B sky130_fd_sc_hd__and2_1
XFILLER_147_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08035_ input40/X _07985_/B _08034_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10679_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09986_ _09925_/A _09924_/B _10131_/A vssd1 vssd1 vccd1 vccd1 _09990_/A sky130_fd_sc_hd__o21ai_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08937_ _10832_/Q _10529_/A vssd1 vssd1 vccd1 vccd1 _08938_/A sky130_fd_sc_hd__and2_1
XFILLER_57_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08868_ input31/X _08819_/X _08820_/X _10822_/Q _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08868_/X sky130_fd_sc_hd__o221a_1
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07819_ _06255_/X _09020_/A _06257_/X _07818_/Y vssd1 vssd1 vccd1 vccd1 _10618_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08799_ _06206_/X _08785_/X _08786_/X _10814_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08799_/X sky130_fd_sc_hd__o221a_1
X_10830_ _10830_/CLK _10830_/D vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10761_ _10935_/CLK _10761_/D vssd1 vssd1 vccd1 vccd1 _10761_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10692_ _10693_/CLK _10692_/D vssd1 vssd1 vccd1 vccd1 _10692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05968__B input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06248__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10347__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10126_ _10126_/A _10126_/B vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__nand2_1
XFILLER_110_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10057_ _10057_/A _10123_/B _10057_/C vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__and3_1
XFILLER_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ _10962_/CLK _10959_/D vssd1 vssd1 vccd1 vccd1 _10959_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10792_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08535__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_3_0_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08779__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06150_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06170_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09440__A2 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10807_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__06254__A2 _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06081_ _08282_/A _05851_/A _08198_/A _08196_/A _06080_/X vssd1 vssd1 vccd1 vccd1
+ _06081_/X sky130_fd_sc_hd__o221a_1
XFILLER_144_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09840_ _09974_/A _09839_/B _09839_/C vssd1 vssd1 vccd1 vccd1 _09841_/B sky130_fd_sc_hd__a21oi_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09771_/A _09771_/B _09771_/C vssd1 vssd1 vccd1 vccd1 _09772_/B sky130_fd_sc_hd__or3_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _07066_/A _07056_/A _10901_/Q _07475_/B vssd1 vssd1 vccd1 vccd1 _07060_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_101_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08722_ _08902_/B vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__clkbuf_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05934_ _08251_/B _05863_/X _05867_/X _05932_/X _05933_/X vssd1 vssd1 vccd1 vccd1
+ _05934_/X sky130_fd_sc_hd__o221a_1
XFILLER_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08653_ _08651_/Y _08649_/C _08652_/X vssd1 vssd1 vccd1 vccd1 _10798_/D sky130_fd_sc_hd__a21oi_1
X_05865_ _05358_/A _05823_/A _10666_/Q vssd1 vssd1 vccd1 vccd1 _05865_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07604_ _07604_/A _07604_/B vssd1 vssd1 vccd1 vccd1 _07605_/B sky130_fd_sc_hd__xor2_4
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08584_ _10780_/Q _08585_/C _08583_/Y vssd1 vssd1 vccd1 vccd1 _10780_/D sky130_fd_sc_hd__o21a_1
XANTENNA__06190__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05796_ _05788_/B _05794_/Y _05795_/Y vssd1 vssd1 vccd1 vccd1 _05796_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07535_ _07535_/A _07535_/B vssd1 vssd1 vccd1 vccd1 _07618_/B sky130_fd_sc_hd__nor2_2
XFILLER_35_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07466_ _07466_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07466_/Y sky130_fd_sc_hd__nand2_1
XFILLER_168_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08445__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06417_ _09356_/A vssd1 vssd1 vccd1 vccd1 _07061_/A sky130_fd_sc_hd__clkbuf_4
X_09205_ _07998_/A _09204_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09205_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07397_ _07397_/A _07397_/B vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__xnor2_1
XFILLER_136_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06348_ _06547_/C vssd1 vssd1 vccd1 vccd1 _06568_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _09136_/A vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _07727_/A _08965_/Y _09036_/X _09063_/X _09066_/X vssd1 vssd1 vccd1 vccd1
+ _09067_/X sky130_fd_sc_hd__a221o_1
XFILLER_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06279_ _06558_/B _06558_/C vssd1 vssd1 vccd1 vccd1 _06338_/A sky130_fd_sc_hd__and2_1
XFILLER_162_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08018_ _08018_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08018_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08180__A _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _09969_/A _09969_/B vssd1 vssd1 vccd1 vccd1 _10039_/A sky130_fd_sc_hd__xnor2_2
XFILLER_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09215__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06181__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _10942_/CLK _10813_/D vssd1 vssd1 vccd1 vccd1 _10813_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10744_ _10770_/CLK _10744_/D vssd1 vssd1 vccd1 vccd1 _10744_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10675_ _10855_/CLK _10675_/D vssd1 vssd1 vccd1 vccd1 _10675_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_127_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10109_ _10109_/A _10109_/B vssd1 vssd1 vccd1 vccd1 _10162_/B sky130_fd_sc_hd__xor2_1
XFILLER_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08161__A2 _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05650_ _10683_/Q vssd1 vssd1 vccd1 vccd1 _05718_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05581_ _10567_/Q _05582_/B vssd1 vssd1 vccd1 vccd1 _05681_/B sky130_fd_sc_hd__nor2_1
X_07320_ _07341_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07488_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08265__A _08267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07251_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__nand2_1
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06202_ input21/X vssd1 vssd1 vccd1 vccd1 _06202_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07182_ _07183_/A _07183_/B vssd1 vssd1 vccd1 vccd1 _07280_/B sky130_fd_sc_hd__and2_1
XFILLER_158_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06133_ _06149_/A vssd1 vssd1 vccd1 vccd1 _06145_/B sky130_fd_sc_hd__buf_4
XFILLER_117_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06064_ _05767_/Y _10675_/Q _06050_/X _09104_/A vssd1 vssd1 vccd1 vccd1 _06069_/C
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08924__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09823_ _10876_/Q _09572_/X _09822_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10876_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09754_ _09754_/A _09754_/B vssd1 vssd1 vccd1 vccd1 _09755_/C sky130_fd_sc_hd__xnor2_1
XFILLER_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06966_ _06966_/A _06966_/B vssd1 vssd1 vccd1 vccd1 _07708_/A sky130_fd_sc_hd__xnor2_4
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08705_ _08808_/A _08705_/B _08725_/A vssd1 vssd1 vccd1 vccd1 _08705_/X sky130_fd_sc_hd__or3_1
X_05917_ _05718_/A _05909_/Y _05911_/Y _05719_/A _05916_/X vssd1 vssd1 vccd1 vccd1
+ _05917_/X sky130_fd_sc_hd__a221o_1
XFILLER_100_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09685_ _09689_/A _09685_/B vssd1 vssd1 vccd1 vccd1 _09686_/C sky130_fd_sc_hd__xnor2_1
X_06897_ _06894_/A _06894_/B _06899_/A _06899_/B vssd1 vssd1 vccd1 vccd1 _06930_/B
+ sky130_fd_sc_hd__a22oi_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08636_ _08638_/B _08638_/C _08592_/A vssd1 vssd1 vccd1 vccd1 _08636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_54_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05848_ _06052_/A _05848_/B _05886_/B vssd1 vssd1 vccd1 vccd1 _05872_/A sky130_fd_sc_hd__or3_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _08432_/Y _08565_/X _08567_/C _08567_/D vssd1 vssd1 vccd1 vccd1 _08568_/A
+ sky130_fd_sc_hd__and4bb_1
X_05779_ _08355_/A _10571_/Q _10572_/Q _05778_/Y vssd1 vssd1 vccd1 vccd1 _05785_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07518_ _07573_/A _07394_/X _07327_/X _07021_/A vssd1 vssd1 vccd1 vccd1 _07519_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08175__A _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08498_ _10785_/Q vssd1 vssd1 vccd1 vccd1 _08498_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07449_ _07562_/C _07573_/C _07373_/A vssd1 vssd1 vccd1 vccd1 _07551_/B sky130_fd_sc_hd__o21ai_2
XFILLER_155_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10460_ _10472_/B vssd1 vssd1 vccd1 vccd1 _10469_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10263__A_N _10939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09119_ _10500_/B vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10391_ _10533_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10391_/X sky130_fd_sc_hd__a21bo_1
XFILLER_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08143__A2 _08086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06154__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10727_ _10804_/CLK _10727_/D vssd1 vssd1 vccd1 vccd1 _10727_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_174_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10658_ _10665_/CLK _10658_/D vssd1 vssd1 vccd1 vccd1 _10658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10589_ _10970_/CLK _10589_/D vssd1 vssd1 vccd1 vccd1 _10589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09159__B2 _05692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06090__B1 _10579_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06820_ _07779_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _06821_/B sky130_fd_sc_hd__xor2_2
XFILLER_68_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07164__A _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06751_ _06748_/X _06772_/A _06771_/B vssd1 vssd1 vccd1 vccd1 _06779_/A sky130_fd_sc_hd__o21ai_1
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05702_ _05702_/A _10556_/Q vssd1 vssd1 vccd1 vccd1 _05702_/X sky130_fd_sc_hd__and2_1
X_09470_ _09520_/A _09470_/B vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__and2_1
X_06682_ _06947_/A _06947_/B vssd1 vssd1 vccd1 vccd1 _06948_/A sky130_fd_sc_hd__or2_1
XFILLER_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08421_ _10763_/Q _10764_/Q _10765_/Q vssd1 vssd1 vccd1 vccd1 _08421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05633_ _10686_/Q vssd1 vssd1 vccd1 vccd1 _05726_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05564_ _05564_/A _05566_/A vssd1 vssd1 vccd1 vccd1 _05564_/Y sky130_fd_sc_hd__xnor2_1
X_08352_ _08352_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08352_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07303_ _07307_/A _07307_/B vssd1 vssd1 vccd1 vccd1 _07349_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ _08274_/Y _08248_/X _08157_/A _08281_/X _08282_/X vssd1 vssd1 vccd1 vccd1
+ _08284_/B sky130_fd_sc_hd__o221a_1
X_05495_ _05495_/A vssd1 vssd1 vccd1 vccd1 _05495_/X sky130_fd_sc_hd__clkbuf_2
X_07234_ _10981_/Q _07382_/A vssd1 vssd1 vccd1 vccd1 _07515_/A sky130_fd_sc_hd__and2_1
XANTENNA__09819__A _09819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ _07196_/A vssd1 vssd1 vccd1 vccd1 _07184_/A sky130_fd_sc_hd__inv_2
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06116_ _08062_/A _08036_/B vssd1 vssd1 vccd1 vccd1 _06117_/D sky130_fd_sc_hd__or2_2
XFILLER_145_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07096_ _07363_/C _07096_/B vssd1 vssd1 vccd1 vccd1 _07355_/A sky130_fd_sc_hd__and2_1
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06081__B1 _08198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06047_ _08209_/A _05702_/A _10704_/Q _08018_/A vssd1 vssd1 vccd1 vccd1 _06047_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09806_ _09807_/A _09856_/C vssd1 vssd1 vccd1 vccd1 _09876_/A sky130_fd_sc_hd__and2_1
XFILLER_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07998_ _07998_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _07998_/X sky130_fd_sc_hd__or2_1
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09737_ _09737_/A vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06949_ _06591_/Y _06949_/B vssd1 vssd1 vccd1 vccd1 _06950_/A sky130_fd_sc_hd__and2b_1
XFILLER_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09669_/B sky130_fd_sc_hd__and2_1
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08619_ _08617_/X _08649_/A _08619_/C vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__and3b_1
XFILLER_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09599_ _09599_/A _09599_/B vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__nand2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09086__A0 _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08833__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10512_ _05982_/A _10497_/B _10510_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10976_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_128_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10443_ _06147_/X _10431_/X _10440_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10950_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08352__B _08352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06153__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _10365_/X _10712_/Q _10368_/X _10372_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10931_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05992__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 _10856_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05280_ _10575_/Q vssd1 vssd1 vccd1 vccd1 _05910_/B sky130_fd_sc_hd__buf_2
XFILLER_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06063__B1 _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08970_ _07715_/C _08943_/X _08967_/Y _08969_/Y vssd1 vssd1 vccd1 vccd1 _08970_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_115_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07921_ _08284_/A _07921_/B vssd1 vssd1 vccd1 vccd1 _10644_/D sky130_fd_sc_hd__nor2_1
XFILLER_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07852_ _10876_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06803_ _07682_/A vssd1 vssd1 vccd1 vccd1 _07780_/C sky130_fd_sc_hd__buf_2
Xinput1 io_ba_match vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
XFILLER_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07783_ _10513_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07785_/A sky130_fd_sc_hd__nand2_1
XFILLER_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _09563_/B _09522_/B vssd1 vssd1 vccd1 vccd1 _09625_/A sky130_fd_sc_hd__and2_1
X_06734_ _06734_/A _06734_/B vssd1 vssd1 vccd1 vccd1 _06735_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06118__A1 _07848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _09390_/A _09488_/A _10964_/Q vssd1 vssd1 vccd1 vccd1 _09454_/C sky130_fd_sc_hd__and3b_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06665_ _06700_/B _06665_/B vssd1 vssd1 vccd1 vccd1 _06903_/A sky130_fd_sc_hd__xnor2_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08404_ _08397_/X _10742_/Q _08394_/X _08403_/X vssd1 vssd1 vccd1 vccd1 _10724_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05616_ _10691_/Q vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09384_ _09417_/A _09810_/A _09424_/A vssd1 vssd1 vccd1 vccd1 _09533_/B sky130_fd_sc_hd__nand3_2
XANTENNA__06238__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06596_ _06599_/A _06599_/B vssd1 vssd1 vccd1 vccd1 _06597_/C sky130_fd_sc_hd__or2_1
XFILLER_101_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08335_ _05574_/X _08339_/C _08092_/A vssd1 vssd1 vccd1 vccd1 _08335_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_51_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05547_ _05547_/A _05637_/B vssd1 vssd1 vccd1 vccd1 _05635_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08266_ _08267_/A _08277_/C vssd1 vssd1 vccd1 vccd1 _08266_/Y sky130_fd_sc_hd__nor2_1
X_05478_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05495_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07217_ _07250_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _07217_/Y sky130_fd_sc_hd__nor2_1
XFILLER_153_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08197_ _08191_/A _08191_/B _05877_/X vssd1 vssd1 vccd1 vccd1 _08197_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_106_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07148_ _07148_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07152_/B sky130_fd_sc_hd__or2_1
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06054__B1 _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07079_ _07163_/B _07312_/A _07149_/C vssd1 vssd1 vccd1 vccd1 _07298_/A sky130_fd_sc_hd__or3b_1
XFILLER_160_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10090_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10091_/C sky130_fd_sc_hd__and2_1
XFILLER_59_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05317__A _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09231__A0 _05598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10426_ _10408_/X _10726_/Q _10424_/X _10425_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10945_/D sky130_fd_sc_hd__o221a_1
XFILLER_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10117__B _10117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10357_ _09634_/A _06746_/A _08494_/X _10924_/Q vssd1 vssd1 vccd1 vccd1 _10924_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_140_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10288_ _10265_/A _10287_/C _10287_/D vssd1 vssd1 vccd1 vccd1 _10289_/B sky130_fd_sc_hd__a21bo_1
XFILLER_111_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06450_ _06468_/A _06450_/B vssd1 vssd1 vccd1 vccd1 _06477_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05401_ _05401_/A _05406_/A vssd1 vssd1 vccd1 vccd1 _05483_/A sky130_fd_sc_hd__xnor2_1
X_06381_ _06895_/A _06895_/B _06381_/C vssd1 vssd1 vccd1 vccd1 _06382_/B sky130_fd_sc_hd__and3_1
XFILLER_159_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05332_ _08021_/A _05844_/B vssd1 vssd1 vccd1 vccd1 _05332_/Y sky130_fd_sc_hd__xnor2_1
X_08120_ _08236_/A vssd1 vssd1 vccd1 vccd1 _08120_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08051_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08052_/A sky130_fd_sc_hd__clkbuf_4
X_07002_ _07562_/C _07573_/C vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__xor2_1
XFILLER_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06036__B1 _05405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08953_ _10914_/Q _10931_/Q _09008_/A vssd1 vssd1 vccd1 vccd1 _08953_/X sky130_fd_sc_hd__mux2_1
XFILLER_131_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07904_ _10608_/Q _07888_/X _07892_/X _07903_/Y vssd1 vssd1 vccd1 vccd1 _07905_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08884_ _08883_/A _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08884_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__10043__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07835_ _10872_/Q _07845_/B vssd1 vssd1 vccd1 vccd1 _07835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07766_ _10504_/A _07766_/B vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09505_ _07066_/A _10887_/Q vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__and2b_1
X_06717_ _06717_/A _06717_/B vssd1 vssd1 vccd1 vccd1 _06718_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07697_ _07637_/A _07637_/B _07696_/X vssd1 vssd1 vccd1 vccd1 _09690_/B sky130_fd_sc_hd__o21a_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09477_/B vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__xnor2_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06648_ _06648_/A _06648_/B vssd1 vssd1 vccd1 vccd1 _06650_/B sky130_fd_sc_hd__xor2_1
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _10888_/Q vssd1 vssd1 vccd1 vccd1 _09367_/Y sky130_fd_sc_hd__inv_2
X_06579_ _06581_/A _06581_/C _06581_/B vssd1 vssd1 vccd1 vccd1 _06579_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08318_ _08318_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08318_/Y sky130_fd_sc_hd__nor2_1
XFILLER_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09298_ hold11/X _09274_/X _09275_/X _09297_/X _09127_/X vssd1 vssd1 vccd1 vccd1
+ _09299_/B sky130_fd_sc_hd__a32o_1
XFILLER_166_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08249_ input26/X _08248_/X _08088_/X _08243_/A _08394_/A vssd1 vssd1 vccd1 vccd1
+ _08249_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10218__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10211_ _10209_/Y _10210_/X _07747_/A _09406_/X vssd1 vssd1 vccd1 vccd1 _10900_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10142_ _10142_/A _10142_/B vssd1 vssd1 vccd1 vccd1 _10143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_97_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10074_/B sky130_fd_sc_hd__nor2_1
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input28_A io_wbs_m2s_data[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10975_ _10976_/CLK _10975_/D vssd1 vssd1 vccd1 vccd1 _10975_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05510__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08007__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ _10427_/B vssd1 vssd1 vccd1 vccd1 _10424_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05950_ _05528_/X _05826_/X _05949_/X vssd1 vssd1 vccd1 vccd1 _05950_/Y sky130_fd_sc_hd__a21oi_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05881_ _06039_/A _10656_/Q _05900_/A vssd1 vssd1 vccd1 vccd1 _05895_/A sky130_fd_sc_hd__or3_1
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07702_/B sky130_fd_sc_hd__xnor2_4
XFILLER_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08268__A _08268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07551_ _07450_/A _07551_/B vssd1 vssd1 vccd1 vccd1 _07585_/A sky130_fd_sc_hd__and2b_1
XFILLER_35_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06502_ _06561_/B _06502_/B _06502_/C _06506_/B vssd1 vssd1 vccd1 vccd1 _06503_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_62_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07482_ _07482_/A _07482_/B vssd1 vssd1 vccd1 vccd1 _07485_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _08235_/A _09220_/X _09226_/S vssd1 vssd1 vccd1 vccd1 _09221_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06433_ _06645_/A _06433_/B vssd1 vssd1 vccd1 vccd1 _06434_/B sky130_fd_sc_hd__or2_1
XANTENNA__09099__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _09112_/X _09147_/Y _09151_/X vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__a21oi_1
X_06364_ _06719_/A _06460_/B vssd1 vssd1 vccd1 vccd1 _06367_/A sky130_fd_sc_hd__nand2_1
XFILLER_159_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08103_ _08117_/B _08102_/Y _06117_/D vssd1 vssd1 vccd1 vccd1 _08103_/Y sky130_fd_sc_hd__a21oi_1
X_05315_ _08352_/A _05827_/A vssd1 vssd1 vccd1 vccd1 _05318_/A sky130_fd_sc_hd__or2_2
XFILLER_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09083_ _09764_/A vssd1 vssd1 vccd1 vccd1 _09908_/A sky130_fd_sc_hd__clkbuf_2
X_06295_ _10922_/Q _10905_/Q vssd1 vssd1 vccd1 vccd1 _06416_/A sky130_fd_sc_hd__or2_1
X_08034_ _08034_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09985_ _09985_/A _10046_/A vssd1 vssd1 vccd1 vccd1 _10021_/A sky130_fd_sc_hd__xnor2_1
XFILLER_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08936_ _08936_/A vssd1 vssd1 vccd1 vccd1 _10832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08867_ _08866_/A _08866_/B _08870_/D vssd1 vssd1 vccd1 vccd1 _08867_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_85_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07818_ _06145_/A _06258_/X _07807_/X _07817_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07818_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08798_ _08803_/D _08798_/B vssd1 vssd1 vccd1 vccd1 _08798_/X sky130_fd_sc_hd__xor2_1
XFILLER_38_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07749_ _09420_/A _07748_/A _07475_/C _07589_/B _07393_/Y vssd1 vssd1 vccd1 vccd1
+ _07750_/B sky130_fd_sc_hd__a311o_1
XFILLER_53_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10760_ _10935_/CLK _10760_/D vssd1 vssd1 vccd1 vccd1 _10760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07810__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ _09336_/A _09336_/B _09333_/A vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__a21o_1
X_10691_ _10693_/CLK _10691_/D vssd1 vssd1 vccd1 vccd1 _10691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05968__C input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10044__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06145__B _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10929_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10125_ _09940_/B _10077_/A _10077_/B _10078_/A vssd1 vssd1 vccd1 vccd1 _10126_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10056_ _10123_/A _10122_/B _10056_/C vssd1 vssd1 vccd1 vccd1 _10057_/C sky130_fd_sc_hd__and3_1
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07704__B _09898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08088__A _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ _10958_/CLK _10958_/D vssd1 vssd1 vccd1 vccd1 _10958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10889_ _10980_/CLK _10889_/D vssd1 vssd1 vccd1 vccd1 _10889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06080_ _05744_/Y _07998_/A _07979_/A _05709_/Y vssd1 vssd1 vccd1 vccd1 _06080_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_156_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07167__A _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09770_ _09771_/A _09771_/B _09771_/C vssd1 vssd1 vccd1 vccd1 _09844_/B sky130_fd_sc_hd__o21ai_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06982_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__or2_2
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08721_ _08888_/B vssd1 vssd1 vccd1 vccd1 _08902_/B sky130_fd_sc_hd__clkbuf_2
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05933_ _05859_/Y _05857_/B _08251_/A vssd1 vssd1 vccd1 vccd1 _05933_/X sky130_fd_sc_hd__a21o_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08652_ _10798_/Q _10797_/Q _08648_/B _08592_/A vssd1 vssd1 vccd1 vccd1 _08652_/X
+ sky130_fd_sc_hd__a31o_1
X_05864_ _10698_/Q vssd1 vssd1 vccd1 vccd1 _08233_/A sky130_fd_sc_hd__buf_2
XFILLER_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07603_ _07603_/A _07711_/B vssd1 vssd1 vccd1 vccd1 _07604_/B sky130_fd_sc_hd__xnor2_4
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08583_ _08583_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _08583_/Y sky130_fd_sc_hd__nor2_1
XFILLER_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05795_ _05732_/D _05734_/X _05732_/C vssd1 vssd1 vccd1 vccd1 _05795_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_35_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07534_ _07534_/A _07534_/B _07534_/C vssd1 vssd1 vccd1 vccd1 _07535_/B sky130_fd_sc_hd__nor3_1
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07465_ _07466_/A _07466_/B vssd1 vssd1 vccd1 vccd1 _07469_/B sky130_fd_sc_hd__xnor2_1
XFILLER_23_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09204_ _08218_/A _07875_/A _09250_/A vssd1 vssd1 vccd1 vccd1 _09204_/X sky130_fd_sc_hd__mux2_1
X_06416_ _06416_/A _06416_/B vssd1 vssd1 vccd1 vccd1 _06420_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08219__A1 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07396_ _07396_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07397_/B sky130_fd_sc_hd__xnor2_1
XFILLER_33_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09135_ _09113_/X _09134_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09135_/Y sky130_fd_sc_hd__o21ai_1
X_06347_ _06561_/C vssd1 vssd1 vccd1 vccd1 _06547_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09066_ _05482_/X _08972_/A _08974_/A _09065_/X vssd1 vssd1 vccd1 vccd1 _09066_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06278_ _10915_/Q _07102_/A vssd1 vssd1 vccd1 vccd1 _06558_/C sky130_fd_sc_hd__or2_1
X_08017_ input31/X _08015_/X _08016_/X _08006_/X vssd1 vssd1 vccd1 vccd1 _10671_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09968_ _10878_/Q _09572_/X _09967_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10878_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_131_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06953__A1 _06769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08919_ hold9/A _08919_/B vssd1 vssd1 vccd1 vccd1 _08920_/B sky130_fd_sc_hd__or2_1
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09899_ _09899_/A _09899_/B vssd1 vssd1 vccd1 vccd1 _09964_/A sky130_fd_sc_hd__xnor2_2
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10812_ _10814_/CLK _10812_/D vssd1 vssd1 vccd1 vccd1 _10812_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10743_ _10770_/CLK _10743_/D vssd1 vssd1 vccd1 vccd1 _10743_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08355__B _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ _10674_/CLK _10674_/D vssd1 vssd1 vccd1 vccd1 _10674_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05995__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10108_ _09961_/A _10037_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _10109_/B sky130_fd_sc_hd__o21ai_1
XFILLER_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10039_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10039_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10141__A _10484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05580_ _05582_/B _05580_/B vssd1 vssd1 vccd1 vccd1 _05580_/X sky130_fd_sc_hd__and2_1
XFILLER_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07250_ _07250_/A _07250_/B vssd1 vssd1 vccd1 vccd1 _07515_/B sky130_fd_sc_hd__xnor2_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05683__A1 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06201_ _06195_/X _06183_/X _06197_/Y _06200_/X vssd1 vssd1 vccd1 vccd1 _10597_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07181_ _07229_/A _07398_/B _07181_/C vssd1 vssd1 vccd1 vccd1 _07183_/B sky130_fd_sc_hd__and3_1
XFILLER_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06132_ _10584_/Q vssd1 vssd1 vccd1 vccd1 _06134_/A sky130_fd_sc_hd__inv_2
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06063_ _05767_/Y _10675_/Q _08298_/A _05782_/Y vssd1 vssd1 vccd1 vccd1 _06063_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09822_ _09822_/A _09822_/B vssd1 vssd1 vccd1 vccd1 _09822_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09753_ _09753_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09754_/B sky130_fd_sc_hd__xnor2_2
X_06965_ _07609_/A _07615_/A _06962_/X _07624_/A vssd1 vssd1 vccd1 vccd1 _06966_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_39_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08137__B1 _08062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _08709_/A _08704_/B _08704_/C vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__nor3_1
XFILLER_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05916_ _05719_/A _05911_/Y _05913_/Y _08082_/C _05915_/X vssd1 vssd1 vccd1 vccd1
+ _05916_/X sky130_fd_sc_hd__o221a_1
X_09684_ _09684_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09685_/B sky130_fd_sc_hd__xnor2_1
X_06896_ _06896_/A _06896_/B vssd1 vssd1 vccd1 vccd1 _06899_/B sky130_fd_sc_hd__nor2_2
XFILLER_66_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ _08635_/A vssd1 vssd1 vccd1 vccd1 _10793_/D sky130_fd_sc_hd__clkbuf_1
X_05847_ _10670_/Q vssd1 vssd1 vccd1 vccd1 _05851_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _10775_/Q _08578_/C vssd1 vssd1 vccd1 vccd1 _08567_/C sky130_fd_sc_hd__or2_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05778_ _10711_/Q vssd1 vssd1 vccd1 vccd1 _05778_/Y sky130_fd_sc_hd__clkinv_2
X_07517_ _07517_/A vssd1 vssd1 vccd1 vccd1 _09303_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_168_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08497_ _10784_/Q _08496_/X _08494_/X _10747_/Q vssd1 vssd1 vccd1 vccd1 _10747_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07448_ _07448_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07450_/A sky130_fd_sc_hd__xnor2_2
XFILLER_168_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10684_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05674__A1 _05598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07379_ _07474_/B _07459_/B _07748_/B vssd1 vssd1 vccd1 vccd1 _07381_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09118_ _09118_/A vssd1 vssd1 vccd1 vccd1 _10500_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10390_ _10936_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10390_/X sky130_fd_sc_hd__and2_1
XFILLER_109_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08191__A _08191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_86_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10986_/CLK sky130_fd_sc_hd__clkbuf_16
X_09049_ _10934_/Q _10394_/C _10430_/B _10950_/Q vssd1 vssd1 vccd1 vccd1 _09049_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07519__B _07519_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09226__S _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input10_A io_wbs_m2s_addr[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10486__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10751_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10865_/CLK sky130_fd_sc_hd__clkbuf_16
X_10726_ _10940_/CLK _10726_/D vssd1 vssd1 vccd1 vccd1 _10726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 _10977_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_146_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10657_ _10657_/CLK _10657_/D vssd1 vssd1 vccd1 vccd1 _10657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10588_ _10968_/CLK _10588_/D vssd1 vssd1 vccd1 vccd1 _10588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07164__B _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ _06758_/A _06776_/A vssd1 vssd1 vccd1 vccd1 _06771_/B sky130_fd_sc_hd__and2_1
XFILLER_36_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05701_ _08206_/A vssd1 vssd1 vccd1 vccd1 _05702_/A sky130_fd_sc_hd__clkinv_2
XFILLER_36_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06681_ _06681_/A _06681_/B vssd1 vssd1 vccd1 vccd1 _06947_/B sky130_fd_sc_hd__or2_1
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08420_ _06143_/X _08419_/B _08419_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10729_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05632_ _10547_/Q _05636_/A vssd1 vssd1 vccd1 vccd1 _05632_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08276__A _08278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07180__A _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08351_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08351_/Y sky130_fd_sc_hd__nand2_1
X_05563_ _10570_/Q _10571_/Q _05576_/A vssd1 vssd1 vccd1 vccd1 _05566_/A sky130_fd_sc_hd__or3_1
XFILLER_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07302_ _07302_/A _07302_/B vssd1 vssd1 vccd1 vccd1 _07307_/B sky130_fd_sc_hd__xor2_2
XFILLER_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08282_ _08282_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08282_/X sky130_fd_sc_hd__or2_1
X_05494_ _05383_/X _05489_/X _05490_/X _05461_/D vssd1 vssd1 vccd1 vccd1 _10549_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_07233_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07236_/A sky130_fd_sc_hd__xnor2_2
XFILLER_149_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07164_ _07166_/A _07164_/B vssd1 vssd1 vccd1 vccd1 _07196_/A sky130_fd_sc_hd__nand2_2
XFILLER_145_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06115_ _06115_/A _06115_/B vssd1 vssd1 vccd1 vccd1 _08036_/B sky130_fd_sc_hd__nor2_1
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07095_ _07284_/A _07095_/B vssd1 vssd1 vccd1 vccd1 _07096_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06046_ _10663_/Q vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08358__B1 _08092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input2_A io_qei_ch_a vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ _09805_/A _09919_/B vssd1 vssd1 vccd1 vccd1 _09856_/C sky130_fd_sc_hd__and2_1
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07997_ _06206_/X _07987_/X _07996_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10663_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06948_ _06948_/A _06948_/B vssd1 vssd1 vccd1 vccd1 _07659_/A sky130_fd_sc_hd__and2_1
X_09736_ _09931_/A _09736_/B _09737_/A _09802_/C vssd1 vssd1 vccd1 vccd1 _09870_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10468__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__nor2_1
X_06879_ _06881_/A _06881_/B _06878_/Y vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__o21a_1
XFILLER_43_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08618_ _08600_/X _08597_/B _08623_/D _10789_/Q vssd1 vssd1 vccd1 vccd1 _08619_/C
+ sky130_fd_sc_hd__a31o_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09598_ _09560_/A _09560_/B _09597_/X vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__o21ai_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08549_/A vssd1 vssd1 vccd1 vccd1 _10770_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06418__B _07061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05647__A1 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10511_ _10529_/A vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10373_ _10412_/A vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09745__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09480__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05513__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09077__A1 _08119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10709_ _10709_/CLK _10709_/D vssd1 vssd1 vccd1 vccd1 _10709_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06063__A1 _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06998__B _07008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07920_ _10612_/Q _07906_/X _07910_/X _07919_/Y vssd1 vssd1 vccd1 vccd1 _07921_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07851_ _10577_/Q vssd1 vssd1 vccd1 vccd1 _07866_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06802_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _06821_/A sky130_fd_sc_hd__xor2_1
XFILLER_96_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput2 io_qei_ch_a vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_8
X_07782_ _07782_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _07786_/A sky130_fd_sc_hd__xnor2_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _09520_/B _09520_/C _09520_/A vssd1 vssd1 vccd1 vccd1 _09522_/B sky130_fd_sc_hd__o21ai_1
XFILLER_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06733_ _06752_/B _06752_/C vssd1 vssd1 vccd1 vccd1 _06745_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06118__A2 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09488_/A sky130_fd_sc_hd__and2_1
XFILLER_24_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06664_ _06695_/A _06695_/B _06661_/A vssd1 vssd1 vccd1 vccd1 _06665_/B sky130_fd_sc_hd__a21oi_2
XFILLER_36_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08403_ _08408_/A _10758_/Q vssd1 vssd1 vccd1 vccd1 _08403_/X sky130_fd_sc_hd__or2_1
X_05615_ _10555_/Q _05664_/A vssd1 vssd1 vccd1 vccd1 _05615_/Y sky130_fd_sc_hd__xnor2_1
X_09383_ _09383_/A vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__clkbuf_2
X_06595_ _06607_/B _06607_/C _06607_/A vssd1 vssd1 vccd1 vccd1 _06599_/B sky130_fd_sc_hd__a21boi_1
XFILLER_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08334_ _08027_/A _08058_/X _08333_/X _06011_/X vssd1 vssd1 vccd1 vccd1 _08334_/X
+ sky130_fd_sc_hd__o211a_1
X_05546_ _05652_/A _05546_/B vssd1 vssd1 vccd1 vccd1 _05637_/B sky130_fd_sc_hd__or2_1
XFILLER_138_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08265_ _08267_/A _08277_/C vssd1 vssd1 vccd1 vccd1 _08276_/B sky130_fd_sc_hd__and2_1
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05477_ _05643_/A vssd1 vssd1 vccd1 vccd1 _05912_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_119_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07216_ _07222_/A _07216_/B vssd1 vssd1 vccd1 vccd1 _07217_/B sky130_fd_sc_hd__nand2_1
XFILLER_137_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08196_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08196_/X sky130_fd_sc_hd__and2_1
XFILLER_119_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07147_ _07147_/A _07147_/B vssd1 vssd1 vccd1 vccd1 _07309_/B sky130_fd_sc_hd__xor2_1
XFILLER_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ _07167_/B vssd1 vssd1 vccd1 vccd1 _07163_/B sky130_fd_sc_hd__inv_2
XFILLER_156_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06029_ _10412_/A _08157_/A _10351_/A _10578_/Q vssd1 vssd1 vccd1 vccd1 _06029_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10504__A _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08200__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__B _10935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09719_ _09599_/A _09760_/B _09903_/A _09805_/A vssd1 vssd1 vccd1 vccd1 _09719_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08644__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _06202_/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10425_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__09475__A _09475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10356_ _10351_/X _06752_/B _10355_/X _10923_/Q vssd1 vssd1 vccd1 vccd1 _10923_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10287_ _10287_/A _10287_/B _10287_/C _10287_/D vssd1 vssd1 vccd1 vccd1 _10289_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09298__B2 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05400_ _05400_/A _05400_/B vssd1 vssd1 vccd1 vccd1 _05485_/A sky130_fd_sc_hd__xnor2_2
X_06380_ _06896_/A _06381_/C vssd1 vssd1 vccd1 vccd1 _06394_/A sky130_fd_sc_hd__nor2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05331_ _10673_/Q vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__clkinv_2
XFILLER_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _10369_/A _08971_/B _08416_/A _10583_/Q vssd1 vssd1 vccd1 vccd1 _08124_/A
+ sky130_fd_sc_hd__a31o_2
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07001_ _07574_/A _07439_/A vssd1 vssd1 vccd1 vccd1 _07573_/C sky130_fd_sc_hd__nand2_2
XFILLER_115_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08952_ _10341_/B _09016_/B vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__nor2_1
XFILLER_130_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07903_ _07903_/A vssd1 vssd1 vccd1 vccd1 _07903_/Y sky130_fd_sc_hd__inv_2
X_08883_ _08883_/A _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08883_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07834_ _07827_/X _05462_/C _07823_/X _07833_/Y vssd1 vssd1 vccd1 vccd1 _10621_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07765_ _10504_/A _07767_/B _06860_/B _06859_/A vssd1 vssd1 vccd1 vccd1 _07769_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_38_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09504_ _09676_/B _09444_/A _09444_/B _09361_/A vssd1 vssd1 vccd1 vccd1 _09507_/A
+ sky130_fd_sc_hd__a31o_2
X_06716_ _06876_/B _06876_/A vssd1 vssd1 vccd1 vccd1 _07794_/A sky130_fd_sc_hd__or2b_1
X_07696_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _07696_/X sky130_fd_sc_hd__or2b_1
XFILLER_53_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09435_ _09471_/A _09435_/B vssd1 vssd1 vccd1 vccd1 _09477_/B sky130_fd_sc_hd__xnor2_2
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06647_ _06647_/A _06647_/B vssd1 vssd1 vccd1 vccd1 _06648_/B sky130_fd_sc_hd__or2_1
XFILLER_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08249__C1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ _09676_/B _09444_/A _09444_/B _09361_/A _09506_/B vssd1 vssd1 vccd1 vccd1
+ _09546_/B sky130_fd_sc_hd__a311o_1
X_06578_ _06578_/A _06578_/B _06578_/C vssd1 vssd1 vccd1 vccd1 _06581_/B sky130_fd_sc_hd__and3_1
X_08317_ _08317_/A _08317_/B vssd1 vssd1 vccd1 vccd1 _08317_/Y sky130_fd_sc_hd__nand2_1
X_05529_ _10572_/Q vssd1 vssd1 vccd1 vccd1 _05564_/A sky130_fd_sc_hd__inv_2
X_09297_ _10679_/Q _09296_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__mux2_1
XFILLER_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08248_ _08248_/A vssd1 vssd1 vccd1 vccd1 _08248_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_126_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08179_ _08191_/B _08178_/X _06117_/D vssd1 vssd1 vccd1 vccd1 _08179_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_134_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10210_ _10202_/X _10203_/X _10208_/X _09480_/X vssd1 vssd1 vccd1 vccd1 _10210_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_106_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10141_ _10484_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10142_/B sky130_fd_sc_hd__nand2_1
XFILLER_106_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05328__A _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__and2_1
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08724__B1 _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10974_ _10976_/CLK _10974_/D vssd1 vssd1 vccd1 vccd1 _10974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05998__A _09090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ _10408_/A vssd1 vssd1 vccd1 vccd1 _10408_/X sky130_fd_sc_hd__clkbuf_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10339_ _10337_/Y _10338_/X _07539_/A _10192_/X vssd1 vssd1 vccd1 vccd1 _10913_/D
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05880_ _10655_/Q _10654_/Q _06038_/A _05906_/A vssd1 vssd1 vccd1 vccd1 _05900_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07550_ _07743_/B _07550_/B vssd1 vssd1 vccd1 vccd1 _07586_/A sky130_fd_sc_hd__or2_1
XFILLER_93_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06501_ _06517_/A _06489_/B _06506_/B _06758_/B vssd1 vssd1 vccd1 vccd1 _06503_/A
+ sky130_fd_sc_hd__a22oi_1
X_07481_ _07489_/A _07481_/B vssd1 vssd1 vccd1 vccd1 _07482_/B sky130_fd_sc_hd__and2_1
XFILLER_62_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09220_ _08233_/A _07882_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06432_ _06645_/A _06433_/B vssd1 vssd1 vccd1 vccd1 _06434_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08284__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09151_ _10809_/Q _08985_/X _08988_/X _10722_/Q _09150_/X vssd1 vssd1 vccd1 vccd1
+ _09151_/X sky130_fd_sc_hd__a221o_1
X_06363_ _06576_/B vssd1 vssd1 vccd1 vccd1 _06460_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08102_ _08098_/A _08098_/B _05728_/X vssd1 vssd1 vccd1 vccd1 _08102_/Y sky130_fd_sc_hd__o21ai_1
X_05314_ _10677_/Q _10676_/Q _05831_/B vssd1 vssd1 vccd1 vccd1 _05827_/A sky130_fd_sc_hd__or3_1
XFILLER_159_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09082_ _10969_/Q vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06294_ _10904_/Q vssd1 vssd1 vccd1 vccd1 _09356_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08033_ input39/X _07985_/B _08032_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10678_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06251__B _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09984_ _09918_/A _09918_/B _09916_/A vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__a21oi_2
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08935_ _08935_/A _10831_/Q vssd1 vssd1 vccd1 vccd1 _08936_/A sky130_fd_sc_hd__and2_1
XFILLER_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08866_ _08866_/A _08866_/B _08870_/D vssd1 vssd1 vccd1 vccd1 _08866_/X sky130_fd_sc_hd__and3_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08182__A1 _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07817_ _10868_/Q _07824_/B vssd1 vssd1 vccd1 vccd1 _07817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08797_ _10813_/Q _08815_/B _08792_/Y vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__a21bo_1
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07748_ _07748_/A _07748_/B vssd1 vssd1 vccd1 vccd1 _07750_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07679_ _09303_/B _07249_/B _07519_/B vssd1 vssd1 vccd1 vccd1 _07680_/B sky130_fd_sc_hd__a21bo_1
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09418_ _09418_/A vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__clkbuf_2
X_10690_ _10693_/CLK _10690_/D vssd1 vssd1 vccd1 vccd1 _10690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09349_ _07013_/A _10891_/Q vssd1 vssd1 vccd1 vccd1 _09372_/B sky130_fd_sc_hd__and2b_1
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06248__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input40_A io_wbs_m2s_data[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _10124_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__xnor2_1
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10055_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10091_/B sky130_fd_sc_hd__nand2_1
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08369__A _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10314__A_N _10944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10957_ _10958_/CLK _10957_/D vssd1 vssd1 vccd1 vccd1 _10957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10888_ _10980_/CLK _10888_/D vssd1 vssd1 vccd1 vccd1 _10888_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _07098_/A _07102_/A vssd1 vssd1 vccd1 vccd1 _07747_/B sky130_fd_sc_hd__or2_2
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08720_ _08840_/B vssd1 vssd1 vccd1 vccd1 _08888_/B sky130_fd_sc_hd__clkbuf_2
X_05932_ _08224_/A _05870_/X _05866_/X _08233_/A _05931_/X vssd1 vssd1 vccd1 vccd1
+ _05932_/X sky130_fd_sc_hd__o221a_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08651_ _10798_/Q vssd1 vssd1 vccd1 vccd1 _08651_/Y sky130_fd_sc_hd__inv_2
X_05863_ _05863_/A _05863_/B vssd1 vssd1 vccd1 vccd1 _05863_/X sky130_fd_sc_hd__and2_1
XFILLER_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07602_ _07502_/A _07502_/B _07455_/A vssd1 vssd1 vccd1 vccd1 _07711_/B sky130_fd_sc_hd__o21ai_4
X_08582_ _10780_/Q _08585_/C vssd1 vssd1 vccd1 vccd1 _08583_/B sky130_fd_sc_hd__and2_1
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05794_ _05794_/A _05794_/B vssd1 vssd1 vccd1 vccd1 _05794_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07533_ _07623_/A _07622_/B vssd1 vssd1 vccd1 vccd1 _07617_/B sky130_fd_sc_hd__or2_1
XFILLER_35_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07464_ _07464_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _07466_/B sky130_fd_sc_hd__nor2_1
XFILLER_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06415_ _10922_/Q _07083_/A vssd1 vssd1 vccd1 vccd1 _06416_/B sky130_fd_sc_hd__nand2_1
X_09203_ _09203_/A vssd1 vssd1 vccd1 vccd1 _09203_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_33_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07395_ _07393_/Y _07394_/X _07386_/B vssd1 vssd1 vccd1 vccd1 _07594_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08219__A2 _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05788__D _05802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ _09114_/X _09133_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06346_ _06346_/A _06346_/B vssd1 vssd1 vccd1 vccd1 _06561_/C sky130_fd_sc_hd__nand2_2
XANTENNA__07978__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09065_ _06038_/X _08995_/X _09064_/X _08981_/A vssd1 vssd1 vccd1 vccd1 _09065_/X
+ sky130_fd_sc_hd__a211o_1
X_06277_ _10898_/Q vssd1 vssd1 vccd1 vccd1 _07102_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_162_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08016_ _08289_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08016_/X sky130_fd_sc_hd__or2_1
XFILLER_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09967_ _09967_/A _09967_/B vssd1 vssd1 vccd1 vccd1 _09967_/Y sky130_fd_sc_hd__xnor2_1
X_08918_ hold9/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07805__B _10117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09898_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _09899_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08189__A _08191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08849_ _08846_/X _08848_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10819_/D sky130_fd_sc_hd__a21oi_1
XFILLER_40_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10811_ _10942_/CLK _10811_/D vssd1 vssd1 vccd1 vccd1 _10811_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10742_ _10776_/CLK _10742_/D vssd1 vssd1 vccd1 vccd1 _10742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10673_ _10674_/CLK _10673_/D vssd1 vssd1 vccd1 vccd1 _10673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09407__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06172__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10107_ _10107_/A _10107_/B vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__xor2_4
XFILLER_122_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10038_ _10039_/A _10039_/B vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06200_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06200_/X sky130_fd_sc_hd__buf_2
XFILLER_158_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07180_ _07197_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07181_/C sky130_fd_sc_hd__nand2_1
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06131_ _06204_/B vssd1 vssd1 vccd1 vccd1 _06131_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06062_ _08282_/A _05851_/A _05388_/A _05726_/A _06061_/X vssd1 vssd1 vccd1 vccd1
+ _06062_/X sky130_fd_sc_hd__a221o_1
XFILLER_172_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07906__A _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09821_ _09754_/A _09754_/B _09757_/B vssd1 vssd1 vccd1 vccd1 _09822_/B sky130_fd_sc_hd__o21ba_1
XFILLER_141_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09752_ _09684_/A _09683_/B _09961_/A vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__a21o_1
X_06964_ _07662_/A vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__buf_2
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08703_ _08709_/A _08704_/B _08704_/C vssd1 vssd1 vccd1 vccd1 _08705_/B sky130_fd_sc_hd__o21a_1
XFILLER_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05915_ _05408_/Y _05912_/B _05813_/X _05914_/X vssd1 vssd1 vccd1 vccd1 _05915_/X
+ sky130_fd_sc_hd__a31o_1
X_09683_ _10066_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06895_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _06896_/B sky130_fd_sc_hd__nor2_1
XFILLER_27_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05846_ _10671_/Q vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__buf_2
X_08634_ _08638_/C _08634_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _08635_/A sky130_fd_sc_hd__and3b_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10930_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_81_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05777_ _06113_/A _10570_/Q _10569_/Q _05766_/Y vssd1 vssd1 vccd1 vccd1 _05785_/A
+ sky130_fd_sc_hd__o22a_1
X_08565_ _10251_/S _10775_/Q _08565_/C vssd1 vssd1 vccd1 vccd1 _08565_/X sky130_fd_sc_hd__and3_1
XFILLER_70_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07516_ _07516_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__and2_1
X_08496_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08496_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__06257__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07447_ _07447_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07448_/B sky130_fd_sc_hd__or2_1
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07378_ _07728_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07378_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06329_ _10913_/Q vssd1 vssd1 vccd1 vccd1 _07112_/A sky130_fd_sc_hd__buf_2
X_09117_ _10939_/Q _09008_/X _09116_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09117_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_109_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08073__B1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09048_ _10369_/B vssd1 vssd1 vccd1 vccd1 _10394_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_136_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10242__A _10937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06167__A input45/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10725_ _10940_/CLK _10725_/D vssd1 vssd1 vccd1 vccd1 _10725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10656_ _10657_/CLK _10656_/D vssd1 vssd1 vccd1 vccd1 _10656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10587_ _10968_/CLK _10587_/D vssd1 vssd1 vccd1 vccd1 _10587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07726__A _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05700_ _10695_/Q vssd1 vssd1 vccd1 vccd1 _08206_/A sky130_fd_sc_hd__clkbuf_2
X_06680_ _06680_/A _06680_/B vssd1 vssd1 vccd1 vccd1 _06681_/B sky130_fd_sc_hd__and2_1
XFILLER_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08557__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05631_ _10687_/Q _05631_/B vssd1 vssd1 vccd1 vccd1 _05631_/X sky130_fd_sc_hd__or2_1
X_08350_ _08350_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08350_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05562_ _10569_/Q _10568_/Q _05769_/A _05582_/B vssd1 vssd1 vccd1 vccd1 _05576_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA_clkbuf_leaf_43_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07301_ _07301_/A _07344_/A vssd1 vssd1 vccd1 vccd1 _07302_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08281_ _08263_/X _08276_/Y _08295_/C _08280_/X _08062_/X vssd1 vssd1 vccd1 vccd1
+ _08281_/X sky130_fd_sc_hd__o32a_1
XFILLER_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05493_ _05385_/Y _05489_/X _05490_/X _05462_/A vssd1 vssd1 vccd1 vccd1 _10548_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07232_ _07232_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__xnor2_2
XFILLER_20_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07163_ _07415_/A _07163_/B _07186_/C vssd1 vssd1 vccd1 vccd1 _07193_/A sky130_fd_sc_hd__or3_2
XANTENNA__10972__D _10972_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06114_ _08351_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _06115_/B sky130_fd_sc_hd__or2_2
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10401__A2 _10719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07094_ _07284_/A _07095_/B vssd1 vssd1 vccd1 vccd1 _07363_/C sky130_fd_sc_hd__or2_1
XFILLER_160_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06045_ _06045_/A _06045_/B vssd1 vssd1 vccd1 vccd1 _06045_/X sky130_fd_sc_hd__or2_1
XANTENNA__06081__A2 _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08358__A1 _05528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09804_ _09870_/B _09804_/B vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__and2b_1
XFILLER_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07996_ _08209_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _07996_/X sky130_fd_sc_hd__or2_1
XFILLER_75_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09735_ _09735_/A _09735_/B vssd1 vssd1 vccd1 vccd1 _09802_/C sky130_fd_sc_hd__xor2_2
XFILLER_28_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06947_ _06947_/A _06947_/B vssd1 vssd1 vccd1 vccd1 _06948_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09666_ _09621_/A _09621_/B _09624_/A vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__o21a_1
X_06878_ _06878_/A _06878_/B vssd1 vssd1 vccd1 vccd1 _06878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08617_ _10789_/Q _08617_/B _08623_/D vssd1 vssd1 vccd1 vccd1 _08617_/X sky130_fd_sc_hd__and3_1
X_05829_ _05318_/A _05831_/C _05827_/Y _08032_/A vssd1 vssd1 vccd1 vccd1 _05829_/X
+ sky130_fd_sc_hd__o22a_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09597_ _09597_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__or2_1
XFILLER_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08580_/B _08548_/B _08553_/B vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__and3_1
XFILLER_168_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08479_ _10780_/Q _10743_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__mux2_1
XFILLER_51_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10510_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10510_/X sky130_fd_sc_hd__or2_1
XFILLER_156_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _10441_/A vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10372_ _06124_/A _10371_/X _10408_/A vssd1 vssd1 vccd1 vccd1 _10372_/X sky130_fd_sc_hd__a21bo_1
XFILLER_163_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10708_ _10859_/CLK _10708_/D vssd1 vssd1 vccd1 vccd1 _10708_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10639_ _10640_/CLK _10639_/D vssd1 vssd1 vccd1 vccd1 _10639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06063__A2 _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07850_ _07850_/A vssd1 vssd1 vccd1 vccd1 _07850_/X sky130_fd_sc_hd__buf_4
XFILLER_96_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_70_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10858_/CLK sky130_fd_sc_hd__clkbuf_16
X_06801_ _10510_/A _06842_/A vssd1 vssd1 vccd1 vccd1 _07774_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07781_ _10502_/A _06857_/B _07780_/X _07635_/A vssd1 vssd1 vccd1 vccd1 _07782_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 io_qei_ch_b vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_49_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09520_ _09520_/A _09520_/B _09520_/C vssd1 vssd1 vccd1 vccd1 _09563_/B sky130_fd_sc_hd__or3_1
X_06732_ _06732_/A _06732_/B vssd1 vssd1 vccd1 vccd1 _06752_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08287__A _08287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09451_ _09489_/A _09451_/B _09579_/A vssd1 vssd1 vccd1 vccd1 _09456_/A sky130_fd_sc_hd__and3_1
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06663_ _06663_/A _06663_/B vssd1 vssd1 vccd1 vccd1 _06695_/B sky130_fd_sc_hd__xnor2_2
XFILLER_51_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_85_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10984_/CLK sky130_fd_sc_hd__clkbuf_16
X_08402_ _08397_/X _10741_/Q _08394_/X _08401_/X vssd1 vssd1 vccd1 vccd1 _10723_/D
+ sky130_fd_sc_hd__o211a_1
X_05614_ _10554_/Q _05663_/B vssd1 vssd1 vccd1 vccd1 _05664_/A sky130_fd_sc_hd__nor2_1
XFILLER_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09382_ _09431_/A _09431_/B vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__xnor2_1
X_06594_ _06594_/A _06594_/B _06579_/Y vssd1 vssd1 vccd1 vccd1 _06607_/A sky130_fd_sc_hd__or3b_1
XFILLER_40_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08333_ _08333_/A _08333_/B _08038_/A vssd1 vssd1 vccd1 vccd1 _08333_/X sky130_fd_sc_hd__or3b_1
X_05545_ _05652_/B _05652_/C vssd1 vssd1 vccd1 vccd1 _05546_/B sky130_fd_sc_hd__nor2_1
X_08264_ _08277_/B vssd1 vssd1 vccd1 vccd1 _08267_/A sky130_fd_sc_hd__clkbuf_2
X_05476_ hold10/X _05471_/X _05474_/Y _05475_/X vssd1 vssd1 vccd1 vccd1 _10541_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07215_ _07248_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07250_/A sky130_fd_sc_hd__nand2_2
XFILLER_165_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08195_ _08196_/A _08196_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__nor2_1
XFILLER_119_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07146_ _07148_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07309_/A sky130_fd_sc_hd__nand2_1
XFILLER_146_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10776_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__06054__A2 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ _07151_/A _07390_/B _07375_/A vssd1 vssd1 vccd1 vccd1 _07091_/B sky130_fd_sc_hd__a21boi_1
XFILLER_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06028_ _08489_/A vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__buf_4
XFILLER_105_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_38_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10864_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07979_ _07979_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07979_/X sky130_fd_sc_hd__or2_1
XFILLER_28_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09718_ _09930_/B _09903_/A vssd1 vssd1 vccd1 vccd1 _09718_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09649_ _09619_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09649_/X sky130_fd_sc_hd__and2b_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08082__D _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _10945_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10424_/X sky130_fd_sc_hd__and2_1
XFILLER_171_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08660__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10377__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10355_ _10355_/A vssd1 vssd1 vccd1 vccd1 _10355_/X sky130_fd_sc_hd__buf_2
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10301_/A _10300_/A vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10430__A _10495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05330_ _10641_/Q vssd1 vssd1 vccd1 vccd1 _07907_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07000_ _09920_/B _07000_/B vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__xnor2_1
XFILLER_174_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06036__A2 _08119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08951_ _09126_/A _09142_/D vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__or2_1
XFILLER_131_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07902_ _07916_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _10639_/D sky130_fd_sc_hd__nor2_1
XFILLER_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08882_ _10824_/Q _08888_/B vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__xor2_1
XFILLER_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07833_ _06160_/A _07828_/X _07829_/X _07831_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07833_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07764_ _07764_/A _07764_/B vssd1 vssd1 vccd1 vccd1 _07803_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09503_ _09448_/A _09879_/B _09678_/A vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__o21ai_4
XFILLER_71_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06715_ _06715_/A _06721_/A vssd1 vssd1 vccd1 vccd1 _06876_/A sky130_fd_sc_hd__xnor2_1
XFILLER_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08497__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07695_ _07693_/A _07693_/B _09576_/A vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__a21bo_2
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _10066_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09435_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06646_ _06646_/A _06646_/B vssd1 vssd1 vccd1 vccd1 _06647_/B sky130_fd_sc_hd__and2_1
XFILLER_52_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08249__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09365_ _10887_/Q _10903_/Q vssd1 vssd1 vccd1 vccd1 _09506_/B sky130_fd_sc_hd__and2b_1
X_06577_ _06578_/A _06578_/B _06578_/C vssd1 vssd1 vccd1 vccd1 _06581_/C sky130_fd_sc_hd__a21oi_1
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08316_ _08305_/A _08315_/C _08317_/A vssd1 vssd1 vccd1 vccd1 _08316_/Y sky130_fd_sc_hd__a21oi_1
X_05528_ _05528_/A vssd1 vssd1 vccd1 vccd1 _05528_/X sky130_fd_sc_hd__clkbuf_4
X_09296_ _06115_/A _10647_/Q _09296_/S vssd1 vssd1 vccd1 vccd1 _09296_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08247_ _08243_/A _08251_/C _08246_/Y vssd1 vssd1 vccd1 vccd1 _08247_/Y sky130_fd_sc_hd__a21oi_1
X_05459_ _05453_/A _09107_/A _09078_/A _05455_/X _05458_/X vssd1 vssd1 vccd1 vccd1
+ _05459_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08480__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _08173_/A _08173_/B _08181_/A vssd1 vssd1 vccd1 vccd1 _08178_/X sky130_fd_sc_hd__a21o_1
X_07129_ _10985_/Q _07229_/B _07376_/A vssd1 vssd1 vccd1 vccd1 _07133_/B sky130_fd_sc_hd__a21boi_2
XFILLER_106_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10515__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _10482_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10142_/A sky130_fd_sc_hd__nand2_1
XFILLER_161_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10071_ _10482_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__and2_1
XFILLER_88_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10973_ _10978_/CLK _10973_/D vssd1 vssd1 vccd1 vccd1 _10973_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10407_ _10389_/X _10721_/Q _10405_/X _10406_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10940_/D sky130_fd_sc_hd__o221a_1
XFILLER_98_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10338_ _10336_/X _10332_/X _10333_/Y _09480_/X vssd1 vssd1 vccd1 vccd1 _10338_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__05777__A1 _06113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05777__B2 _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _10252_/A _10247_/A _10261_/A _10268_/Y vssd1 vssd1 vccd1 vccd1 _10287_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08176__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07518__A2 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06500_ _06502_/B vssd1 vssd1 vccd1 vccd1 _06758_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07480_ _07480_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__xnor2_1
XFILLER_35_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08565__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06431_ _06431_/A _06431_/B vssd1 vssd1 vccd1 vccd1 _06433_/B sky130_fd_sc_hd__xor2_1
XFILLER_22_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06362_ _06587_/A vssd1 vssd1 vccd1 vccd1 _06576_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09150_ _07979_/A _09123_/X _09127_/X _09149_/X vssd1 vssd1 vccd1 vccd1 _09150_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05313_ _05329_/A vssd1 vssd1 vccd1 vccd1 _05831_/B sky130_fd_sc_hd__clkbuf_2
X_08101_ _08097_/X _08099_/X _08100_/X vssd1 vssd1 vccd1 vccd1 _10684_/D sky130_fd_sc_hd__o21a_1
X_06293_ _06293_/A _06293_/B vssd1 vssd1 vccd1 vccd1 _06805_/A sky130_fd_sc_hd__nor2_2
X_09081_ _08974_/X _09077_/X _09078_/Y _09036_/X _09080_/X vssd1 vssd1 vccd1 vccd1
+ _09081_/X sky130_fd_sc_hd__a32o_1
X_08032_ _08032_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 io_wbs_m2s_we vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_4
XFILLER_116_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10980__D _10980_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10210__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05768__A1 _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09983_ _09983_/A _09983_/B vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__xor2_1
XFILLER_89_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05768__B2 _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ _08934_/A vssd1 vssd1 vccd1 vccd1 _10831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08706__A1 _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08167__C1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08865_ _10822_/Q _08865_/B vssd1 vssd1 vccd1 vccd1 _08870_/D sky130_fd_sc_hd__xor2_1
XFILLER_85_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07816_ _06255_/X _08994_/A _06257_/X _07815_/Y vssd1 vssd1 vccd1 vccd1 _10617_/D
+ sky130_fd_sc_hd__o211a_1
X_08796_ _10814_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08803_/D sky130_fd_sc_hd__xor2_1
XFILLER_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07747_ _07747_/A _07747_/B vssd1 vssd1 vccd1 vccd1 _07748_/A sky130_fd_sc_hd__nor2_1
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07678_ _07678_/A _09303_/B vssd1 vssd1 vccd1 vccd1 _07680_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09417_ _09417_/A _09810_/A vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__or2_1
X_06629_ _06800_/A _06719_/C vssd1 vssd1 vccd1 vccd1 _06630_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09348_ _10891_/Q _10907_/Q vssd1 vssd1 vccd1 vccd1 _09371_/A sky130_fd_sc_hd__and2b_1
XFILLER_138_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _09289_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09280_/A sky130_fd_sc_hd__and2_2
XFILLER_138_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09198__B2 _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__nand2_1
XFILLER_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input33_A io_wbs_m2s_data[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _10055_/A _10055_/B vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__or2_1
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10956_ _10958_/CLK _10956_/D vssd1 vssd1 vccd1 vccd1 _10956_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08385__A _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05802__A _05802_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10887_ _10980_/CLK _10887_/D vssd1 vssd1 vccd1 vccd1 _10887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07436__A1 _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07436__B2 _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07729__A _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09189__B2 _05877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ _10899_/Q vssd1 vssd1 vccd1 vccd1 _07098_/A sky130_fd_sc_hd__clkbuf_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05931_ _08218_/A _05872_/X _05870_/X _08224_/A _05930_/X vssd1 vssd1 vccd1 vccd1
+ _05931_/X sky130_fd_sc_hd__a221o_1
XFILLER_67_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08650_ _08650_/A vssd1 vssd1 vccd1 vccd1 _10797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05862_ _05350_/B _05854_/B _08244_/A vssd1 vssd1 vccd1 vccd1 _05863_/A sky130_fd_sc_hd__o21ai_1
XFILLER_67_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07601_ _07601_/A _07601_/B vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__xnor2_2
XFILLER_82_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08581_ _08581_/A vssd1 vssd1 vccd1 vccd1 _10779_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05793_ _05732_/B _05741_/Y _05742_/B vssd1 vssd1 vccd1 vccd1 _05794_/B sky130_fd_sc_hd__a21oi_1
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07532_ _07628_/A _07627_/B vssd1 vssd1 vccd1 vccd1 _07622_/B sky130_fd_sc_hd__or2_1
XANTENNA__06808__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10975__D _10975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07463_ _07473_/A _07463_/B vssd1 vssd1 vccd1 vccd1 _07464_/B sky130_fd_sc_hd__and2_1
XFILLER_50_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09202_ _09202_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _10849_/D sky130_fd_sc_hd__nor2_4
X_06414_ _10905_/Q vssd1 vssd1 vccd1 vccd1 _07083_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_167_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07394_ _07394_/A vssd1 vssd1 vccd1 vccd1 _07394_/X sky130_fd_sc_hd__buf_2
XFILLER_148_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _10940_/Q _09008_/X _09132_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09133_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06345_ _06343_/A _06736_/A _06371_/C vssd1 vssd1 vccd1 vccd1 _06346_/B sky130_fd_sc_hd__o21ai_1
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06276_ _06276_/A _06276_/B vssd1 vssd1 vccd1 vccd1 _06352_/A sky130_fd_sc_hd__nand2_2
X_09064_ _05462_/C _08978_/A _06129_/B _05728_/X _09179_/A vssd1 vssd1 vccd1 vccd1
+ _09064_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08015_ _08015_/A vssd1 vssd1 vccd1 vccd1 _08015_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_38_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _09893_/Y _09896_/B _09894_/A vssd1 vssd1 vccd1 vccd1 _09967_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08917_ _08814_/X _08915_/Y _08916_/X vssd1 vssd1 vccd1 vccd1 _10828_/D sky130_fd_sc_hd__o21a_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07805__C _10117_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09897_ _10877_/Q _09572_/X _09896_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10877_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08848_ input28/X _08672_/X _08674_/X _08847_/X vssd1 vssd1 vccd1 vccd1 _08848_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06166__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _06191_/X _08728_/X _08729_/X _08771_/A vssd1 vssd1 vccd1 vccd1 _08779_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _10942_/CLK _10810_/D vssd1 vssd1 vccd1 vccd1 _10810_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _10776_/CLK _10741_/D vssd1 vssd1 vccd1 vccd1 _10741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10672_ _10674_/CLK _10672_/D vssd1 vssd1 vccd1 vccd1 _10672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10106_ _10035_/A _10035_/B _10105_/X vssd1 vssd1 vccd1 vccd1 _10107_/B sky130_fd_sc_hd__a21o_2
XFILLER_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07715__C _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05770__A1_N _05767_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10037_ _10037_/A _10037_/B vssd1 vssd1 vccd1 vccd1 _10039_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06157__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10939_ _10940_/CLK _10939_/D vssd1 vssd1 vccd1 vccd1 _10939_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_143_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06130_ _06149_/A vssd1 vssd1 vccd1 vccd1 _06204_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_157_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06061_ _06061_/A _08000_/A vssd1 vssd1 vccd1 vccd1 _06061_/X sky130_fd_sc_hd__xor2_1
XFILLER_173_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08909__A1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09031__A0 _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09820_ _09820_/A _09820_/B vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06810__B _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09751_ _10066_/A vssd1 vssd1 vccd1 vccd1 _09961_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_113_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06963_ _07675_/A vssd1 vssd1 vccd1 vccd1 _07662_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_140_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10332__B _10946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ _08691_/B _08693_/B _08689_/Y vssd1 vssd1 vccd1 vccd1 _08704_/C sky130_fd_sc_hd__a21o_1
XFILLER_67_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05914_ _10681_/Q _05913_/Y _05814_/X vssd1 vssd1 vccd1 vccd1 _05914_/X sky130_fd_sc_hd__a21bo_1
XFILLER_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _09682_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06894_ _06894_/A _06894_/B vssd1 vssd1 vccd1 vccd1 _06899_/A sky130_fd_sc_hd__xor2_4
XFILLER_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08633_ _08633_/A vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__buf_4
X_05845_ _05845_/A _05941_/B vssd1 vssd1 vccd1 vccd1 _05940_/B sky130_fd_sc_hd__and2_1
XFILLER_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08564_ _10774_/Q _08559_/X _08562_/X _08563_/X vssd1 vssd1 vccd1 vccd1 _10774_/D
+ sky130_fd_sc_hd__o211a_1
X_05776_ _08297_/A _05772_/Y _05564_/A _06115_/A _05807_/A vssd1 vssd1 vccd1 vccd1
+ _05786_/C sky130_fd_sc_hd__o221a_1
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07515_ _07515_/A _07515_/B vssd1 vssd1 vccd1 vccd1 _07516_/B sky130_fd_sc_hd__or2_1
X_08495_ _10783_/Q _08491_/X _08494_/X _10746_/Q vssd1 vssd1 vccd1 vccd1 _10746_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07446_ _07714_/S _07445_/B _07445_/C vssd1 vssd1 vccd1 vccd1 _07447_/B sky130_fd_sc_hd__a21oi_1
XFILLER_168_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07377_ _07377_/A vssd1 vssd1 vccd1 vccd1 _07728_/A sky130_fd_sc_hd__buf_2
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09116_ _10955_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09116_/Y sky130_fd_sc_hd__nor2_1
X_06328_ _06288_/X _06851_/A _06851_/B _06850_/A vssd1 vssd1 vccd1 vccd1 _06342_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06084__B1 _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ _10432_/A _09142_/C _09142_/D _10341_/B vssd1 vssd1 vccd1 vccd1 _10369_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06259_ _10978_/Q vssd1 vssd1 vccd1 vccd1 _06436_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09477__A_N _09436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09949_ _09949_/A vssd1 vssd1 vccd1 vccd1 _09949_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07832__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09089__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08836__B1 _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ _10940_/CLK _10724_/D vssd1 vssd1 vccd1 vccd1 _10724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10655_ _10655_/CLK _10655_/D vssd1 vssd1 vccd1 vccd1 _10655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08064__A1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10586_ _10968_/CLK _10586_/D vssd1 vssd1 vccd1 vccd1 _10586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05527__A _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05630_ _05630_/A _05630_/B vssd1 vssd1 vccd1 vccd1 _05631_/B sky130_fd_sc_hd__and2_1
XFILLER_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05561_ _10566_/Q _05588_/A vssd1 vssd1 vccd1 vccd1 _05582_/B sky130_fd_sc_hd__or2_1
X_07300_ _07349_/B _07300_/B vssd1 vssd1 vccd1 vccd1 _07307_/A sky130_fd_sc_hd__or2_1
Xclkbuf_opt_2_1_clock clkbuf_opt_2_1_clock/A vssd1 vssd1 vccd1 vccd1 _10863_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_60_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08280_ _05851_/A _08235_/B _08278_/Y _08279_/X vssd1 vssd1 vccd1 vccd1 _08280_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05492_ _05389_/Y _05489_/X _05490_/X _05462_/B vssd1 vssd1 vccd1 vccd1 _10547_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_149_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07231_ _07231_/A _07231_/B vssd1 vssd1 vccd1 vccd1 _07258_/A sky130_fd_sc_hd__xnor2_1
XFILLER_30_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09252__A0 _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ _07211_/A _07166_/B vssd1 vssd1 vccd1 vccd1 _07186_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08055__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08055__B2 _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06113_ _06113_/A _08333_/A vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__nand2_1
XFILLER_161_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07093_ _07363_/B _07093_/B vssd1 vssd1 vccd1 vccd1 _07095_/B sky130_fd_sc_hd__nand2_1
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06044_ _05749_/A _10671_/Q _05408_/Y _08082_/D vssd1 vssd1 vccd1 vccd1 _06045_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07917__A _08462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10343__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09803_ _10069_/A _09802_/B _09930_/C _09932_/A vssd1 vssd1 vccd1 vccd1 _09804_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07995_ _07995_/A vssd1 vssd1 vccd1 vccd1 _08005_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09734_ _09734_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09735_/B sky130_fd_sc_hd__xnor2_2
XFILLER_68_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06946_ _06946_/A _06948_/A vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__xnor2_1
X_09665_ _09665_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__xor2_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06877_ _06878_/A _06878_/B vssd1 vssd1 vccd1 vccd1 _06881_/B sky130_fd_sc_hd__xnor2_2
XFILLER_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08616_ _08614_/Y _08612_/C _08623_/D _08617_/B _08630_/A vssd1 vssd1 vccd1 vccd1
+ _10788_/D sky130_fd_sc_hd__a221oi_1
X_05828_ _10678_/Q vssd1 vssd1 vccd1 vccd1 _08032_/A sky130_fd_sc_hd__inv_2
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__xnor2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ _08547_/A _08547_/B vssd1 vssd1 vccd1 vccd1 _08553_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05759_ _06061_/A vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__inv_2
XFILLER_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08478_ _08478_/A vssd1 vssd1 vccd1 vccd1 _10742_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08483__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07429_ _07429_/A _07429_/B vssd1 vssd1 vccd1 vccd1 _07430_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ _10950_/Q _10440_/B vssd1 vssd1 vccd1 vccd1 _10440_/X sky130_fd_sc_hd__or2_1
XFILLER_137_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10371_ _10371_/A vssd1 vssd1 vccd1 vccd1 _10371_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07827__A _07848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07562__A _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06178__A input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_7_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10859_/CLK _10707_/D vssd1 vssd1 vccd1 vccd1 _10707_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10638_ _10640_/CLK _10638_/D vssd1 vssd1 vccd1 vccd1 _10638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ _10855_/CLK _10569_/D vssd1 vssd1 vccd1 vccd1 _10569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_4_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10981_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06800_ _06800_/A vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_84_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07780_ _06855_/A _07780_/B _07780_/C vssd1 vssd1 vccd1 vccd1 _07780_/X sky130_fd_sc_hd__and3b_1
XFILLER_96_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput4 io_wbs_m2s_addr[0] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_6
X_06731_ _06731_/A _06731_/B vssd1 vssd1 vccd1 vccd1 _06752_/B sky130_fd_sc_hd__xnor2_4
XFILLER_49_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09450_ _09555_/A _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__and3_1
XFILLER_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06662_ _06692_/A _06692_/B _06621_/A vssd1 vssd1 vccd1 vccd1 _06663_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08401_ _08408_/A _10757_/Q vssd1 vssd1 vccd1 vccd1 _08401_/X sky130_fd_sc_hd__or2_1
X_05613_ _10694_/Q vssd1 vssd1 vccd1 vccd1 _05877_/A sky130_fd_sc_hd__buf_2
X_09381_ _09381_/A _10897_/Q vssd1 vssd1 vccd1 vccd1 _09431_/B sky130_fd_sc_hd__xor2_4
XFILLER_91_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06593_ _06593_/A _06593_/B _06593_/C vssd1 vssd1 vccd1 vccd1 _06607_/C sky130_fd_sc_hd__and3_1
XFILLER_101_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08332_ _08332_/A _08332_/B vssd1 vssd1 vccd1 vccd1 _08333_/B sky130_fd_sc_hd__and2_1
X_05544_ _05910_/B _05737_/B _05543_/Y vssd1 vssd1 vccd1 vccd1 _05652_/C sky130_fd_sc_hd__a21oi_1
XFILLER_20_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10983__D _10983_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08263_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08263_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05475_ _10648_/Q vssd1 vssd1 vccd1 vccd1 _05475_/X sky130_fd_sc_hd__buf_4
X_07214_ _07214_/A _07214_/B vssd1 vssd1 vccd1 vccd1 _07232_/A sky130_fd_sc_hd__and2_1
XANTENNA__08028__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09225__A0 _08242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08194_ _08190_/X _08192_/X _08193_/X vssd1 vssd1 vccd1 vccd1 _10693_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07145_ _07145_/A _07145_/B vssd1 vssd1 vccd1 vccd1 _07148_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07076_ _07137_/A _07076_/B vssd1 vssd1 vccd1 vccd1 _07375_/A sky130_fd_sc_hd__nand2_1
XFILLER_160_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06027_ _08201_/A _09403_/B vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__and2_1
XFILLER_160_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08200__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _06178_/X _07965_/X _07976_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10657_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09717_ _09717_/A vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06929_ _06937_/A _06937_/B _06928_/Y vssd1 vssd1 vccd1 vccd1 _06936_/B sky130_fd_sc_hd__a21o_2
XFILLER_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09648_ _09649_/B _09619_/A vssd1 vssd1 vccd1 vccd1 _09648_/X sky130_fd_sc_hd__or2b_1
XFILLER_76_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10423_ _10408_/X _10725_/Q _10421_/X _10422_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10944_/D sky130_fd_sc_hd__o221a_1
XFILLER_136_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10354_ _09634_/A _06732_/B _08494_/X _10922_/Q vssd1 vssd1 vccd1 vccd1 _10922_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10285_ _10957_/Q _10941_/Q vssd1 vssd1 vccd1 vccd1 _10300_/A sky130_fd_sc_hd__and2b_1
XANTENNA__08727__C1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09758__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08950_ _09142_/A _09142_/B vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__or2_1
XFILLER_142_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07901_ _10607_/Q _07888_/X _07892_/X _07900_/Y vssd1 vssd1 vccd1 vccd1 _07902_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_69_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _10823_/D sky130_fd_sc_hd__nor2_1
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07832_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07832_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08298__A _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07941__A0 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10978__D _10978_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ _07763_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07764_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ _09501_/B _09501_/C _09501_/A vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__a21o_1
X_06714_ _06722_/A _06714_/B vssd1 vssd1 vccd1 vccd1 _06721_/A sky130_fd_sc_hd__xnor2_1
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08280__A2_N _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07694_ _09575_/B _09575_/C _09575_/A vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10190__B_N _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07930__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06645_ _06645_/A _06645_/B vssd1 vssd1 vccd1 vccd1 _06648_/A sky130_fd_sc_hd__or2_1
XFILLER_80_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08249__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09364_ _09336_/A _09336_/B _09421_/B _09333_/A vssd1 vssd1 vccd1 vccd1 _09444_/B
+ sky130_fd_sc_hd__a211o_1
X_06576_ _10974_/Q _06576_/B _06951_/A vssd1 vssd1 vccd1 vccd1 _06578_/C sky130_fd_sc_hd__and3_1
XANTENNA__05450__A _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08315_ _08315_/A _08315_/B _08315_/C vssd1 vssd1 vccd1 vccd1 _08327_/B sky130_fd_sc_hd__and3_1
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05527_ _06115_/A vssd1 vssd1 vccd1 vccd1 _05528_/A sky130_fd_sc_hd__buf_2
X_09295_ _09295_/A vssd1 vssd1 vccd1 vccd1 _10864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06265__B _10898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05468__D1 _05467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _08243_/A _08251_/C _08067_/X vssd1 vssd1 vccd1 vccd1 _08246_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05458_ _05455_/X _09078_/A _05283_/Y _09020_/A _05457_/X vssd1 vssd1 vccd1 vccd1
+ _05458_/X sky130_fd_sc_hd__o221a_1
X_08177_ _08172_/X _08174_/X _08176_/X vssd1 vssd1 vccd1 vccd1 _10691_/D sky130_fd_sc_hd__o21a_1
XFILLER_118_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05389_ _05389_/A _05389_/B vssd1 vssd1 vccd1 vccd1 _05389_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07128_ _07137_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _07376_/A sky130_fd_sc_hd__nand2_1
XFILLER_137_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07059_ _07560_/A _07076_/B vssd1 vssd1 vccd1 vccd1 _07357_/C sky130_fd_sc_hd__nand2_1
XFILLER_121_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10531__A _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__A_N _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10972_ _10978_/CLK _10972_/D vssd1 vssd1 vccd1 vccd1 _10972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_opt_6_0_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 clkbuf_opt_6_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10406_ _06178_/X _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10406_/X sky130_fd_sc_hd__a21bo_1
XFILLER_171_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06191__A input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_84_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10980_/CLK sky130_fd_sc_hd__clkbuf_16
X_10337_ _10332_/X _10333_/Y _10336_/X vssd1 vssd1 vccd1 vccd1 _10337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09117__A1_N _10939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _10268_/A vssd1 vssd1 vccd1 vccd1 _10268_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10441__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10199_ _10197_/Y _10198_/Y _09757_/A vssd1 vssd1 vccd1 vccd1 _10199_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10160__B _10160_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06083__A2_N _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08479__A1 _10743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10782_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06430_ _06631_/A _06430_/B vssd1 vssd1 vccd1 vccd1 _06431_/B sky130_fd_sc_hd__or2_1
XFILLER_50_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06361_ _06281_/B _06359_/Y _06360_/X vssd1 vssd1 vccd1 vccd1 _06587_/A sky130_fd_sc_hd__o21a_1
XANTENNA__06085__B _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ _10531_/A _08047_/X _08052_/X _08098_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08100_/X sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_37_clock _10856_/CLK vssd1 vssd1 vccd1 vccd1 _10848_/CLK sky130_fd_sc_hd__clkbuf_16
X_05312_ _10675_/Q _05834_/A vssd1 vssd1 vccd1 vccd1 _05329_/A sky130_fd_sc_hd__or2_1
XFILLER_148_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09080_ _10718_/Q _09079_/X _09037_/Y _10805_/Q vssd1 vssd1 vccd1 vccd1 _09080_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06292_ _10927_/Q _06993_/A vssd1 vssd1 vccd1 vccd1 _06293_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08031_ input37/X _07985_/B _08029_/Y _08030_/X vssd1 vssd1 vccd1 vccd1 _10677_/D
+ sky130_fd_sc_hd__o211a_1
Xinput40 io_wbs_m2s_data[31] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_6
XFILLER_156_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 reset vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_6
XFILLER_174_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07197__A _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09982_ _09982_/A _09982_/B vssd1 vssd1 vccd1 vccd1 _09983_/B sky130_fd_sc_hd__xnor2_1
XFILLER_107_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08933_ _08935_/A input2/X vssd1 vssd1 vccd1 vccd1 _08934_/A sky130_fd_sc_hd__and2_1
XFILLER_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08864_ _08881_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _10821_/D sky130_fd_sc_hd__nor2_1
XANTENNA__10351__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07815_ _06140_/A _06258_/X _07807_/X _07814_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07815_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_85_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08795_ _08793_/X _08794_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10813_/D sky130_fd_sc_hd__o21a_1
XFILLER_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07746_ _07746_/A _07746_/B vssd1 vssd1 vccd1 vccd1 _07755_/A sky130_fd_sc_hd__xnor2_1
XFILLER_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07677_ _07677_/A _07677_/B vssd1 vssd1 vccd1 vccd1 _07681_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09416_ _10964_/Q _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09427_/A sky130_fd_sc_hd__and3_1
XFILLER_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06628_ _06841_/A _06408_/B _06409_/C vssd1 vssd1 vccd1 vccd1 _06633_/A sky130_fd_sc_hd__a21boi_1
XFILLER_53_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_34_clock_A _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ _09863_/A _09797_/A vssd1 vssd1 vccd1 vccd1 _09372_/A sky130_fd_sc_hd__nand2_1
X_06559_ _06281_/B _06359_/Y _06360_/X _06558_/X _06502_/B vssd1 vssd1 vccd1 vccd1
+ _07676_/A sky130_fd_sc_hd__o2111a_1
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09278_ hold12/X _09274_/X _09275_/X _09277_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09279_/B sky130_fd_sc_hd__a32o_1
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08229_ _06117_/C _08074_/A _08228_/Y _08044_/A _08000_/A vssd1 vssd1 vccd1 vccd1
+ _08229_/X sky130_fd_sc_hd__a32o_1
XFILLER_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10526__A _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10122_ _10491_/A _10122_/B vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__nand2_1
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10053_ _10148_/A _10053_/B vssd1 vssd1 vccd1 vccd1 _10055_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A io_wbs_m2s_data[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07570__A _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10955_ _10958_/CLK _10955_/D vssd1 vssd1 vccd1 vccd1 _10955_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08330__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10886_ _10984_/CLK _10886_/D vssd1 vssd1 vccd1 vccd1 _10886_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05930_ _08206_/A _05876_/X _05872_/X _08224_/B _05929_/X vssd1 vssd1 vccd1 vccd1
+ _05930_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05861_ _10667_/Q vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07600_ _07598_/Y _07451_/B _07599_/X vssd1 vssd1 vccd1 vccd1 _07601_/B sky130_fd_sc_hd__o21a_1
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08580_ _08585_/C _08580_/B _08580_/C vssd1 vssd1 vccd1 vccd1 _08581_/A sky130_fd_sc_hd__and3b_1
X_05792_ _05747_/X _05761_/X _05749_/X vssd1 vssd1 vccd1 vccd1 _05792_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_82_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07531_ _07633_/A _07632_/B vssd1 vssd1 vccd1 vccd1 _07627_/B sky130_fd_sc_hd__or2_1
XFILLER_81_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ _07462_/A _07462_/B vssd1 vssd1 vccd1 vccd1 _07466_/A sky130_fd_sc_hd__nor2_1
X_09201_ _09112_/A _09197_/Y _09200_/X vssd1 vssd1 vccd1 vccd1 _09202_/B sky130_fd_sc_hd__a21oi_1
X_06413_ _06736_/A _06732_/A vssd1 vssd1 vccd1 vccd1 _06421_/A sky130_fd_sc_hd__nor2_1
XANTENNA__05686__B2 _05570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07393_ _07592_/A vssd1 vssd1 vccd1 vccd1 _07393_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09132_ _10956_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09132_/Y sky130_fd_sc_hd__nor2_1
X_06344_ _06352_/C vssd1 vssd1 vccd1 vccd1 _06736_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09063_ _10717_/Q _08999_/X _09037_/Y _10804_/Q vssd1 vssd1 vccd1 vccd1 _09063_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06275_ _06275_/A _06275_/B vssd1 vssd1 vccd1 vccd1 _06276_/B sky130_fd_sc_hd__or2_1
XANTENNA__10346__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08014_ input30/X _08002_/X _08013_/Y _08006_/X vssd1 vssd1 vccd1 vccd1 _10670_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07358__C _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09965_ _09965_/A _09964_/X vssd1 vssd1 vccd1 vccd1 _09967_/A sky130_fd_sc_hd__or2b_1
X_08916_ input37/X _08819_/X _08820_/X _10828_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08916_/X sky130_fd_sc_hd__o221a_1
XFILLER_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _09896_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__xnor2_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _10819_/Q vssd1 vssd1 vccd1 vccd1 _08847_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_40_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08778_ _08778_/A _08778_/B _08778_/C vssd1 vssd1 vccd1 vccd1 _08778_/X sky130_fd_sc_hd__and3_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07390__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _07729_/A _07729_/B vssd1 vssd1 vccd1 vccd1 _07730_/B sky130_fd_sc_hd__nand2_1
XFILLER_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _10776_/CLK _10740_/D vssd1 vssd1 vccd1 vccd1 _10740_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08863__A1 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10671_ _10671_/CLK _10671_/D vssd1 vssd1 vccd1 vccd1 _10671_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08933__B input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10422__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08379__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10186__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09040__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10105_ _10033_/B _10105_/B vssd1 vssd1 vccd1 vccd1 _10105_/X sky130_fd_sc_hd__and2b_1
XFILLER_110_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07715__D _07715_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10036_ _09961_/B _09962_/A _09961_/A vssd1 vssd1 vccd1 vccd1 _10037_/B sky130_fd_sc_hd__a21o_1
XFILLER_76_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08551__B1 _08462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05813__A _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10938_ _10940_/CLK _10938_/D vssd1 vssd1 vccd1 vccd1 _10938_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10869_ _10967_/CLK _10869_/D vssd1 vssd1 vccd1 vccd1 _10869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06060_ _08315_/A _08023_/A _08256_/A _05751_/Y _06059_/X vssd1 vssd1 vccd1 vccd1
+ _06070_/A sky130_fd_sc_hd__o221a_1
XFILLER_145_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07475__A _07728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08790__B1 _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _09815_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__or2_1
X_06962_ _07620_/A _06962_/B vssd1 vssd1 vccd1 vccd1 _06962_/X sky130_fd_sc_hd__and2_1
XFILLER_86_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08701_ _08701_/A _08732_/B vssd1 vssd1 vccd1 vccd1 _08704_/B sky130_fd_sc_hd__nor2_1
X_05913_ _05913_/A _05913_/B vssd1 vssd1 vccd1 vccd1 _05913_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09681_ _09681_/A _09802_/B vssd1 vssd1 vccd1 vccd1 _09684_/A sky130_fd_sc_hd__xor2_1
XFILLER_95_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06893_ _06893_/A _06893_/B vssd1 vssd1 vccd1 vccd1 _06894_/B sky130_fd_sc_hd__xor2_4
X_08632_ _08600_/X _08642_/D _10793_/Q vssd1 vssd1 vccd1 vccd1 _08634_/B sky130_fd_sc_hd__a21o_1
X_05844_ _05844_/A _05844_/B _05844_/C vssd1 vssd1 vccd1 vccd1 _05941_/B sky130_fd_sc_hd__or3_1
XFILLER_94_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06819__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10986__D _10986_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08563_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08563_/X sky130_fd_sc_hd__buf_4
X_05775_ _06113_/A _10570_/Q _10571_/Q _08355_/A vssd1 vssd1 vccd1 vccd1 _05807_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_42_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07514_ _07514_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__and2_1
XFILLER_81_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08494_ _10355_/A vssd1 vssd1 vccd1 vccd1 _08494_/X sky130_fd_sc_hd__buf_2
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07445_ _07714_/S _07445_/B _07445_/C vssd1 vssd1 vccd1 vccd1 _07447_/A sky130_fd_sc_hd__and3_1
XFILLER_23_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07376_ _07376_/A vssd1 vssd1 vccd1 vccd1 _07459_/B sky130_fd_sc_hd__clkbuf_2
X_09115_ _09194_/B vssd1 vssd1 vccd1 vccd1 _09164_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06327_ _10929_/Q _10912_/Q vssd1 vssd1 vccd1 vccd1 _06850_/A sky130_fd_sc_hd__and2_1
XFILLER_109_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09046_ _09930_/B vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__06084__B2 _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06258_ _07849_/A vssd1 vssd1 vccd1 vccd1 _06258_/X sky130_fd_sc_hd__buf_4
XFILLER_159_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09022__A1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06189_ _06189_/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08230__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08781__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ _09810_/B _09744_/B _09769_/B _10493_/A vssd1 vssd1 vccd1 vccd1 _09949_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_58_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09879_ _10129_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09880_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10274__B_N _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _10784_/CLK _10723_/D vssd1 vssd1 vccd1 vccd1 _10723_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10654_ _10654_/CLK _10654_/D vssd1 vssd1 vccd1 vccd1 _10654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10585_ _10968_/CLK _10585_/D vssd1 vssd1 vccd1 vccd1 _10585_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08064__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_3_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10841__CLK _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10019_ _10089_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10021_/B sky130_fd_sc_hd__and2_1
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05560_ _10565_/Q _10564_/Q _05593_/A vssd1 vssd1 vccd1 vccd1 _05588_/A sky130_fd_sc_hd__or3_1
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05491_ _05393_/B _05489_/X _05490_/X _05462_/C vssd1 vssd1 vccd1 vccd1 _10546_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_07230_ _07231_/A _07231_/B vssd1 vssd1 vccd1 vccd1 _07230_/X sky130_fd_sc_hd__and2_1
XFILLER_20_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07161_ _10982_/Q vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__inv_2
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06112_ _08339_/B _08332_/B vssd1 vssd1 vccd1 vccd1 _08333_/A sky130_fd_sc_hd__nor2_1
XFILLER_157_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09685__A _09689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07092_ _07402_/A _07091_/B _07091_/C vssd1 vssd1 vccd1 vccd1 _07093_/B sky130_fd_sc_hd__o21ai_1
XFILLER_106_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06043_ _10680_/Q vssd1 vssd1 vccd1 vccd1 _08082_/D sky130_fd_sc_hd__buf_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09802_ _09931_/A _09802_/B _09802_/C _09932_/A vssd1 vssd1 vccd1 vccd1 _09870_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07994_ _06202_/X _07987_/X _07991_/Y _07993_/X vssd1 vssd1 vccd1 vccd1 _10662_/D
+ sky130_fd_sc_hd__o211a_1
X_06945_ _06945_/A _06945_/B vssd1 vssd1 vccd1 vccd1 _06946_/A sky130_fd_sc_hd__nor2_1
X_09733_ _09371_/B _09733_/B vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__and2b_1
XFILLER_68_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09664_ _09779_/A _09779_/B vssd1 vssd1 vccd1 vccd1 _09728_/B sky130_fd_sc_hd__xor2_1
X_06876_ _06876_/A _06876_/B vssd1 vssd1 vccd1 vccd1 _06878_/B sky130_fd_sc_hd__xnor2_2
XFILLER_131_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05827_ _05827_/A _05831_/C vssd1 vssd1 vccd1 vccd1 _05827_/Y sky130_fd_sc_hd__nor2_1
X_08615_ _10788_/Q _10787_/Q _10786_/Q _10785_/Q vssd1 vssd1 vccd1 vccd1 _08623_/D
+ sky130_fd_sc_hd__and4_1
X_09595_ _09593_/Y _09595_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__and2b_1
XFILLER_55_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _10769_/Q _08543_/B _10770_/Q vssd1 vssd1 vccd1 vccd1 _08548_/B sky130_fd_sc_hd__a21o_1
X_05758_ _08224_/A vssd1 vssd1 vccd1 vccd1 _06061_/A sky130_fd_sc_hd__buf_2
XFILLER_23_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08477_ _08477_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08478_/A sky130_fd_sc_hd__or2_1
XFILLER_126_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05689_ _05528_/X _05564_/Y _05687_/B _08350_/A _05688_/X vssd1 vssd1 vccd1 vccd1
+ _05689_/X sky130_fd_sc_hd__a221o_1
XFILLER_51_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07428_ _07428_/A _07428_/B _07428_/C vssd1 vssd1 vccd1 vccd1 _07429_/B sky130_fd_sc_hd__nand3_1
XFILLER_168_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07359_ _07359_/A _07359_/B vssd1 vssd1 vccd1 vccd1 _07407_/A sky130_fd_sc_hd__xnor2_1
XFILLER_137_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10370_ _10399_/A vssd1 vssd1 vccd1 vccd1 _10371_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ _09716_/A vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__buf_2
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08939__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09482__B2 _09406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _10860_/CLK _10706_/D vssd1 vssd1 vccd1 vccd1 _10706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10637_ _10666_/CLK _10637_/D vssd1 vssd1 vccd1 vccd1 _10637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10568_ _10855_/CLK _10568_/D vssd1 vssd1 vccd1 vccd1 _10568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08993__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10499_ _06124_/X _10496_/X _10497_/Y _10498_/X vssd1 vssd1 vccd1 vccd1 _10971_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10193__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06730_ _06730_/A _06730_/B _06730_/C vssd1 vssd1 vccd1 vccd1 _06731_/A sky130_fd_sc_hd__nand3_2
XFILLER_65_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 io_wbs_m2s_addr[10] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06661_ _06661_/A _06661_/B vssd1 vssd1 vccd1 vccd1 _06695_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08400_ _08397_/X _10740_/Q _08394_/X _08399_/X vssd1 vssd1 vccd1 vccd1 _10722_/D
+ sky130_fd_sc_hd__o211a_1
X_05612_ _05612_/A _05612_/B vssd1 vssd1 vccd1 vccd1 _05612_/X sky130_fd_sc_hd__and2_1
X_09380_ _09338_/X _10065_/C _10063_/B _10062_/A vssd1 vssd1 vccd1 vccd1 _09431_/A
+ sky130_fd_sc_hd__a31o_2
X_06592_ _06949_/B _06952_/A _06591_/Y vssd1 vssd1 vccd1 vccd1 _06593_/C sky130_fd_sc_hd__a21o_1
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08331_ _08157_/X _08326_/X _08329_/Y _08330_/X vssd1 vssd1 vccd1 vccd1 _10707_/D
+ sky130_fd_sc_hd__o31a_1
X_05543_ _05454_/A _10543_/Q _05641_/A vssd1 vssd1 vccd1 vccd1 _05543_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08262_ _08262_/A vssd1 vssd1 vccd1 vccd1 _10700_/D sky130_fd_sc_hd__clkbuf_1
X_05474_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05474_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_165_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07213_ _07186_/A _07125_/A _07222_/B _07211_/A vssd1 vssd1 vccd1 vccd1 _07214_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08028__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08193_ _06195_/X _08164_/X _08165_/X _08191_/A _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08193_/X sky130_fd_sc_hd__o221a_1
XFILLER_158_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07144_ _07144_/A _07144_/B vssd1 vssd1 vccd1 vccd1 _07148_/A sky130_fd_sc_hd__and2_1
XFILLER_134_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07075_ _07377_/A _07151_/A _07076_/B _07390_/B vssd1 vssd1 vccd1 vccd1 _07402_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06026_ _10581_/Q _10582_/Q vssd1 vssd1 vccd1 vccd1 _09403_/B sky130_fd_sc_hd__and2b_4
XFILLER_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07977_ _07977_/A vssd1 vssd1 vccd1 vccd1 _07977_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09716_ _09716_/A _09760_/B vssd1 vssd1 vccd1 vccd1 _09716_/Y sky130_fd_sc_hd__nand2_1
X_06928_ _06928_/A _06928_/B vssd1 vssd1 vccd1 vccd1 _06928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09647_ _09647_/A _09647_/B vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__xnor2_1
XFILLER_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06859_ _06859_/A _06859_/B vssd1 vssd1 vccd1 vccd1 _06860_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09578_ _09563_/A _09563_/B _09564_/A vssd1 vssd1 vccd1 vccd1 _09623_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08494__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08529_ _06008_/A _10394_/B _08418_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _08529_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_169_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10529__A _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10422_ input20/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10422_/X sky130_fd_sc_hd__a21bo_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10353_ _10351_/X _06412_/A _10346_/X _10921_/Q vssd1 vssd1 vccd1 vccd1 _10921_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10284_ _10941_/Q _10957_/Q vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__and2b_1
XFILLER_97_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_opt_2_0_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_1_clock/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08669__A _10799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10174__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09963__A _09964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07900_ _07900_/A vssd1 vssd1 vccd1 vccd1 _07900_/Y sky130_fd_sc_hd__inv_2
X_08880_ _08814_/A _08891_/A _08878_/X _08879_/Y vssd1 vssd1 vccd1 vccd1 _08881_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_116_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07831_ _10871_/Q _07845_/B vssd1 vssd1 vccd1 vccd1 _07831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07941__A1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ _06871_/A _06871_/B _07761_/X vssd1 vssd1 vccd1 vccd1 _07763_/B sky130_fd_sc_hd__o21a_1
X_09501_ _09501_/A _09501_/B _09501_/C vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__nand3_1
X_06713_ _06719_/B _06635_/B _06634_/A vssd1 vssd1 vccd1 vccd1 _06714_/B sky130_fd_sc_hd__o21a_1
X_07693_ _07693_/A _07693_/B vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__xor2_1
XFILLER_65_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08939__D_N input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09432_ _09432_/A vssd1 vssd1 vccd1 vccd1 _10066_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06644_ _06841_/A _06408_/B _06408_/C vssd1 vssd1 vccd1 vccd1 _06645_/B sky130_fd_sc_hd__a21oi_1
XFILLER_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09363_ _09420_/A _10885_/Q vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__nor2_1
X_06575_ _10973_/Q _06575_/B vssd1 vssd1 vccd1 vccd1 _06951_/A sky130_fd_sc_hd__nand2_1
X_08314_ input34/X vssd1 vssd1 vccd1 vccd1 _08314_/Y sky130_fd_sc_hd__inv_2
X_05526_ _10711_/Q vssd1 vssd1 vccd1 vccd1 _06115_/A sky130_fd_sc_hd__clkbuf_4
X_09294_ _10343_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__and2_1
XFILLER_20_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08245_ _06105_/B _08058_/X _08243_/Y _08244_/Y _08062_/X vssd1 vssd1 vccd1 vccd1
+ _08245_/Y sky130_fd_sc_hd__a311oi_1
XFILLER_166_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05457_ _09020_/A _05283_/Y _05286_/B _08994_/A vssd1 vssd1 vccd1 vccd1 _05457_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_119_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07658__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08176_ _06187_/X _08164_/X _08165_/X _05692_/A _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08176_/X sky130_fd_sc_hd__o221a_1
X_05388_ _05388_/A _05392_/A vssd1 vssd1 vccd1 vccd1 _05389_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07127_ _07748_/B _07147_/A vssd1 vssd1 vccd1 vccd1 _07133_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07058_ _07197_/B vssd1 vssd1 vccd1 vccd1 _07076_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_161_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_30_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06009_ _10579_/Q vssd1 vssd1 vccd1 vccd1 _08236_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07393__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10971_ _10971_/CLK _10971_/D vssd1 vssd1 vccd1 vccd1 _10971_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08893__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10976_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07999__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06120__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07568__A _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10405_ _10940_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10405_/X sky130_fd_sc_hd__and2_1
XFILLER_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10336_ _10291_/S _10324_/A _10334_/Y _10335_/Y _10334_/A vssd1 vssd1 vccd1 vccd1
+ _10336_/X sky130_fd_sc_hd__o32a_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10266_/X _10259_/X _10257_/B vssd1 vssd1 vccd1 vccd1 _10268_/A sky130_fd_sc_hd__a21o_1
XFILLER_97_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08176__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08176__B2 _05692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10198_ _10198_/A _10198_/B vssd1 vssd1 vccd1 vccd1 _10198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06360_ _06360_/A _09302_/B _06736_/A vssd1 vssd1 vccd1 vccd1 _06360_/X sky130_fd_sc_hd__or3_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08100__A1 _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05311_ _10674_/Q _10673_/Q _05844_/B vssd1 vssd1 vccd1 vccd1 _05834_/A sky130_fd_sc_hd__or3_1
XANTENNA__08100__B2 _08098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06291_ _10910_/Q vssd1 vssd1 vccd1 vccd1 _06993_/A sky130_fd_sc_hd__buf_2
X_08030_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08030_/X sky130_fd_sc_hd__buf_4
Xinput30 io_wbs_m2s_data[22] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_4
XFILLER_163_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput41 io_wbs_m2s_data[3] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_8
XFILLER_155_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09981_ _09907_/A _09907_/B _09911_/A vssd1 vssd1 vccd1 vccd1 _09982_/B sky130_fd_sc_hd__o21a_1
XFILLER_103_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08932_ _08929_/Y _08930_/X _08931_/X vssd1 vssd1 vccd1 vccd1 _10830_/D sky130_fd_sc_hd__o21a_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08167__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08863_ _08658_/X _08860_/X _08866_/B _08862_/X vssd1 vssd1 vccd1 vccd1 _08864_/B
+ sky130_fd_sc_hd__a31oi_1
X_07814_ _10867_/Q _07824_/B vssd1 vssd1 vccd1 vccd1 _07814_/Y sky130_fd_sc_hd__nand2_1
XFILLER_84_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08794_ _06202_/X _08728_/X _08729_/X _10813_/Q vssd1 vssd1 vccd1 vccd1 _08794_/X
+ sky130_fd_sc_hd__a22o_1
X_07745_ _07745_/A _07745_/B vssd1 vssd1 vccd1 vccd1 _07746_/B sky130_fd_sc_hd__xnor2_1
XFILLER_72_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07677_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09415_ _09443_/B _09487_/A _09411_/A _09449_/A _10964_/Q vssd1 vssd1 vccd1 vccd1
+ _09454_/A sky130_fd_sc_hd__o2111a_1
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06627_ _06841_/A _06627_/B vssd1 vssd1 vccd1 vccd1 _06719_/B sky130_fd_sc_hd__nand2_2
XFILLER_25_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09346_ _09346_/A _09346_/B vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__nor2_2
X_06558_ _10972_/Q _06558_/B _06558_/C vssd1 vssd1 vccd1 vccd1 _06558_/X sky130_fd_sc_hd__and3_1
XFILLER_166_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05509_ _05350_/X _05503_/X _05506_/X _07885_/A vssd1 vssd1 vccd1 vccd1 _10560_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _08025_/A _09276_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09277_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06489_ _06600_/A _06489_/B vssd1 vssd1 vccd1 vccd1 _06541_/C sky130_fd_sc_hd__nand2_2
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08228_ _08228_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08228_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_154_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08159_ _08158_/X _08160_/B _08058_/A vssd1 vssd1 vccd1 vccd1 _08159_/X sky130_fd_sc_hd__a21bo_1
XFILLER_106_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10121_ _10120_/X _10101_/A _10121_/S vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10052_ _10052_/A _10051_/A vssd1 vssd1 vccd1 vccd1 _10053_/B sky130_fd_sc_hd__or2b_1
XFILLER_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07851__A _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input19_A io_wbs_m2s_data[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07570__B _09920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10954_ _10954_/CLK _10954_/D vssd1 vssd1 vccd1 vccd1 _10954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08330__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08330__B2 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10885_ _10984_/CLK _10885_/D vssd1 vssd1 vccd1 vccd1 _10885_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _10317_/X _10318_/Y _10329_/S vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__mux2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05860_ _08251_/A _05859_/Y _05857_/B _05858_/Y _10701_/Q vssd1 vssd1 vccd1 vccd1
+ _05860_/X sky130_fd_sc_hd__a32o_1
XFILLER_66_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05791_ _05791_/A _05791_/B vssd1 vssd1 vccd1 vccd1 _05791_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07530_ _07638_/B _07639_/A vssd1 vssd1 vccd1 vccd1 _07632_/B sky130_fd_sc_hd__or2b_1
XFILLER_35_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07461_ _07461_/A _07461_/B _07471_/A vssd1 vssd1 vccd1 vccd1 _07462_/B sky130_fd_sc_hd__nor3_1
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06412_ _06412_/A _06412_/B vssd1 vssd1 vccd1 vccd1 _06732_/A sky130_fd_sc_hd__nor2_1
X_09200_ _10814_/Q _09168_/X _09079_/X _10727_/Q _09199_/X vssd1 vssd1 vccd1 vccd1
+ _09200_/X sky130_fd_sc_hd__a221o_1
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07392_ _07391_/A _07163_/B _07588_/A vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__o21ai_1
XFILLER_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06343_ _06343_/A _06371_/C _06352_/C vssd1 vssd1 vccd1 vccd1 _06346_/A sky130_fd_sc_hd__or3_1
X_09131_ _09153_/A _09131_/B vssd1 vssd1 vccd1 vccd1 _10842_/D sky130_fd_sc_hd__nor2_4
XFILLER_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09821__A1 _09754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09062_ _09056_/X _09061_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10838_/D sky130_fd_sc_hd__o21a_4
X_06274_ _06305_/A _06274_/B vssd1 vssd1 vccd1 vccd1 _06371_/A sky130_fd_sc_hd__xor2_4
XFILLER_163_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08013_ _08013_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08013_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09964_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__or2_1
XFILLER_134_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08915_ _08921_/A _08915_/B vssd1 vssd1 vccd1 vccd1 _08915_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_131_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _09820_/B _09822_/B _09820_/A vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__o21bai_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08846_ _08844_/A _08844_/B _08845_/Y _08814_/A vssd1 vssd1 vccd1 vccd1 _08846_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08778_/C sky130_fd_sc_hd__nand2_1
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09101__A1_N _10938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05989_ input51/X vssd1 vssd1 vccd1 vccd1 _08462_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _07728_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07730_/A sky130_fd_sc_hd__nand2_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08312__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07659_ _07659_/A _07659_/B vssd1 vssd1 vccd1 vccd1 _07688_/B sky130_fd_sc_hd__xor2_1
XFILLER_14_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_83_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10926_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10670_ _10671_/CLK _10670_/D vssd1 vssd1 vccd1 vccd1 _10670_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _09329_/A _09329_/B vssd1 vssd1 vccd1 vccd1 _09400_/B sky130_fd_sc_hd__xnor2_4
XFILLER_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10537__A _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10256__B _10938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10186__A1 _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clock _10856_/CLK vssd1 vssd1 vccd1 vccd1 _10770_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10104_ _10104_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__05366__A _08198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10035_ _10035_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08551__A1 _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10937_ _10940_/CLK _10937_/D vssd1 vssd1 vccd1 vccd1 _10937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _10881_/CLK _10868_/D vssd1 vssd1 vccd1 vccd1 _10868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09301__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10799_ _10942_/CLK _10799_/D vssd1 vssd1 vccd1 vccd1 _10799_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10413__A2 _10722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07475__B _07475_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06250__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_77_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ _07625_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _06962_/B sky130_fd_sc_hd__and2_1
XFILLER_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08700_ _10803_/Q vssd1 vssd1 vccd1 vccd1 _08701_/A sky130_fd_sc_hd__clkbuf_2
X_05912_ _10648_/Q _05912_/B vssd1 vssd1 vccd1 vccd1 _05913_/B sky130_fd_sc_hd__xor2_1
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09680_ _09867_/B _09737_/A vssd1 vssd1 vccd1 vccd1 _09802_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06892_ _06902_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _06894_/A sky130_fd_sc_hd__xor2_4
XFILLER_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08631_ _10793_/Q _10792_/Q _08631_/C vssd1 vssd1 vccd1 vccd1 _08638_/C sky130_fd_sc_hd__and3_1
X_05843_ _05844_/B _05844_/C _05844_/A vssd1 vssd1 vccd1 vccd1 _05845_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__06553__B1 _10497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08562_ _08531_/X _08565_/C _10774_/Q _08531_/A vssd1 vssd1 vccd1 vccd1 _08562_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_05774_ _10710_/Q vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__inv_2
XFILLER_70_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07513_ _07513_/A _07516_/A vssd1 vssd1 vccd1 vccd1 _07514_/B sky130_fd_sc_hd__nand2_1
X_08493_ _08633_/A vssd1 vssd1 vccd1 vccd1 _10355_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07444_ _07717_/A _07444_/B vssd1 vssd1 vccd1 vccd1 _07445_/C sky130_fd_sc_hd__nor2_1
XFILLER_23_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07375_ _07375_/A vssd1 vssd1 vccd1 vccd1 _07391_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09114_ _09114_/A vssd1 vssd1 vccd1 vccd1 _09114_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06326_ _10928_/Q _10911_/Q _06805_/A _06805_/B _06293_/A vssd1 vssd1 vccd1 vccd1
+ _06851_/B sky130_fd_sc_hd__a221o_1
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09045_ _09599_/A vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__clkbuf_2
X_06257_ _08557_/A vssd1 vssd1 vccd1 vccd1 _06257_/X sky130_fd_sc_hd__buf_2
XFILLER_136_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10168__A1 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06188_ _10595_/Q vssd1 vssd1 vccd1 vccd1 _06189_/A sky130_fd_sc_hd__inv_2
XFILLER_116_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09947_ _10129_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _10023_/B sky130_fd_sc_hd__nand2_1
XFILLER_77_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _09953_/A _09878_/B vssd1 vssd1 vccd1 vccd1 _09882_/A sky130_fd_sc_hd__xor2_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08829_ _08841_/A _08841_/B _08827_/X _08828_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08829_/X sky130_fd_sc_hd__o311a_1
XFILLER_18_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09861__B_N _07008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _10784_/CLK _10722_/D vssd1 vssd1 vccd1 vccd1 _10722_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06745__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10653_ _10653_/CLK _10653_/D vssd1 vssd1 vccd1 vccd1 _10653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10584_ _10962_/CLK _10584_/D vssd1 vssd1 vccd1 vccd1 _10584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10018_ _10017_/A _10017_/B _10016_/Y vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__o21bai_1
XFILLER_110_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10331__A1 _09379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08288__B1 _08287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05490_ _05490_/A vssd1 vssd1 vccd1 vccd1 _05490_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10177__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07160_ _07280_/A _07159_/X vssd1 vssd1 vccd1 vccd1 _07200_/A sky130_fd_sc_hd__or2b_1
XFILLER_157_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06111_ _10707_/Q _08324_/B vssd1 vssd1 vccd1 vccd1 _08332_/B sky130_fd_sc_hd__or2_1
XFILLER_30_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07091_ _07402_/A _07091_/B _07091_/C vssd1 vssd1 vccd1 vccd1 _07363_/B sky130_fd_sc_hd__or3_1
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06042_ _10705_/Q _08021_/A _05475_/X _05736_/A vssd1 vssd1 vccd1 vccd1 _06045_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ _09801_/A vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__inv_2
XANTENNA__08763__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07993_ _08563_/A vssd1 vssd1 vccd1 vccd1 _07993_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09732_ _09432_/A _09679_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__o21a_1
X_06944_ _06944_/A _06944_/B vssd1 vssd1 vccd1 vccd1 _07645_/A sky130_fd_sc_hd__nand2_2
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09663_ _09661_/X _09663_/B vssd1 vssd1 vccd1 vccd1 _09779_/B sky130_fd_sc_hd__and2b_1
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06875_ _06875_/A _06875_/B vssd1 vssd1 vccd1 vccd1 _06878_/A sky130_fd_sc_hd__xnor2_2
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05453__B _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08614_ _10788_/Q vssd1 vssd1 vccd1 vccd1 _08614_/Y sky130_fd_sc_hd__inv_2
X_05826_ _05525_/B _08034_/A _05831_/C vssd1 vssd1 vccd1 vccd1 _05826_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09594_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09595_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08545_ _08545_/A vssd1 vssd1 vccd1 vccd1 _10769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05757_ _08242_/A _05752_/Y _10559_/Q _08232_/A vssd1 vssd1 vccd1 vccd1 _05765_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08476_ _10779_/Q _10742_/Q _08476_/S vssd1 vssd1 vccd1 vccd1 _08477_/B sky130_fd_sc_hd__mux2_1
X_05688_ _05570_/X _05571_/X _05686_/X _05687_/X vssd1 vssd1 vccd1 vccd1 _05688_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07427_ _07428_/A _07428_/B _07428_/C vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__a21o_1
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07358_ _07070_/A _07398_/B _07562_/A vssd1 vssd1 vccd1 vccd1 _07359_/B sky130_fd_sc_hd__and3b_1
XANTENNA__08780__A _08992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06309_ _06734_/A _06309_/B vssd1 vssd1 vccd1 vccd1 _06731_/B sky130_fd_sc_hd__nand2_2
XFILLER_164_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07289_ _07289_/A _07305_/B _07304_/B vssd1 vssd1 vccd1 vccd1 _07289_/X sky130_fd_sc_hd__or3b_1
X_09028_ _09805_/A vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08754__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08939__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10313__A1 _09920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _10860_/CLK _10705_/D vssd1 vssd1 vccd1 vccd1 _10705_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10636_ _10666_/CLK _10636_/D vssd1 vssd1 vccd1 vccd1 _10636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10567_ _10855_/CLK _10567_/D vssd1 vssd1 vccd1 vccd1 _10567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10498_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06205__C1 _06200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput6 io_wbs_m2s_addr[11] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_37_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09170__B2 _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06660_ _06660_/A _06660_/B vssd1 vssd1 vccd1 vccd1 _06661_/B sky130_fd_sc_hd__nor2_1
XFILLER_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05611_ _10555_/Q _05663_/A _05663_/B _10556_/Q vssd1 vssd1 vccd1 vccd1 _05612_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06591_ _06591_/A _06591_/B vssd1 vssd1 vccd1 vccd1 _06591_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__05731__A1 _05728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08330_ input35/X _08248_/X _08088_/X _08324_/A _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08330_/X sky130_fd_sc_hd__o221a_1
X_05542_ _05482_/X _05741_/B _05541_/X vssd1 vssd1 vccd1 vccd1 _05641_/A sky130_fd_sc_hd__o21ai_1
XFILLER_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08261_ _08259_/X _08261_/B vssd1 vssd1 vccd1 vccd1 _08262_/A sky130_fd_sc_hd__and2b_1
X_05473_ _05479_/A vssd1 vssd1 vccd1 vccd1 _05517_/A sky130_fd_sc_hd__clkbuf_4
X_07212_ _07415_/A _07244_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07214_/A sky130_fd_sc_hd__or3b_1
XFILLER_165_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08192_ _06117_/C _08074_/X _08191_/Y _08044_/A _07988_/A vssd1 vssd1 vccd1 vccd1
+ _08192_/X sky130_fd_sc_hd__a32o_1
XFILLER_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ _10985_/Q _07327_/A _07490_/A vssd1 vssd1 vccd1 vccd1 _07144_/B sky130_fd_sc_hd__a21bo_1
XFILLER_118_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07074_ _07186_/B vssd1 vssd1 vccd1 vccd1 _07390_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_173_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08105__A _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06025_ _08096_/A vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__buf_4
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07976_ _07976_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07976_/X sky130_fd_sc_hd__or2_1
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09715_ _09780_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__xnor2_1
XFILLER_101_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06927_ _06938_/A _06938_/B _06926_/X vssd1 vssd1 vccd1 vccd1 _06937_/B sky130_fd_sc_hd__a21o_1
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09646_ _09695_/B _09646_/B vssd1 vssd1 vccd1 vccd1 _09647_/B sky130_fd_sc_hd__xnor2_2
X_06858_ _07780_/C _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06859_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05809_ _05787_/B _05791_/Y _05792_/Y _05802_/Y _05808_/X vssd1 vssd1 vccd1 vccd1
+ _05809_/X sky130_fd_sc_hd__a311o_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09623_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06789_ _06741_/A _06834_/B _06788_/X vssd1 vssd1 vccd1 vccd1 _06832_/A sky130_fd_sc_hd__o21ai_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _10765_/Q _08419_/B _08527_/X vssd1 vssd1 vccd1 vccd1 _10765_/D sky130_fd_sc_hd__a21o_1
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08121__C1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08459_ _10774_/Q _10737_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__mux2_1
XFILLER_50_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10421_ _10944_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__and2_1
XFILLER_137_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10352_ _10351_/X _06387_/B _10346_/X _10920_/Q vssd1 vssd1 vccd1 vccd1 _10920_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08015__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10264__B _10939_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_140_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10283_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10283_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input49_A io_wbs_m2s_stb vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10534__A1 _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10619_ _10652_/CLK _10619_/D vssd1 vssd1 vccd1 vccd1 _10619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08966__A1 _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10525__A1 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07830_ _10577_/Q vssd1 vssd1 vccd1 vccd1 _07845_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07761_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _07761_/X sky130_fd_sc_hd__or2_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09500_ _09542_/B _09499_/B _09499_/C vssd1 vssd1 vccd1 vccd1 _09501_/C sky130_fd_sc_hd__a21o_1
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06712_ _06718_/B _06712_/B vssd1 vssd1 vccd1 vccd1 _06722_/A sky130_fd_sc_hd__and2_1
X_07692_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09575_/C sky130_fd_sc_hd__and2b_1
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09431_ _09431_/A _09431_/B vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__xor2_4
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06643_ _06643_/A _06643_/B vssd1 vssd1 vccd1 vccd1 _06702_/B sky130_fd_sc_hd__xor2_4
XFILLER_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09362_ _09420_/A _10885_/Q vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__nand2_1
X_06574_ _06585_/A _06585_/B _06573_/C vssd1 vssd1 vccd1 vccd1 _06578_/B sky130_fd_sc_hd__a21o_1
XFILLER_80_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08313_ _09154_/A vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__buf_4
X_05525_ _05525_/A _05525_/B vssd1 vssd1 vccd1 vccd1 _10572_/D sky130_fd_sc_hd__nor2_1
XANTENNA__07457__A1 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09293_ hold9/X _09274_/X _09275_/X _09292_/X _09270_/X vssd1 vssd1 vccd1 vccd1 _09294_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08244_ _08244_/A _08306_/B vssd1 vssd1 vccd1 vccd1 _08244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05456_ _10618_/Q vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06843__A _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08175_ _08175_/A vssd1 vssd1 vccd1 vccd1 _08175_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_146_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05387_ _10622_/Q vssd1 vssd1 vccd1 vccd1 _05462_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07126_ _10985_/Q _07474_/B vssd1 vssd1 vccd1 vccd1 _07147_/A sky130_fd_sc_hd__nand2_1
XFILLER_134_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ _07166_/B vssd1 vssd1 vccd1 vccd1 _07197_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_06008_ _06008_/A vssd1 vssd1 vccd1 vccd1 _06008_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10516__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07959_ _08443_/A _07959_/B vssd1 vssd1 vccd1 vccd1 _07960_/A sky130_fd_sc_hd__or2_1
XANTENNA__05943__A1 _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10970_ _10970_/CLK _10970_/D vssd1 vssd1 vccd1 vccd1 _10970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09629_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09630_/B sky130_fd_sc_hd__and2_1
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08645__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05459__B1 _09078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06120__A1 _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10275__A _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _10389_/X _10720_/Q _10402_/X _10403_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10939_/D sky130_fd_sc_hd__o221a_1
XFILLER_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10335_ _10324_/A _10327_/A _10279_/S vssd1 vssd1 vccd1 vccd1 _10335_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10266_ _10938_/Q _10954_/Q vssd1 vssd1 vccd1 vccd1 _10266_/X sky130_fd_sc_hd__or2b_1
XFILLER_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10507__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10197_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09125__B2 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05310_ _05336_/A vssd1 vssd1 vccd1 vccd1 _05844_/B sky130_fd_sc_hd__clkbuf_2
X_06290_ _10927_/Q _10910_/Q vssd1 vssd1 vccd1 vccd1 _06293_/A sky130_fd_sc_hd__and2_1
XFILLER_174_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput20 io_wbs_m2s_data[13] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_4
Xinput31 io_wbs_m2s_data[23] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_4
XFILLER_128_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput42 io_wbs_m2s_data[4] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_8
XFILLER_162_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05279__A _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09980_ _09980_/A _09980_/B vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__xnor2_1
XFILLER_104_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08931_ input40/X _08819_/X _08820_/X hold11/A _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08931_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ input30/X _08830_/A _08831_/A hold4/A vssd1 vssd1 vccd1 vccd1 _08862_/X sky130_fd_sc_hd__a22o_1
XFILLER_112_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07813_ _06255_/X hold10/A _06257_/X _07812_/Y vssd1 vssd1 vccd1 vccd1 _10616_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08793_ _08803_/C _08790_/X _08791_/X _08792_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08793_/X sky130_fd_sc_hd__o311a_1
XFILLER_84_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07744_ _07744_/A _07744_/B vssd1 vssd1 vccd1 vccd1 _07745_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07675_ _07675_/A _07675_/B vssd1 vssd1 vccd1 vccd1 _07677_/A sky130_fd_sc_hd__nor2_1
X_09414_ _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09487_/A sky130_fd_sc_hd__and2_1
X_06626_ _06626_/A vssd1 vssd1 vccd1 vccd1 _06841_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09345_ _09344_/B _10892_/Q vssd1 vssd1 vccd1 vccd1 _09346_/B sky130_fd_sc_hd__and2b_1
XFILLER_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06557_ _06561_/B _07675_/B vssd1 vssd1 vccd1 vccd1 _06587_/C sky130_fd_sc_hd__and2_1
XFILLER_166_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05508_ _05353_/X _05503_/X _05506_/X _07882_/A vssd1 vssd1 vccd1 vccd1 _10559_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09276_ _08324_/A _07914_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09276_/X sky130_fd_sc_hd__mux2_1
X_06488_ _06567_/A vssd1 vssd1 vccd1 vccd1 _06600_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08227_ _08092_/X _08232_/B _08226_/X _08096_/X vssd1 vssd1 vccd1 vccd1 _08227_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_166_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05439_ _10642_/Q vssd1 vssd1 vccd1 vccd1 _07911_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06292__B _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ _08160_/A vssd1 vssd1 vccd1 vccd1 _08158_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_107_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07109_ _07215_/B vssd1 vssd1 vccd1 vccd1 _07125_/A sky130_fd_sc_hd__buf_2
XFILLER_106_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08089_ _10528_/A _08086_/X _08088_/X _05733_/X _08166_/A vssd1 vssd1 vccd1 vccd1
+ _08090_/B sky130_fd_sc_hd__o221a_1
XFILLER_107_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10120_ _10102_/A _10102_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _10120_/X sky130_fd_sc_hd__a21bo_1
XFILLER_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10051_ _10051_/A _10052_/A vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__or2b_1
XFILLER_88_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _10954_/CLK _10953_/D vssd1 vssd1 vccd1 vccd1 _10953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10884_ _10984_/CLK _10884_/D vssd1 vssd1 vccd1 vccd1 _10884_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09291__A0 _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10318_ _10307_/A _10309_/Y _10307_/B vssd1 vssd1 vccd1 vccd1 _10318_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10249_ _10249_/A vssd1 vssd1 vccd1 vccd1 _10249_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05790_ _05765_/C _05789_/X _05765_/B vssd1 vssd1 vccd1 vccd1 _05791_/B sky130_fd_sc_hd__a21bo_1
XFILLER_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07460_ _07460_/A _07460_/B vssd1 vssd1 vccd1 vccd1 _07746_/A sky130_fd_sc_hd__xnor2_2
XFILLER_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06411_ _06717_/A _06411_/B vssd1 vssd1 vccd1 vccd1 _06431_/A sky130_fd_sc_hd__or2_1
XFILLER_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07391_ _07391_/A _07391_/B vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__nand2_1
X_09130_ _09112_/X _09122_/Y _09129_/X vssd1 vssd1 vccd1 vccd1 _09131_/B sky130_fd_sc_hd__a21oi_1
X_06342_ _06342_/A _06342_/B vssd1 vssd1 vccd1 vccd1 _06352_/C sky130_fd_sc_hd__xor2_2
XANTENNA__08085__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08085__B2 _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ _10487_/A _10474_/B _10495_/B _10508_/A _09060_/X vssd1 vssd1 vccd1 vccd1
+ _09061_/X sky130_fd_sc_hd__a221o_1
X_06273_ _06263_/Y _06270_/A _06276_/A _06272_/Y vssd1 vssd1 vccd1 vccd1 _06274_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ input29/X _08002_/X _08011_/X _08006_/X vssd1 vssd1 vccd1 vccd1 _10669_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09585__A1 _10968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__B2 _10967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_2_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10978_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08793__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__and2_1
XFILLER_103_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08914_ _08927_/A _08921_/B vssd1 vssd1 vccd1 vccd1 _08915_/B sky130_fd_sc_hd__or2_1
XFILLER_98_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _09894_/A _09893_/Y vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__or2b_1
XFILLER_85_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08845_ _08845_/A vssd1 vssd1 vccd1 vccd1 _08845_/Y sky130_fd_sc_hd__inv_2
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08778_/B sky130_fd_sc_hd__or2_1
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05988_ _09078_/A _05975_/X _05987_/Y _05977_/X vssd1 vssd1 vccd1 vccd1 _10575_/D
+ sky130_fd_sc_hd__a211oi_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05472__A _05490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07731_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07658_ _07670_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07659_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06609_ _06758_/A vssd1 vssd1 vccd1 vccd1 _06856_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07589_ _07589_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07593_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09328_ _09312_/X _09325_/Y _09402_/B _09327_/X vssd1 vssd1 vccd1 vccd1 _10867_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_167_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08076__B2 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06087__B1 _05813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ _09259_/A _09259_/B vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__and2_4
XFILLER_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08023__A _08023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09328__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _10029_/A _10029_/B _10022_/A vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__o21ai_2
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input31_A io_wbs_m2s_data[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10034_ _09955_/A _09955_/B _09960_/A vssd1 vssd1 vccd1 vccd1 _10035_/B sky130_fd_sc_hd__o21ai_2
XFILLER_75_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10936_ _10940_/CLK _10936_/D vssd1 vssd1 vccd1 vccd1 _10936_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _10967_/CLK _10867_/D vssd1 vssd1 vccd1 vccd1 _10867_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10798_/CLK _10798_/D vssd1 vssd1 vccd1 vccd1 _10798_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06960_ _07630_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__and2b_1
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05911_ _05911_/A _05911_/B vssd1 vssd1 vccd1 vccd1 _05911_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_67_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06891_ _06891_/A _06891_/B vssd1 vssd1 vccd1 vccd1 _06930_/A sky130_fd_sc_hd__xnor2_4
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08630_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _10792_/D sky130_fd_sc_hd__nor2_1
X_05842_ _10673_/Q vssd1 vssd1 vccd1 vccd1 _05844_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _10773_/Q _08559_/B _08560_/X _08030_/X vssd1 vssd1 vccd1 vccd1 _10773_/D
+ sky130_fd_sc_hd__o211a_1
X_05773_ _10709_/Q vssd1 vssd1 vccd1 vccd1 _06113_/A sky130_fd_sc_hd__inv_2
X_07512_ _07522_/B _07512_/B vssd1 vssd1 vccd1 vccd1 _07657_/A sky130_fd_sc_hd__nor2_1
XFILLER_35_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08492_ input51/X _09403_/B vssd1 vssd1 vccd1 vccd1 _08633_/A sky130_fd_sc_hd__nor2_1
XFILLER_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07443_ _07715_/C _07726_/B _07732_/B _07442_/X vssd1 vssd1 vccd1 vccd1 _07444_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_11_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07374_ _07374_/A _07374_/B vssd1 vssd1 vccd1 vccd1 _07456_/A sky130_fd_sc_hd__xor2_2
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09113_ _09113_/A vssd1 vssd1 vccd1 vccd1 _09113_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06325_ _06734_/B _06318_/X _06735_/A _06322_/X _06324_/X vssd1 vssd1 vccd1 vccd1
+ _06805_/B sky130_fd_sc_hd__o311ai_4
XFILLER_129_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09044_ _09489_/A vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06256_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08557_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10373__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06187_ input18/X vssd1 vssd1 vccd1 vccd1 _06187_/X sky130_fd_sc_hd__buf_4
XFILLER_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08230__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08230__B2 _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09946_ _10031_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__xnor2_1
XFILLER_132_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _09943_/B _09877_/B vssd1 vssd1 vccd1 vccd1 _09878_/B sky130_fd_sc_hd__or2_1
XFILLER_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _08841_/B _08827_/X _08841_/A vssd1 vssd1 vccd1 vccd1 _08828_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ _08759_/A _08759_/B vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__and2_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10940_/CLK _10721_/D vssd1 vssd1 vccd1 vccd1 _10721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09246__A0 _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10652_ _10652_/CLK _10652_/D vssd1 vssd1 vccd1 vccd1 _10652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _10657_/CLK _10583_/D vssd1 vssd1 vccd1 vccd1 _10583_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10283__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_21_clock_A _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08688__A _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07592__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10017_ _10017_/A _10017_/B _10016_/Y vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__or3b_1
XFILLER_76_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08288__A1 _08278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05840__A _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09312__A _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10919_ _10981_/CLK _10919_/D vssd1 vssd1 vccd1 vccd1 _10919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09237__A0 _08267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06110_ _10706_/Q _08317_/B vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__or2_1
XANTENNA__07767__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07090_ _07359_/A _07090_/B vssd1 vssd1 vccd1 vccd1 _07091_/C sky130_fd_sc_hd__or2_1
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06041_ _08105_/A _06038_/X _06040_/X vssd1 vssd1 vccd1 vccd1 _06071_/A sky130_fd_sc_hd__o21ai_1
XFILLER_161_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09800_ _09867_/B _09937_/A vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_82_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10909_/CLK sky130_fd_sc_hd__clkbuf_16
X_07992_ _10441_/A vssd1 vssd1 vccd1 vccd1 _08563_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__08598__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09731_ _09731_/A _09731_/B vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__xnor2_2
X_06943_ _06943_/A _06943_/B _06943_/C vssd1 vssd1 vccd1 vccd1 _06944_/B sky130_fd_sc_hd__nand3_1
XFILLER_101_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09662_ _09662_/A _09662_/B _09660_/Y vssd1 vssd1 vccd1 vccd1 _09663_/B sky130_fd_sc_hd__or3b_1
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06874_ _06874_/A _06874_/B vssd1 vssd1 vccd1 vccd1 _06881_/A sky130_fd_sc_hd__or2_2
XFILLER_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08613_ _08613_/A vssd1 vssd1 vccd1 vccd1 _10787_/D sky130_fd_sc_hd__clkbuf_1
X_05825_ _05844_/C vssd1 vssd1 vccd1 vccd1 _05831_/C sky130_fd_sc_hd__clkbuf_2
X_09593_ _09594_/A _09594_/B vssd1 vssd1 vccd1 vccd1 _09593_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08544_ _08580_/B _08544_/B _08544_/C vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__and3_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08279__A1 _08278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05756_ _05756_/A vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_70_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_clock _10856_/CLK vssd1 vssd1 vccd1 vccd1 _10833_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08475_ _08475_/A vssd1 vssd1 vccd1 vccd1 _10741_/D sky130_fd_sc_hd__clkbuf_1
X_05687_ _08350_/A _05687_/B vssd1 vssd1 vccd1 vccd1 _05687_/X sky130_fd_sc_hd__or2_1
XANTENNA__10368__A _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07426_ _07426_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07428_/C sky130_fd_sc_hd__xnor2_1
XFILLER_51_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07357_ _07377_/A _07390_/B _07357_/C vssd1 vssd1 vccd1 vccd1 _07360_/A sky130_fd_sc_hd__and3_1
XFILLER_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_clock _10856_/CLK vssd1 vssd1 vccd1 vccd1 _10830_/CLK sky130_fd_sc_hd__clkbuf_16
X_06308_ _10923_/Q _10906_/Q vssd1 vssd1 vccd1 vccd1 _06309_/B sky130_fd_sc_hd__or2_1
XFILLER_109_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07288_ _07302_/A _07344_/A _07279_/B vssd1 vssd1 vccd1 vccd1 _07304_/B sky130_fd_sc_hd__o21ai_1
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ _09555_/A vssd1 vssd1 vccd1 vccd1 _09805_/A sky130_fd_sc_hd__clkbuf_2
X_06239_ _06253_/B vssd1 vssd1 vccd1 vccd1 _06249_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_151_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09892__A _09893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09340__A_N _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09929_ _09929_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _10704_/CLK _10704_/D vssd1 vssd1 vccd1 vccd1 _10704_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10635_ _10666_/CLK _10635_/D vssd1 vssd1 vccd1 vccd1 _10635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07587__A _07592_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10566_ _10674_/CLK _10566_/D vssd1 vssd1 vccd1 vccd1 _10566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10497_/Y sky130_fd_sc_hd__nand2_1
XFILLER_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 io_wbs_m2s_addr[1] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XFILLER_65_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05610_ _05610_/A _05610_/B vssd1 vssd1 vccd1 vccd1 _05610_/X sky130_fd_sc_hd__and2_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06590_ _06951_/A _06951_/B vssd1 vssd1 vccd1 vccd1 _06952_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05570__A _08339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05541_ _05643_/A _05539_/Y _05540_/X vssd1 vssd1 vccd1 vccd1 _05541_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08260_ input28/X _08212_/X _08124_/X _05598_/X _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08261_/B sky130_fd_sc_hd__o221a_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05472_ _05490_/A _05472_/B vssd1 vssd1 vccd1 vccd1 _05479_/A sky130_fd_sc_hd__or2_1
XANTENNA__08881__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07211_ _07211_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07244_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08191_ _08191_/A _08191_/B vssd1 vssd1 vccd1 vccd1 _08191_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_119_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07142_ _10986_/Q _07142_/B vssd1 vssd1 vccd1 vccd1 _07490_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08433__A1 _10218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07073_ _07137_/A vssd1 vssd1 vccd1 vccd1 _07377_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06024_ _06024_/A vssd1 vssd1 vccd1 vccd1 _08096_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08197__B1 _05877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07944__A0 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07975_ _06172_/X _07965_/X _07974_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10656_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09714_ _09553_/A _09656_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09715_/B sky130_fd_sc_hd__a21oi_1
X_06926_ _06925_/B _06926_/B vssd1 vssd1 vccd1 vccd1 _06926_/X sky130_fd_sc_hd__and2b_1
XFILLER_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09645_ _09596_/A _09595_/B _09593_/Y vssd1 vssd1 vccd1 vccd1 _09646_/B sky130_fd_sc_hd__a21oi_2
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06857_ _07682_/A _06857_/B _06857_/C vssd1 vssd1 vccd1 vccd1 _06859_/A sky130_fd_sc_hd__and3_1
XFILLER_82_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05808_ _05785_/B _05807_/Y _05528_/A _05564_/A vssd1 vssd1 vccd1 vccd1 _05808_/X
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__nand2_4
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _10506_/A _07784_/B _07773_/B _06900_/A vssd1 vssd1 vccd1 vccd1 _06788_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08527_ _06124_/A _10394_/B _08418_/B _07899_/A vssd1 vssd1 vccd1 vccd1 _08527_/X
+ sky130_fd_sc_hd__a31o_1
X_05739_ _08132_/A _05739_/B vssd1 vssd1 vccd1 vccd1 _05742_/C sky130_fd_sc_hd__nor2_1
X_08458_ _08476_/S vssd1 vssd1 vccd1 vccd1 _08473_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07409_ _07540_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07410_/B sky130_fd_sc_hd__xor2_1
XFILLER_136_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08389_ _08383_/X _10736_/Q _08380_/X _08388_/X vssd1 vssd1 vccd1 vccd1 _10718_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10420_ _10408_/X _10724_/Q _10418_/X _10419_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10943_/D sky130_fd_sc_hd__o221a_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10351_ _10351_/A vssd1 vssd1 vccd1 vccd1 _10351_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_136_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10282_ _07013_/A _10253_/A _10281_/Y _08563_/X vssd1 vssd1 vccd1 vccd1 _10907_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09127__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05410__A1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09688__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07870__A _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08360__B1 _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06910__A1 _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06910__B2 _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08663__A1 _10799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10618_ _10652_/CLK _10618_/D vssd1 vssd1 vccd1 vccd1 _10618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10549_ _10554_/CLK _10549_/D vssd1 vssd1 vccd1 vccd1 _10549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09128__C1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ _06393_/A _06393_/B _07801_/A vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__a21o_1
XFILLER_38_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06711_ _06711_/A _06711_/B vssd1 vssd1 vccd1 vccd1 _06712_/B sky130_fd_sc_hd__or2_1
X_07691_ _09483_/A _09483_/B _07654_/A vssd1 vssd1 vccd1 vccd1 _09532_/B sky130_fd_sc_hd__o21ai_2
XFILLER_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09430_ _09430_/A _09430_/B vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06642_ _06642_/A _06642_/B vssd1 vssd1 vccd1 vccd1 _06885_/A sky130_fd_sc_hd__nor2_2
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06901__A1 _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ _09361_/A _09361_/B vssd1 vssd1 vccd1 vccd1 _09676_/B sky130_fd_sc_hd__nor2_4
XFILLER_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06573_ _06585_/A _06585_/B _06573_/C vssd1 vssd1 vccd1 vccd1 _06578_/A sky130_fd_sc_hd__nand3_1
X_08312_ _08157_/X _08307_/X _08309_/Y _08311_/X vssd1 vssd1 vccd1 vccd1 _10705_/D
+ sky130_fd_sc_hd__o31a_1
X_05524_ _10647_/Q vssd1 vssd1 vccd1 vccd1 _05525_/A sky130_fd_sc_hd__inv_2
X_09292_ _08352_/A _09291_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09292_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08243_ _08243_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _08243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05455_ _10619_/Q vssd1 vssd1 vccd1 vccd1 _05455_/X sky130_fd_sc_hd__buf_2
XFILLER_166_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08174_ _06117_/C _08074_/X _08173_/Y _08044_/X _07981_/A vssd1 vssd1 vccd1 vccd1
+ _08174_/X sky130_fd_sc_hd__a32o_1
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05386_ _10623_/Q vssd1 vssd1 vccd1 vccd1 _05462_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08116__A _08117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07125_ _07125_/A vssd1 vssd1 vccd1 vccd1 _07474_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07056_ _07056_/A _07056_/B vssd1 vssd1 vccd1 vccd1 _07166_/B sky130_fd_sc_hd__xor2_4
XFILLER_122_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06007_ input27/X vssd1 vssd1 vccd1 vccd1 _06008_/A sky130_fd_sc_hd__buf_6
XFILLER_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_68_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07958_ _10535_/A _08119_/A _07983_/A vssd1 vssd1 vccd1 vccd1 _07959_/B sky130_fd_sc_hd__mux2_1
XFILLER_29_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06909_ _09302_/B _06367_/A _06368_/B vssd1 vssd1 vccd1 vccd1 _06914_/A sky130_fd_sc_hd__o21a_2
X_07889_ _07889_/A vssd1 vssd1 vccd1 vccd1 _07889_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09628_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09559_ _09516_/A _09516_/C _09516_/B vssd1 vssd1 vccd1 vccd1 _09560_/B sky130_fd_sc_hd__a21boi_1
XFILLER_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09410__A _10966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10403_ _06172_/X _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__a21bo_1
XFILLER_152_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10334_ _10334_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10334_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07865__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10287_/A sky130_fd_sc_hd__nor2_2
XFILLER_127_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10196_ _10196_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _10197_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09291__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07105__A _10985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput10 io_wbs_m2s_addr[4] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_4
XFILLER_174_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput21 io_wbs_m2s_data[14] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_4
XFILLER_163_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput32 io_wbs_m2s_data[24] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_6
XFILLER_156_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput43 io_wbs_m2s_data[5] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_6
XFILLER_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09061__A1 _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09061__B2 _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08930_ _08920_/A _08927_/X _08928_/X _08814_/A vssd1 vssd1 vccd1 vccd1 _08930_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_115_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08861_ _08870_/C _08861_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07812_ _06134_/A _06258_/X _07807_/X _07809_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07812_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08792_ _08790_/X _08791_/X _08803_/C vssd1 vssd1 vccd1 vccd1 _08792_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07743_ _07743_/A _07743_/B _07743_/C vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__or3_1
XFILLER_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07674_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _09329_/A sky130_fd_sc_hd__nand2_2
XFILLER_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05689__A1 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07015__A _10982_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _09494_/B _09413_/B vssd1 vssd1 vccd1 vccd1 _09429_/A sky130_fd_sc_hd__or2_1
X_06625_ _06643_/A _06643_/B vssd1 vssd1 vccd1 vccd1 _06641_/B sky130_fd_sc_hd__nor2_1
XFILLER_13_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _10892_/Q _09344_/B vssd1 vssd1 vccd1 vccd1 _09346_/A sky130_fd_sc_hd__and2b_1
X_06556_ _10971_/Q _06575_/B vssd1 vssd1 vccd1 vccd1 _07675_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06854__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05507_ _05358_/X _05503_/X _05506_/X _07878_/A vssd1 vssd1 vccd1 vccd1 _10558_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09275_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09275_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06487_ _10973_/Q vssd1 vssd1 vccd1 vccd1 _06567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08226_ _08216_/X _08208_/A _08207_/B _06061_/A vssd1 vssd1 vccd1 vccd1 _08226_/X
+ sky130_fd_sc_hd__a31o_1
X_05438_ _07907_/A _05332_/Y _05437_/X vssd1 vssd1 vccd1 vccd1 _05438_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08157_/A vssd1 vssd1 vccd1 vccd1 _08157_/X sky130_fd_sc_hd__buf_2
X_05369_ _05369_/A _05369_/B vssd1 vssd1 vccd1 vccd1 _05369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07108_ _07747_/A _07108_/B vssd1 vssd1 vccd1 vccd1 _07215_/B sky130_fd_sc_hd__xnor2_4
X_08088_ _08355_/B vssd1 vssd1 vccd1 vccd1 _08088_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07039_ _07416_/A _07472_/A _07039_/C vssd1 vssd1 vccd1 vccd1 _07424_/A sky130_fd_sc_hd__and3_1
XFILLER_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10050_ _10050_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__xnor2_1
XFILLER_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09405__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _10954_/CLK _10952_/D vssd1 vssd1 vccd1 vccd1 _10952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10883_ _10986_/CLK _10883_/D vssd1 vssd1 vccd1 vccd1 _10883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10425__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09286__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10317_ _10307_/A _10310_/X _10307_/B vssd1 vssd1 vccd1 vccd1 _10317_/X sky130_fd_sc_hd__o21ba_1
XFILLER_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _10224_/A _10935_/Q _10233_/X _10235_/B _10247_/Y vssd1 vssd1 vccd1 vccd1
+ _10249_/A sky130_fd_sc_hd__o311a_1
XFILLER_140_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10179_ _06997_/B _10174_/X _10177_/X _10890_/Q vssd1 vssd1 vccd1 vccd1 _10890_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_94_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10113__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06410_ _06626_/A _06428_/B _06872_/A vssd1 vssd1 vccd1 vccd1 _06411_/B sky130_fd_sc_hd__a21oi_1
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07390_ _07592_/A _07390_/B vssd1 vssd1 vccd1 vccd1 _07391_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06341_ _06371_/B vssd1 vssd1 vccd1 vccd1 _06343_/A sky130_fd_sc_hd__inv_2
XANTENNA__10416__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09060_ _10935_/Q _10394_/C _10430_/B _10951_/Q vssd1 vssd1 vccd1 vccd1 _09060_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06272_ _10918_/Q _10901_/Q vssd1 vssd1 vccd1 vccd1 _06272_/Y sky130_fd_sc_hd__nor2_1
XFILLER_163_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08011_ _08268_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08011_/X sky130_fd_sc_hd__or2_1
XFILLER_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09962_ _09962_/A _09962_/B vssd1 vssd1 vccd1 vccd1 _09964_/B sky130_fd_sc_hd__xnor2_1
XFILLER_143_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08913_ _10828_/Q _08919_/B vssd1 vssd1 vccd1 vccd1 _08921_/B sky130_fd_sc_hd__and2_1
XFILLER_103_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09893_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _08844_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _08845_/A sky130_fd_sc_hd__or2_1
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05987_ _05992_/B _05986_/X _05993_/S vssd1 vssd1 vccd1 vccd1 _05987_/Y sky130_fd_sc_hd__a21oi_1
X_08775_ _08804_/A _08804_/B _08804_/C _08806_/A vssd1 vssd1 vccd1 vccd1 _08777_/B
+ sky130_fd_sc_hd__a31oi_1
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _07726_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07734_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08848__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07657_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09879__B _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06608_ _06607_/A _06607_/B _06607_/C vssd1 vssd1 vccd1 vccd1 _06614_/B sky130_fd_sc_hd__a21o_1
X_07588_ _07588_/A _07588_/B vssd1 vssd1 vccd1 vccd1 _07589_/B sky130_fd_sc_hd__xor2_1
XFILLER_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09327_ _10867_/Q _10283_/A vssd1 vssd1 vccd1 vccd1 _09327_/X sky130_fd_sc_hd__and2_1
X_06539_ _06532_/A _06532_/B _06538_/X vssd1 vssd1 vccd1 vccd1 _06542_/A sky130_fd_sc_hd__o21ba_1
XFILLER_22_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06087__A1 _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06087__B2 _05721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09258_ _08876_/A _09243_/X _09244_/X _09257_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09259_/B sky130_fd_sc_hd__a32o_1
XFILLER_139_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08209_ _08209_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08209_/Y sky130_fd_sc_hd__nor2_1
X_09189_ _05460_/B _09136_/A _09148_/X _05877_/X _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09189_/X sky130_fd_sc_hd__a221o_1
XFILLER_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08784__B1 _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08023__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10102_ _10102_/A _10102_/B vssd1 vssd1 vccd1 vccd1 _10104_/A sky130_fd_sc_hd__xnor2_4
XFILLER_161_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10033_ _10105_/B _10033_/B vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__xnor2_2
XFILLER_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input24_A io_wbs_m2s_data[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10935_ _10935_/CLK _10935_/D vssd1 vssd1 vccd1 vccd1 _10935_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05522__B1 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06494__A _10971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10866_ _10881_/CLK _10866_/D vssd1 vssd1 vccd1 vccd1 _10866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10797_ _10798_/CLK _10797_/D vssd1 vssd1 vccd1 vccd1 _10797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06250__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08527__B1 _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05910_ _06065_/A _05910_/B vssd1 vssd1 vccd1 vccd1 _05911_/B sky130_fd_sc_hd__xnor2_1
X_06890_ _06932_/B _06890_/B vssd1 vssd1 vccd1 vccd1 _06935_/A sky130_fd_sc_hd__xnor2_4
XFILLER_95_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05841_ _05337_/B _08018_/A _05844_/C vssd1 vssd1 vccd1 vccd1 _05841_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05772_ _10565_/Q vssd1 vssd1 vccd1 vccd1 _05772_/Y sky130_fd_sc_hd__inv_2
X_08560_ _08531_/X _08559_/X _10773_/Q _08531_/A vssd1 vssd1 vccd1 vccd1 _08560_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_07511_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07512_/B sky130_fd_sc_hd__nor2_1
X_08491_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08491_/X sky130_fd_sc_hd__buf_2
XFILLER_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07442_ _07573_/A vssd1 vssd1 vccd1 vccd1 _07442_/X sky130_fd_sc_hd__buf_2
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07373_ _07373_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07374_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06324_ _06323_/Y _06317_/A _06313_/A vssd1 vssd1 vccd1 vccd1 _06324_/X sky130_fd_sc_hd__o21a_1
X_09112_ _09112_/A vssd1 vssd1 vccd1 vccd1 _09112_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09043_ _10966_/Q vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06255_ _07848_/A vssd1 vssd1 vccd1 vccd1 _06255_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06186_ _06182_/X _06183_/X _06185_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10594_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08124__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06241__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09945_ _09945_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__xnor2_1
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08518__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07682__B _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09876_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09877_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _10816_/Q hold13/A _08928_/B vssd1 vssd1 vccd1 vccd1 _08827_/X sky130_fd_sc_hd__o21a_1
XFILLER_161_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _08758_/A _08758_/B vssd1 vssd1 vccd1 vccd1 _08804_/A sky130_fd_sc_hd__and2_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _10045_/A _10045_/B _07708_/X vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__o21ai_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _10802_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _10940_/CLK _10720_/D vssd1 vssd1 vccd1 vccd1 _10720_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10651_ _10651_/CLK _10651_/D vssd1 vssd1 vccd1 vccd1 _10651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10582_ _10814_/CLK _10582_/D vssd1 vssd1 vccd1 vccd1 _10582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08034__A _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06232__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07873__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07980__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10016_ _09945_/A _09945_/B _09929_/B vssd1 vssd1 vccd1 vccd1 _10016_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10918_ _10981_/CLK _10918_/D vssd1 vssd1 vccd1 vccd1 _10918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__A _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849_ _10850_/CLK _10849_/D vssd1 vssd1 vccd1 vccd1 _10849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10474__A _10495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05568__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06040_ _05749_/A _08289_/A _07976_/A _05711_/Y vssd1 vssd1 vccd1 vccd1 _06040_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07783__A _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07991_ _07991_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _07991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09730_ _09793_/B _09730_/B vssd1 vssd1 vccd1 vccd1 _09731_/B sky130_fd_sc_hd__xnor2_2
XFILLER_113_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06942_ _06942_/A _06942_/B vssd1 vssd1 vccd1 vccd1 _07641_/A sky130_fd_sc_hd__or2_1
XFILLER_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09661_ _09662_/A _09662_/B _09660_/Y vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__o21ba_1
X_06873_ _06383_/C _06873_/B vssd1 vssd1 vccd1 vccd1 _06874_/B sky130_fd_sc_hd__and2b_1
XFILLER_67_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08612_ _10355_/A _08612_/B _08612_/C vssd1 vssd1 vccd1 vccd1 _08613_/A sky130_fd_sc_hd__and3_1
X_05824_ _05854_/B vssd1 vssd1 vccd1 vccd1 _05844_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09592_ _09640_/A _09592_/B vssd1 vssd1 vccd1 vccd1 _09594_/B sky130_fd_sc_hd__or2_1
XFILLER_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08543_ _10769_/Q _08543_/B vssd1 vssd1 vccd1 vccd1 _08544_/C sky130_fd_sc_hd__nand2_1
XFILLER_39_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05755_ _10698_/Q vssd1 vssd1 vccd1 vccd1 _05756_/A sky130_fd_sc_hd__inv_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05686_ _05574_/X _05576_/X _05571_/X _05570_/X _05685_/X vssd1 vssd1 vccd1 vccd1
+ _05686_/X sky130_fd_sc_hd__a221o_1
X_08474_ _08477_/A _08474_/B vssd1 vssd1 vccd1 vccd1 _08475_/A sky130_fd_sc_hd__or2_1
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08119__A _08119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07425_ _07425_/A _07425_/B vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__or2_1
XFILLER_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07356_ _07560_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07406_/A sky130_fd_sc_hd__nand2_2
XFILLER_136_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06307_ _10923_/Q _10906_/Q vssd1 vssd1 vccd1 vccd1 _06734_/A sky130_fd_sc_hd__nand2_2
XFILLER_137_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07287_ _07287_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _07305_/B sky130_fd_sc_hd__xnor2_1
XFILLER_137_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06238_ _06238_/A vssd1 vssd1 vccd1 vccd1 _06238_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09026_ _10965_/Q vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__05478__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06169_ _10591_/Q vssd1 vssd1 vccd1 vccd1 _06170_/A sky130_fd_sc_hd__inv_2
XFILLER_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09928_ _10056_/C _10069_/B vssd1 vssd1 vccd1 vccd1 _09929_/B sky130_fd_sc_hd__or2_1
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09859_ _09859_/A vssd1 vssd1 vccd1 vccd1 _09859_/Y sky130_fd_sc_hd__inv_2
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05941__A _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _10703_/CLK _10703_/D vssd1 vssd1 vccd1 vccd1 _10703_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10634_ _10666_/CLK _10634_/D vssd1 vssd1 vccd1 vccd1 _10634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10565_ _10674_/CLK _10565_/D vssd1 vssd1 vccd1 vccd1 _10565_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05388__A _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07650__B1 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10496_ _10497_/B vssd1 vssd1 vccd1 vccd1 _10496_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06205__A1 _06202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output55_A _10987_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 io_wbs_m2s_addr[2] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_6
XFILLER_64_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05851__A _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09323__A _09323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05540_ _10574_/Q _10542_/Q vssd1 vssd1 vccd1 vccd1 _05540_/X sky130_fd_sc_hd__xor2_1
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05471_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05471_/X sky130_fd_sc_hd__clkbuf_4
X_07210_ _07210_/A _07260_/A vssd1 vssd1 vccd1 vccd1 _07275_/A sky130_fd_sc_hd__xnor2_1
X_08190_ _08092_/X _08196_/B _08189_/X _08096_/X vssd1 vssd1 vccd1 vccd1 _08190_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07141_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07296_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08433__A2 _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07072_ _10986_/Q vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06023_ _10583_/Q _06023_/B vssd1 vssd1 vccd1 vccd1 _06024_/A sky130_fd_sc_hd__nand2_2
XANTENNA__08197__A1 _08191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07944__A1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07974_ _07974_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07974_/X sky130_fd_sc_hd__or2_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09713_ _09713_/A _09713_/B vssd1 vssd1 vccd1 vccd1 _09723_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06925_ _06926_/B _06925_/B vssd1 vssd1 vccd1 vccd1 _06938_/B sky130_fd_sc_hd__xnor2_2
X_09644_ _09644_/A _09769_/C vssd1 vssd1 vccd1 vccd1 _09695_/B sky130_fd_sc_hd__xor2_2
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06856_ _06856_/A _07766_/B _06856_/C vssd1 vssd1 vccd1 vccd1 _06857_/C sky130_fd_sc_hd__and3_1
XFILLER_56_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05807_ _05807_/A _05807_/B vssd1 vssd1 vccd1 vccd1 _05807_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09575_ _09575_/A _09575_/B _09575_/C vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__or3_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06787_ _10506_/A _07773_/B vssd1 vssd1 vccd1 vccd1 _06834_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10379__A _10933_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _08526_/A vssd1 vssd1 vccd1 vccd1 _10764_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05738_ _08130_/A vssd1 vssd1 vccd1 vccd1 _08132_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08457_ _08457_/A vssd1 vssd1 vccd1 vccd1 _10736_/D sky130_fd_sc_hd__clkbuf_1
X_05669_ _10695_/Q _05612_/X _05610_/X _08224_/B _05668_/X vssd1 vssd1 vccd1 vccd1
+ _05669_/X sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_64_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07408_ _07543_/A _07361_/B _07407_/X vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__a21bo_1
X_08388_ _08395_/A _10752_/Q vssd1 vssd1 vccd1 vccd1 _08388_/X sky130_fd_sc_hd__or2_1
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07339_ _07528_/B _07339_/B vssd1 vssd1 vccd1 vccd1 _07526_/A sky130_fd_sc_hd__nand2_2
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10350_ _09312_/X _06371_/A _10346_/X _10919_/Q vssd1 vssd1 vccd1 vccd1 _10919_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09009_ _10948_/Q _10432_/C _09008_/X _10932_/Q vssd1 vssd1 vccd1 vccd1 _09009_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10281_ _10276_/Y _10279_/X _10280_/Y vssd1 vssd1 vccd1 vccd1 _10281_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09408__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09137__B1 _06212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09176__A1_N _10944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__A1 _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08360__A1 _05528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_81_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10925_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_70_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08663__A2 _08658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10617_ _10652_/CLK _10617_/D vssd1 vssd1 vccd1 vccd1 _10617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10548_ _10654_/CLK _10548_/D vssd1 vssd1 vccd1 vccd1 _10548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_170_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06007__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10479_ _06124_/X _10475_/X _10478_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10963_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06710_ _06711_/A _06711_/B vssd1 vssd1 vccd1 vccd1 _06718_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_34_clock _10856_/CLK vssd1 vssd1 vccd1 vccd1 _10821_/CLK sky130_fd_sc_hd__clkbuf_16
X_07690_ _07687_/A _07687_/B _07688_/B _09442_/A vssd1 vssd1 vccd1 vccd1 _09483_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_65_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06641_ _06641_/A _06641_/B _06641_/C vssd1 vssd1 vccd1 vccd1 _06642_/B sky130_fd_sc_hd__nor3_1
XFILLER_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09360_ _10902_/Q _10886_/Q vssd1 vssd1 vccd1 vccd1 _09361_/B sky130_fd_sc_hd__and2b_1
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06572_ _06571_/A _06571_/C _06571_/B vssd1 vssd1 vccd1 vccd1 _06594_/B sky130_fd_sc_hd__a21oi_1
X_08311_ input33/X _08248_/X _08088_/X _08305_/A _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08311_/X sky130_fd_sc_hd__o221a_1
XFILLER_21_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05523_ _05318_/X _05517_/X _05471_/X _07925_/A vssd1 vssd1 vccd1 vccd1 _10571_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09291_ _08351_/A _07925_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09291_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_49_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10860_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08242_ _08242_/A vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_05454_ _05454_/A vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__buf_2
XFILLER_166_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05385_ _10655_/Q _05389_/A vssd1 vssd1 vccd1 vccd1 _05385_/Y sky130_fd_sc_hd__xnor2_2
X_08173_ _08173_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08173_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_146_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08406__A2 _10743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07124_ _07137_/A _07229_/B vssd1 vssd1 vccd1 vccd1 _07748_/B sky130_fd_sc_hd__nand2_2
XFILLER_107_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07055_ _07113_/A _07475_/B _07112_/A vssd1 vssd1 vccd1 vccd1 _07056_/B sky130_fd_sc_hd__o21a_2
XFILLER_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06006_ _06006_/A vssd1 vssd1 vccd1 vccd1 _10578_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07971__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _08445_/A vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06908_ _06928_/A _06928_/B vssd1 vssd1 vccd1 vccd1 _06937_/A sky130_fd_sc_hd__xor2_4
XFILLER_56_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07888_ _07906_/A vssd1 vssd1 vccd1 vccd1 _07888_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_44_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09627_ _09682_/A _09627_/B vssd1 vssd1 vccd1 vccd1 _09629_/B sky130_fd_sc_hd__xor2_1
X_06839_ _06839_/A _06839_/B vssd1 vssd1 vccd1 vccd1 _06840_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09558_ _09597_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09560_/A sky130_fd_sc_hd__xnor2_1
XFILLER_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10437__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08509_ _10177_/A vssd1 vssd1 vccd1 vccd1 _08509_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09489_ _09489_/A _09555_/A _09642_/A _09492_/A vssd1 vssd1 vccd1 vccd1 _09618_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05459__A2 _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10402_ _10939_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10402_/X sky130_fd_sc_hd__and2_1
XFILLER_171_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ _10962_/Q _10946_/Q vssd1 vssd1 vccd1 vccd1 _10333_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10264_ _10955_/Q _10939_/Q vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08042__A _08062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _10932_/Q _10948_/Q vssd1 vssd1 vccd1 vccd1 _10196_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07881__A _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput11 io_wbs_m2s_addr[5] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput22 io_wbs_m2s_data[15] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput33 io_wbs_m2s_data[25] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput44 io_wbs_m2s_data[6] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_4
XFILLER_156_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10482__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_12_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08860_ _08870_/C _08861_/B vssd1 vssd1 vccd1 vccd1 _08860_/X sky130_fd_sc_hd__or2_1
XFILLER_112_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07811_ _07874_/A vssd1 vssd1 vccd1 vccd1 _07811_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08791_ _08778_/B _08803_/B vssd1 vssd1 vccd1 vccd1 _08791_/X sky130_fd_sc_hd__and2b_1
X_07742_ _07406_/A _07544_/A _07753_/A vssd1 vssd1 vccd1 vccd1 _07743_/C sky130_fd_sc_hd__a21oi_1
XFILLER_65_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07673_ _07673_/A _07673_/B vssd1 vssd1 vccd1 vccd1 _07674_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09412_ _09489_/A _09536_/B _09579_/A _10965_/Q vssd1 vssd1 vccd1 vccd1 _09413_/B
+ sky130_fd_sc_hd__a22oi_1
X_06624_ _06624_/A _06650_/A _06624_/C vssd1 vssd1 vccd1 vccd1 _06643_/B sky130_fd_sc_hd__and3_2
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09511__A _09599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09343_ _09343_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__nor2_1
X_06555_ _06555_/A _06555_/B vssd1 vssd1 vccd1 vccd1 _06585_/A sky130_fd_sc_hd__xnor2_2
XFILLER_34_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05506_ _05513_/A vssd1 vssd1 vccd1 vccd1 _05506_/X sky130_fd_sc_hd__clkbuf_1
X_09274_ _09274_/A vssd1 vssd1 vccd1 vccd1 _09274_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06486_ _06486_/A _06486_/B vssd1 vssd1 vccd1 vccd1 _06643_/A sky130_fd_sc_hd__xnor2_4
XFILLER_166_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08225_ _08233_/B vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__inv_2
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05437_ _10641_/Q _05332_/Y _05337_/X _05436_/X vssd1 vssd1 vccd1 vccd1 _05437_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08156_ _08156_/A vssd1 vssd1 vccd1 vccd1 _10689_/D sky130_fd_sc_hd__clkbuf_1
X_05368_ _10660_/Q _05886_/A _10661_/Q vssd1 vssd1 vccd1 vccd1 _05369_/B sky130_fd_sc_hd__o21a_1
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07107_ _10913_/Q _07747_/B vssd1 vssd1 vccd1 vccd1 _07108_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08260__B1 _08124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10392__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05299_ _05374_/A vssd1 vssd1 vccd1 vccd1 _05886_/A sky130_fd_sc_hd__clkbuf_2
X_08087_ _08124_/A vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07038_ _07428_/B _07038_/B vssd1 vssd1 vccd1 vccd1 _07051_/A sky130_fd_sc_hd__and2_1
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08990_/C sky130_fd_sc_hd__nand2_1
XFILLER_29_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ _10971_/CLK _10951_/D vssd1 vssd1 vccd1 vccd1 _10951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10882_ _10986_/CLK _10882_/D vssd1 vssd1 vccd1 vccd1 _10882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08079__B1 _05733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10316_ _10316_/A _10316_/B vssd1 vssd1 vccd1 vccd1 _10320_/A sky130_fd_sc_hd__nor2_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10247_ _10247_/A vssd1 vssd1 vccd1 vccd1 _10247_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10178_ _07083_/A _10174_/X _10177_/X _10889_/Q vssd1 vssd1 vccd1 vccd1 _10889_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10361__A1 _08491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06340_ _06459_/B vssd1 vssd1 vccd1 vccd1 _07682_/B sky130_fd_sc_hd__buf_2
XFILLER_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06271_ _06275_/A _06275_/B vssd1 vssd1 vccd1 vccd1 _06276_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08010_ input28/X _08002_/X _08009_/Y _08006_/X vssd1 vssd1 vccd1 vccd1 _10668_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09399__A_N _09400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09961_ _09961_/A _09961_/B vssd1 vssd1 vccd1 vccd1 _09962_/B sky130_fd_sc_hd__nor2_1
XFILLER_104_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08912_ _10828_/Q _08918_/B vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09894_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08843_ _08871_/A _08873_/A vssd1 vssd1 vccd1 vccd1 _08844_/B sky130_fd_sc_hd__nor2_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08774_ _10810_/Q _10809_/Q _10808_/Q _08748_/X _08801_/B vssd1 vssd1 vccd1 vccd1
+ _08806_/A sky130_fd_sc_hd__o41a_1
X_05986_ input44/X input43/X vssd1 vssd1 vccd1 vccd1 _05986_/X sky130_fd_sc_hd__or2_1
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ _07726_/A _07732_/B _07577_/B _07576_/A vssd1 vssd1 vccd1 vccd1 _07735_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07656_ _07657_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__and2_1
XFILLER_25_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06607_ _06607_/A _06607_/B _06607_/C vssd1 vssd1 vccd1 vccd1 _06614_/A sky130_fd_sc_hd__nand3_1
X_07587_ _07592_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07588_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09326_ _09326_/A _09326_/B vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__or2_1
X_06538_ _06533_/A _06538_/B vssd1 vssd1 vccd1 vccd1 _06538_/X sky130_fd_sc_hd__and2b_1
XFILLER_166_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06087__A2 _08023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ _08298_/A _09256_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09257_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06469_ _06448_/B _06469_/B vssd1 vssd1 vccd1 vccd1 _06470_/B sky130_fd_sc_hd__and2b_1
XFILLER_154_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08208_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08208_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09188_ _09113_/A _09187_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09188_/Y sky130_fd_sc_hd__o21ai_1
X_08139_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08140_/B sky130_fd_sc_hd__and2_1
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10101_ _10101_/A _10101_/B vssd1 vssd1 vccd1 vccd1 _10102_/B sky130_fd_sc_hd__and2_1
XFILLER_108_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10032_ _10030_/X _09952_/B _10031_/X vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__o21a_1
XFILLER_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input17_A io_wbs_m2s_data[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05770__B2 _08317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10934_ _10940_/CLK _10934_/D vssd1 vssd1 vccd1 vccd1 _10934_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _10865_/CLK _10865_/D vssd1 vssd1 vccd1 vccd1 _10865_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _10935_/CLK _10796_/D vssd1 vssd1 vccd1 vccd1 _10796_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09297__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07027__A1 _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06015__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08527__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05840_ _08298_/A vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__inv_2
XFILLER_95_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05771_ _05771_/A vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__buf_2
XFILLER_48_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07510_ _07510_/A _07510_/B vssd1 vssd1 vccd1 vccd1 _07633_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08490_ _10181_/A vssd1 vssd1 vccd1 vccd1 _08514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07441_ _07574_/A vssd1 vssd1 vccd1 vccd1 _07715_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07372_ _07373_/A _07374_/A _07373_/B vssd1 vssd1 vccd1 vccd1 _07454_/B sky130_fd_sc_hd__and3_1
XFILLER_148_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09111_ _09111_/A vssd1 vssd1 vccd1 vccd1 _10841_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06323_ _10926_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _06323_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09042_ _07732_/A _08965_/Y _09036_/X _09038_/X _09041_/X vssd1 vssd1 vccd1 vccd1
+ _09042_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06254_ input40/X _06145_/B _06253_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10615_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06185_ _06185_/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_116_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _10012_/A _09944_/B vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__or2_1
XFILLER_86_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09236__A _09236_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input9_A io_wbs_m2s_addr[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _09876_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09943_/B sky130_fd_sc_hd__and2_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08817_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08841_/B sky130_fd_sc_hd__and2b_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09191__B2 _10726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _10809_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08758_/B sky130_fd_sc_hd__or2_1
XFILLER_173_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05969_ _08414_/A _08939_/C vssd1 vssd1 vccd1 vccd1 _06126_/D sky130_fd_sc_hd__or2_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _07708_/A _07605_/B vssd1 vssd1 vccd1 vccd1 _07708_/X sky130_fd_sc_hd__or2b_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08688_ _08688_/A vssd1 vssd1 vccd1 vccd1 _08688_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _07639_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _07693_/A sky130_fd_sc_hd__xor2_2
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10650_ _10651_/CLK _10650_/D vssd1 vssd1 vccd1 vccd1 _10650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ _09313_/B _09310_/C _09396_/A vssd1 vssd1 vccd1 vccd1 _09309_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10581_ _10914_/CLK _10581_/D vssd1 vssd1 vccd1 vccd1 _10581_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_167_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08315__A _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08034__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06217__C1 _06200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_59_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10017_/B sky130_fd_sc_hd__and2_1
XFILLER_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10917_ _10980_/CLK _10917_/D vssd1 vssd1 vccd1 vccd1 _10917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08209__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10848_ _10848_/CLK _10848_/D vssd1 vssd1 vccd1 vccd1 _10848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10779_ _10782_/CLK _10779_/D vssd1 vssd1 vccd1 vccd1 _10779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08996__A1 _05721_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07990_ _08015_/A vssd1 vssd1 vccd1 vccd1 _08021_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_99_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06941_ _06941_/A _06941_/B _06944_/A vssd1 vssd1 vccd1 vccd1 _06942_/B sky130_fd_sc_hd__and3_1
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09660_ _09713_/A _09713_/B vssd1 vssd1 vccd1 vccd1 _09660_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06872_ _06872_/A _06872_/B vssd1 vssd1 vccd1 vccd1 _06873_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08611_ _10787_/Q _08611_/B vssd1 vssd1 vccd1 vccd1 _08612_/C sky130_fd_sc_hd__nand2_1
X_05823_ _05823_/A vssd1 vssd1 vccd1 vccd1 _05854_/B sky130_fd_sc_hd__clkbuf_2
X_09591_ _09590_/B _09591_/B vssd1 vssd1 vccd1 vccd1 _09592_/B sky130_fd_sc_hd__and2b_1
XFILLER_94_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05734__B2 _05728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08542_ _10769_/Q _08543_/B vssd1 vssd1 vccd1 vccd1 _08544_/B sky130_fd_sc_hd__or2_1
X_05754_ _05751_/Y _10561_/Q _05752_/Y _08242_/A vssd1 vssd1 vccd1 vccd1 _05765_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08473_ _10778_/Q _10741_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08474_/B sky130_fd_sc_hd__mux2_1
X_05685_ _05679_/X _05683_/X _05576_/X _08339_/B _05684_/X vssd1 vssd1 vccd1 vccd1
+ _05685_/X sky130_fd_sc_hd__o221a_1
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08119__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _07424_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _07425_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07355_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07366_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06306_ _06263_/Y _06270_/A _06276_/A _06305_/X _06272_/Y vssd1 vssd1 vccd1 vccd1
+ _06730_/C sky130_fd_sc_hd__a311o_1
XANTENNA__05759__A _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07286_ _07286_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _07287_/B sky130_fd_sc_hd__nor2_1
XFILLER_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09025_ _10714_/Q _08990_/C _09024_/X vssd1 vssd1 vccd1 vccd1 _09025_/X sky130_fd_sc_hd__o21a_1
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06237_ input32/X _06225_/X _06236_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10608_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07974__A _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06168_ _10537_/A vssd1 vssd1 vccd1 vccd1 _06168_/X sky130_fd_sc_hd__buf_4
XFILLER_85_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06099_ _10689_/Q _08150_/B vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__or2_2
XFILLER_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09927_ _10056_/C _10069_/B vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_60_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09858_ _10076_/A _09858_/B vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _08804_/Y _08806_/Y _08801_/X _08802_/Y vssd1 vssd1 vccd1 vccd1 _08817_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09848_/B _09789_/B vssd1 vssd1 vccd1 vccd1 _09827_/B sky130_fd_sc_hd__and2_2
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08029__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ _10704_/CLK _10702_/D vssd1 vssd1 vccd1 vccd1 _10702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ _10666_/CLK _10633_/D vssd1 vssd1 vccd1 vccd1 _10633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10564_ _10640_/CLK _10564_/D vssd1 vssd1 vccd1 vccd1 _10564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10495_ _10495_/A _10495_/B vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__nand2_2
XFILLER_114_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 io_wbs_m2s_addr[3] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_8
XFILLER_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05470_ _05470_/A _05470_/B vssd1 vssd1 vccd1 vccd1 _05513_/A sky130_fd_sc_hd__nor2_2
XANTENNA__06963__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06141__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10485__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08969__A1 _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07140_ _07151_/A _07474_/B _07147_/B _07139_/X vssd1 vssd1 vccd1 vccd1 _07295_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07071_ _07357_/C _07283_/B vssd1 vssd1 vccd1 vccd1 _07284_/A sky130_fd_sc_hd__or2_1
XFILLER_118_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06022_ _08837_/A vssd1 vssd1 vccd1 vccd1 _10412_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_141_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07973_ _08027_/B vssd1 vssd1 vccd1 vccd1 _07988_/B sky130_fd_sc_hd__clkbuf_1
X_09712_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09723_/A sky130_fd_sc_hd__or2_1
XFILLER_68_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06924_ _06914_/A _06914_/B _06923_/X vssd1 vssd1 vccd1 vccd1 _06925_/B sky130_fd_sc_hd__a21oi_1
XFILLER_142_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09643_ _09764_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09769_/C sky130_fd_sc_hd__nand2_1
X_06855_ _06855_/A _06855_/B vssd1 vssd1 vccd1 vccd1 _06857_/B sky130_fd_sc_hd__xnor2_1
XFILLER_95_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05806_ _05768_/X _05805_/X _05785_/A vssd1 vssd1 vccd1 vccd1 _05807_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09574_ _09570_/A _09574_/B vssd1 vssd1 vccd1 vccd1 _09631_/B sky130_fd_sc_hd__and2b_1
X_06786_ _06786_/A vssd1 vssd1 vccd1 vccd1 _07773_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_83_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08525_ _10763_/Q _10529_/A vssd1 vssd1 vccd1 vccd1 _08526_/A sky130_fd_sc_hd__and2_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05737_ _08082_/B _05737_/B vssd1 vssd1 vccd1 vccd1 _05742_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08456_ _08460_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__or2_1
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05668_ _05877_/A _05615_/Y _05612_/X _10695_/Q _05667_/X vssd1 vssd1 vccd1 vccd1
+ _05668_/X sky130_fd_sc_hd__o221a_1
X_07407_ _07407_/A _07360_/A vssd1 vssd1 vccd1 vccd1 _07407_/X sky130_fd_sc_hd__or2b_1
XFILLER_23_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08409__B1 _08992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08387_ _08383_/X _10735_/Q _08380_/X _08386_/X vssd1 vssd1 vccd1 vccd1 _10717_/D
+ sky130_fd_sc_hd__o211a_1
X_05599_ _10561_/Q _05602_/A vssd1 vssd1 vccd1 vccd1 _05599_/X sky130_fd_sc_hd__xor2_1
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07338_ _07338_/A _07338_/B vssd1 vssd1 vccd1 vccd1 _07339_/B sky130_fd_sc_hd__or2_1
XFILLER_136_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07269_ _07269_/A _07269_/B _07514_/A vssd1 vssd1 vccd1 vccd1 _07270_/B sky130_fd_sc_hd__and3_1
XFILLER_137_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09008_ _09008_/A vssd1 vssd1 vccd1 vccd1 _09008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10280_ _10276_/Y _10279_/X _10253_/A vssd1 vssd1 vccd1 vccd1 _10280_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_133_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05946__A1 _08339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06113__A _06113_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05946__B2 _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09137__B2 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08345__C1 _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05952__A _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10616_ _10652_/CLK _10616_/D vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_2
XFILLER_174_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10547_ _10654_/CLK _10547_/D vssd1 vssd1 vccd1 vccd1 _10547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10478_ _10478_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10478_/X sky130_fd_sc_hd__or2_1
XFILLER_136_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06023__A _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09128__A1 _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07780__C _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06640_ _06641_/A _06641_/B _06641_/C vssd1 vssd1 vccd1 vccd1 _06642_/A sky130_fd_sc_hd__o21a_1
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06571_ _06571_/A _06571_/B _06571_/C vssd1 vssd1 vccd1 vccd1 _06594_/A sky130_fd_sc_hd__and3_1
XFILLER_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08310_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08310_/X sky130_fd_sc_hd__clkbuf_4
X_05522_ _05324_/X _05517_/X _05471_/X _07922_/A vssd1 vssd1 vccd1 vccd1 _10570_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_33_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09290_ _09290_/A vssd1 vssd1 vccd1 vccd1 _10863_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08241_ _08241_/A vssd1 vssd1 vccd1 vccd1 _10698_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_162_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05453_ _05453_/A _09107_/A vssd1 vssd1 vccd1 vccd1 _05453_/X sky130_fd_sc_hd__or2_1
XFILLER_159_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08172_ _08092_/X _08181_/B _08171_/X _08096_/X vssd1 vssd1 vccd1 vccd1 _08172_/X
+ sky130_fd_sc_hd__a31o_1
X_05384_ _10624_/Q vssd1 vssd1 vccd1 vccd1 _05461_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_119_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07123_ _07144_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07134_/A sky130_fd_sc_hd__xnor2_2
XFILLER_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_opt_2_0_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07054_ _07151_/A vssd1 vssd1 vccd1 vccd1 _07560_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08413__A _10495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06005_ _08483_/A _06005_/B vssd1 vssd1 vccd1 vccd1 _06006_/A sky130_fd_sc_hd__and2_1
XFILLER_130_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07956_ _07956_/A vssd1 vssd1 vccd1 vccd1 _10653_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__07971__B _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09244__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06907_ _06904_/X _06922_/B _06906_/X vssd1 vssd1 vccd1 vccd1 _06928_/B sky130_fd_sc_hd__a21oi_2
X_07887_ _07898_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _10635_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09626_ _09626_/A _09682_/B vssd1 vssd1 vccd1 vccd1 _09627_/B sky130_fd_sc_hd__nand2_1
XFILLER_44_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06838_ _06839_/A _06839_/B vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__or2_1
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ _09652_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__or2_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06769_ _06769_/A vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09898__B _09898_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08508_ _10790_/Q _08506_/X _08502_/X _10753_/Q vssd1 vssd1 vccd1 vccd1 _10753_/D
+ sky130_fd_sc_hd__a22o_1
X_09488_ _09488_/A vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08439_ _08443_/A _08439_/B vssd1 vssd1 vccd1 vccd1 _08440_/A sky130_fd_sc_hd__or2_1
XFILLER_157_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10401_ _10389_/X _10719_/Q _10398_/X _10400_/X _10392_/X vssd1 vssd1 vccd1 vccd1
+ _10938_/D sky130_fd_sc_hd__o221a_1
XFILLER_165_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05947__A _08339_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10332_ _10962_/Q _10946_/Q vssd1 vssd1 vccd1 vccd1 _10332_/X sky130_fd_sc_hd__or2_1
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08323__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10263_ _10939_/Q _10955_/Q vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__and2b_1
XFILLER_79_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08042__B _08352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input47_A io_wbs_m2s_data[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _10948_/Q _10932_/Q vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__and2b_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09154__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06018__A _06023_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 io_wbs_m2s_addr[6] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 io_wbs_m2s_data[16] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_4
Xinput34 io_wbs_m2s_data[26] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_8
Xinput45 io_wbs_m2s_data[7] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_2
XFILLER_155_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05857__A _08268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08233__A _08233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07810_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07874_/A sky130_fd_sc_hd__buf_4
X_08790_ _10812_/Q _08771_/A _08918_/B vssd1 vssd1 vccd1 vccd1 _08790_/X sky130_fd_sc_hd__o21a_1
XFILLER_112_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07741_ _07741_/A _07741_/B vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__xnor2_2
XFILLER_38_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07672_ _07673_/A _07673_/B vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__or2_1
XFILLER_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09411_ _09411_/A vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06623_ _06541_/C _06542_/A _06528_/Y vssd1 vssd1 vccd1 vccd1 _06624_/C sky130_fd_sc_hd__a21o_1
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09342_ _07028_/A _10893_/Q vssd1 vssd1 vccd1 vccd1 _09343_/B sky130_fd_sc_hd__and2b_1
X_06554_ _10972_/Q _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06555_/B sky130_fd_sc_hd__and3_1
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05505_ _05360_/X _05503_/X _05495_/X _07875_/A vssd1 vssd1 vccd1 vccd1 _10557_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09273_ _09273_/A vssd1 vssd1 vccd1 vccd1 _10860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06485_ _06486_/A _06486_/B vssd1 vssd1 vccd1 vccd1 _06641_/A sky130_fd_sc_hd__and2_1
XFILLER_138_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08224_ _08224_/A _08224_/B _08224_/C vssd1 vssd1 vccd1 vccd1 _08233_/B sky130_fd_sc_hd__and3_1
X_05436_ _07900_/A _05340_/X _05337_/B _10640_/Q _05435_/X vssd1 vssd1 vccd1 vccd1
+ _05436_/X sky130_fd_sc_hd__a221o_1
XFILLER_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08156_/A sky130_fd_sc_hd__and2_1
XFILLER_119_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05367_ _10629_/Q vssd1 vssd1 vccd1 vccd1 _05460_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07106_ _07384_/A _07137_/C vssd1 vssd1 vccd1 vccd1 _07144_/A sky130_fd_sc_hd__or2_2
XFILLER_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09239__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08260__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08086_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08086_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08260__B2 _05598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05298_ _10659_/Q _05373_/B vssd1 vssd1 vccd1 vccd1 _05374_/A sky130_fd_sc_hd__or2_1
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07037_ _07555_/B _07037_/B vssd1 vssd1 vccd1 vccd1 _07038_/B sky130_fd_sc_hd__nand2_1
XFILLER_122_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08012__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_80_clock _10977_/CLK vssd1 vssd1 vccd1 vccd1 _10971_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08988_ _09079_/A vssd1 vssd1 vccd1 vccd1 _08988_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07939_ _07939_/A vssd1 vssd1 vccd1 vccd1 _10648_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09512__B2 _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _10954_/CLK _10950_/D vssd1 vssd1 vccd1 vccd1 _10950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09609_ _09867_/A _09610_/C _09717_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09611_/A
+ sky130_fd_sc_hd__a22oi_1
X_10881_ _10881_/CLK _10881_/D vssd1 vssd1 vccd1 vccd1 _10881_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09276__A0 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__A _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10822_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ _10960_/Q _10944_/Q vssd1 vssd1 vccd1 vccd1 _10316_/B sky130_fd_sc_hd__and2b_1
XFILLER_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07892__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ _10246_/A _10246_/B _10246_/C vssd1 vssd1 vccd1 vccd1 _10247_/A sky130_fd_sc_hd__and3_1
XFILLER_140_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10177_ _10177_/A vssd1 vssd1 vccd1 vccd1 _10177_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08711__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06270_ _06270_/A _06270_/B vssd1 vssd1 vccd1 vccd1 _06275_/B sky130_fd_sc_hd__and2_1
XANTENNA__09019__B1 _08992_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10493__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09960_ _09960_/A _09960_/B vssd1 vssd1 vccd1 vccd1 _09962_/A sky130_fd_sc_hd__nand2_1
XFILLER_171_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08911_ _08904_/B _08907_/B _08904_/A vssd1 vssd1 vccd1 vccd1 _08921_/A sky130_fd_sc_hd__o21bai_1
XFILLER_131_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09961_/B _09891_/B vssd1 vssd1 vccd1 vccd1 _09893_/B sky130_fd_sc_hd__or2_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08842_ _10818_/Q hold3/A _10816_/Q hold13/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08873_/A
+ sky130_fd_sc_hd__o41a_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08773_ _08773_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05985_ input44/X input43/X vssd1 vssd1 vccd1 vccd1 _05992_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07724_ _07724_/A _07724_/B vssd1 vssd1 vccd1 vccd1 _07740_/A sky130_fd_sc_hd__or2_1
XFILLER_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07655_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07657_/B sky130_fd_sc_hd__and2_1
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06606_ _06680_/A _06680_/B vssd1 vssd1 vccd1 vccd1 _06681_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _07586_/A _07586_/B vssd1 vssd1 vccd1 vccd1 _07751_/A sky130_fd_sc_hd__xnor2_1
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09325_ _09326_/A _09326_/B vssd1 vssd1 vccd1 vccd1 _09325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06537_ _06621_/A _06663_/A _06536_/A vssd1 vssd1 vccd1 vccd1 _06544_/B sky130_fd_sc_hd__a21oi_1
XFILLER_166_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09256_ _08297_/A _07903_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09256_/X sky130_fd_sc_hd__mux2_1
X_06468_ _06468_/A _06468_/B vssd1 vssd1 vccd1 vccd1 _06474_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08207_ _08208_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08207_/Y sky130_fd_sc_hd__nor2_1
X_05419_ _10625_/Q _05380_/Y _05383_/X _05461_/D _05418_/X vssd1 vssd1 vccd1 vccd1
+ _05419_/X sky130_fd_sc_hd__a221o_1
X_09187_ _09114_/A _09186_/X _10500_/B vssd1 vssd1 vccd1 vccd1 _09187_/X sky130_fd_sc_hd__o21a_1
X_06399_ _10975_/Q vssd1 vssd1 vccd1 vccd1 _06441_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05497__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08138_ _08139_/A _08139_/B vssd1 vssd1 vccd1 vccd1 _08148_/B sky130_fd_sc_hd__nor2_1
XFILLER_134_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08069_ _06008_/A _08047_/X _08052_/X _08059_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08069_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10100_ _10100_/A _10100_/B _10100_/C vssd1 vssd1 vccd1 vccd1 _10101_/B sky130_fd_sc_hd__nand3_1
XFILLER_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10031_ _10031_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__or2_1
XFILLER_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06121__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05960__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10933_ _10958_/CLK _10933_/D vssd1 vssd1 vccd1 vccd1 _10933_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10864_ _10864_/CLK _10864_/D vssd1 vssd1 vccd1 vccd1 _10864_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_25_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10795_ _10798_/CLK _10795_/D vssd1 vssd1 vccd1 vccd1 _10795_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_55_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10229_ _10202_/X _10203_/X _10226_/X _10228_/Y vssd1 vssd1 vccd1 vccd1 _10246_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_67_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05770_ _05767_/Y _10568_/Q _05769_/Y _08317_/A vssd1 vssd1 vccd1 vccd1 _05770_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_63_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07440_ _07573_/A _07574_/A _07726_/B _07732_/B vssd1 vssd1 vccd1 vccd1 _07717_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07371_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07373_/B sky130_fd_sc_hd__or2_1
X_09110_ _09228_/A _09110_/B vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__and2_2
XFILLER_148_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06322_ _06734_/A _06320_/Y _06321_/A _06318_/X vssd1 vssd1 vccd1 vccd1 _06322_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_31_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09041_ _10577_/Q _08972_/X _08974_/A _09040_/X vssd1 vssd1 vccd1 vccd1 _09041_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07928__A2_N _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06253_ _10615_/Q _06253_/B vssd1 vssd1 vccd1 vccd1 _06253_/X sky130_fd_sc_hd__or2_1
XFILLER_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06184_ _10594_/Q vssd1 vssd1 vccd1 vccd1 _06185_/A sky130_fd_sc_hd__inv_2
XANTENNA__06206__A input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09943_ _09943_/A _09943_/B _09943_/C vssd1 vssd1 vccd1 vccd1 _09944_/B sky130_fd_sc_hd__nor3_1
XFILLER_104_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _09943_/A _09874_/B vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__nor2_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08825_ _08825_/A _08825_/B vssd1 vssd1 vccd1 vccd1 _08841_/A sky130_fd_sc_hd__and2_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05968_ input14/X input49/X input1/X vssd1 vssd1 vccd1 vccd1 _08939_/C sky130_fd_sc_hd__nand3b_2
X_08756_ _10809_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08758_/A sky130_fd_sc_hd__nand2_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07707_ _09969_/A _09969_/B _07706_/X vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__a21oi_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08687_ _08808_/A vssd1 vssd1 vccd1 vccd1 _08688_/A sky130_fd_sc_hd__buf_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05899_ _05388_/A _05904_/A _05295_/A vssd1 vssd1 vccd1 vccd1 _05900_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10398__A _10938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _07715_/D _07638_/B vssd1 vssd1 vccd1 vccd1 _07639_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07569_ _10912_/Q vssd1 vssd1 vccd1 vccd1 _09379_/B sky130_fd_sc_hd__buf_2
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09308_ _09449_/A _09443_/B vssd1 vssd1 vccd1 vccd1 _09396_/A sky130_fd_sc_hd__nand2_2
XFILLER_142_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _10693_/CLK _10583_/Q vssd1 vssd1 vccd1 vccd1 _10580_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09239_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09239_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06116__A _08062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09954__B2 _09882_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05955__A _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10017_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10916_ _10981_/CLK _10916_/D vssd1 vssd1 vccd1 vccd1 _10916_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _10847_/CLK _10847_/D vssd1 vssd1 vccd1 vccd1 _10847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10778_ _10782_/CLK _10778_/D vssd1 vssd1 vccd1 vccd1 _10778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08996__A2 _06212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06940_ _06940_/A _06940_/B vssd1 vssd1 vccd1 vccd1 _07636_/A sky130_fd_sc_hd__xnor2_2
XFILLER_140_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06871_ _06871_/A _06871_/B vssd1 vssd1 vccd1 vccd1 _07799_/A sky130_fd_sc_hd__xnor2_4
XFILLER_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08610_ _10786_/Q _08498_/X _08600_/A _08597_/B _10787_/Q vssd1 vssd1 vccd1 vccd1
+ _08612_/B sky130_fd_sc_hd__a41o_1
X_05822_ _05886_/B vssd1 vssd1 vccd1 vccd1 _05823_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09590_ _09591_/B _09590_/B vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__and2b_1
XFILLER_82_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05753_ _08251_/B vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__clkbuf_2
X_08541_ _08541_/A vssd1 vssd1 vccd1 vccd1 _10768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08472_ _08472_/A vssd1 vssd1 vccd1 vccd1 _10740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05684_ _08327_/A _05684_/B vssd1 vssd1 vccd1 vccd1 _05684_/X sky130_fd_sc_hd__or2_1
XANTENNA__08684__A1 _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09881__B1 _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07423_ _07424_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _07425_/A sky130_fd_sc_hd__and2_1
XFILLER_50_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07354_ _07461_/B _07471_/A _07461_/A vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__o21a_1
XFILLER_148_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06305_ _06305_/A _06374_/B _06305_/C vssd1 vssd1 vccd1 vccd1 _06305_/X sky130_fd_sc_hd__or3_1
XFILLER_164_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07285_ _07285_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07286_/B sky130_fd_sc_hd__and2_1
X_09024_ _10198_/A _08418_/B _09168_/A _10801_/Q _08999_/X vssd1 vssd1 vccd1 vccd1
+ _09024_/X sky130_fd_sc_hd__a221o_1
X_06236_ _10608_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06236_/X sky130_fd_sc_hd__or2_1
XFILLER_85_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06167_ input45/X vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__buf_4
XANTENNA__07947__A0 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06098_ _10688_/Q _10687_/Q _08132_/B vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__or3_1
XFILLER_172_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09926_ _10068_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__nand2_1
XFILLER_104_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07990__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _09930_/B _09919_/B _09930_/C _09716_/A vssd1 vssd1 vccd1 vccd1 _09858_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _08808_/A vssd1 vssd1 vccd1 vccd1 _08814_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09787_/A _09787_/B _09787_/C vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__o21ai_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _08688_/X _08736_/X _08738_/X vssd1 vssd1 vccd1 vccd1 _10806_/D sky130_fd_sc_hd__o21a_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10701_ _10703_/CLK _10701_/D vssd1 vssd1 vccd1 vccd1 _10701_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _10666_/CLK _10632_/D vssd1 vssd1 vccd1 vccd1 _10632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10563_ _10674_/CLK _10563_/D vssd1 vssd1 vccd1 vccd1 _10563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _06168_/X _10489_/B _10493_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10970_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10473__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09091__A1 _07393_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07070_ _07070_/A _07070_/B vssd1 vssd1 vccd1 vccd1 _07283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06021_ _08201_/A vssd1 vssd1 vccd1 vccd1 _08837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07972_ _07995_/A vssd1 vssd1 vccd1 vccd1 _08027_/B sky130_fd_sc_hd__buf_2
X_09711_ _09711_/A _09711_/B vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__nor2_1
X_06923_ _06913_/A _06923_/B vssd1 vssd1 vccd1 vccd1 _06923_/X sky130_fd_sc_hd__and2b_1
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09642_ _09642_/A vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06854_ _07675_/A _07780_/B vssd1 vssd1 vccd1 vccd1 _06855_/B sky130_fd_sc_hd__or2_1
XFILLER_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05805_ _05783_/X _05804_/X _05770_/X vssd1 vssd1 vccd1 vccd1 _05805_/X sky130_fd_sc_hd__o21ba_1
XFILLER_27_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09573_ _09567_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09631_/A sky130_fd_sc_hd__and2b_1
X_06785_ _06785_/A vssd1 vssd1 vccd1 vccd1 _10506_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _08524_/A vssd1 vssd1 vccd1 vccd1 _10763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05736_ _05736_/A _10541_/Q vssd1 vssd1 vccd1 vccd1 _05742_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09530__A _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10464__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05667_ _05662_/X _05665_/X _05666_/X vssd1 vssd1 vccd1 vccd1 _05667_/X sky130_fd_sc_hd__a21o_1
X_08455_ _10773_/Q _10736_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08456_/B sky130_fd_sc_hd__mux2_1
X_07406_ _07406_/A vssd1 vssd1 vccd1 vccd1 _07543_/A sky130_fd_sc_hd__inv_2
XFILLER_51_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08386_ _08395_/A _10751_/Q vssd1 vssd1 vccd1 vccd1 _08386_/X sky130_fd_sc_hd__or2_1
XFILLER_149_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05598_ _08251_/A vssd1 vssd1 vccd1 vccd1 _05598_/X sky130_fd_sc_hd__buf_2
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ _07522_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07525_/B sky130_fd_sc_hd__nand2_1
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07268_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07330_/A sky130_fd_sc_hd__xnor2_1
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09007_ _09124_/C _09098_/B vssd1 vssd1 vccd1 vccd1 _10432_/C sky130_fd_sc_hd__nor2_2
X_06219_ input24/X _06207_/X _06218_/X _06200_/X vssd1 vssd1 vccd1 vccd1 _10601_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_151_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07199_ _07277_/A _07277_/B vssd1 vssd1 vccd1 vccd1 _07301_/A sky130_fd_sc_hd__or2b_1
XFILLER_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09909_ _09910_/A _10049_/C vssd1 vssd1 vccd1 vccd1 _09911_/A sky130_fd_sc_hd__or2_1
XFILLER_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08345__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10455__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10615_ _10864_/CLK _10615_/D vssd1 vssd1 vccd1 vccd1 _10615_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09073__A1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__B2 _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10546_ _10654_/CLK _10546_/D vssd1 vssd1 vccd1 vccd1 _10546_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_4_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10477_ _10493_/B vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__08033__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06023__B _06023_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06570_ _06570_/A _06570_/B vssd1 vssd1 vccd1 vccd1 _06599_/A sky130_fd_sc_hd__xnor2_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05521_ _05326_/X _05517_/X _05471_/X _07919_/A vssd1 vssd1 vccd1 vccd1 _10569_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08240_ _08238_/X _08240_/B vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05452_ _05452_/A vssd1 vssd1 vccd1 vccd1 _09107_/A sky130_fd_sc_hd__buf_2
XFILLER_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08171_ _08158_/X _08150_/A _08148_/B _05692_/A vssd1 vssd1 vccd1 vccd1 _08171_/X
+ sky130_fd_sc_hd__a31o_1
X_05383_ _05383_/A _05383_/B vssd1 vssd1 vccd1 vccd1 _05383_/X sky130_fd_sc_hd__and2_1
XANTENNA__09064__B2 _05728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07122_ _07135_/A _07136_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07123_/B sky130_fd_sc_hd__o21bai_4
XFILLER_106_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07053_ _10985_/Q vssd1 vssd1 vccd1 vccd1 _07151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06004_ input38/X _10578_/Q _06120_/S vssd1 vssd1 vccd1 vccd1 _06005_/B sky130_fd_sc_hd__mux2_1
XFILLER_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_opt_6_0_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07955_ _07955_/A _07955_/B vssd1 vssd1 vccd1 vccd1 _07956_/A sky130_fd_sc_hd__or2_1
X_06906_ _06921_/A _06921_/B vssd1 vssd1 vccd1 vccd1 _06906_/X sky130_fd_sc_hd__and2_1
XFILLER_96_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07886_ _10603_/Q _07870_/X _07874_/X _07885_/Y vssd1 vssd1 vccd1 vccd1 _07887_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09625_ _09625_/A _09625_/B _09566_/A vssd1 vssd1 vccd1 vccd1 _09682_/B sky130_fd_sc_hd__or3b_1
X_06837_ _06828_/A _06828_/B _06836_/Y _06796_/B _06796_/A vssd1 vssd1 vccd1 vccd1
+ _06839_/B sky130_fd_sc_hd__o32a_1
XFILLER_71_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09556_ _09554_/C _09600_/A vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__and2b_1
XFILLER_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06768_ _06774_/B vssd1 vssd1 vccd1 vccd1 _06842_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09260__A _09260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10437__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08507_ _10789_/Q _08506_/X _08502_/X _10752_/Q vssd1 vssd1 vccd1 vccd1 _10752_/D
+ sky130_fd_sc_hd__a22o_1
X_05719_ _05719_/A vssd1 vssd1 vccd1 vccd1 _08082_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09487_ _09487_/A vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06699_ _06916_/A _06912_/B _06698_/X vssd1 vssd1 vccd1 vccd1 _06903_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08438_ _10768_/Q _10731_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08439_/B sky130_fd_sc_hd__mux2_1
XFILLER_169_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09055__A1 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10251_/S sky130_fd_sc_hd__buf_2
XFILLER_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10400_ _10537_/A _10399_/X _10395_/X vssd1 vssd1 vccd1 vccd1 _10400_/X sky130_fd_sc_hd__a21bo_1
XFILLER_165_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10331_ _09379_/B _10283_/X _10330_/Y _10293_/X vssd1 vssd1 vccd1 vccd1 _10912_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _07083_/A _10115_/X _10261_/X _10043_/X vssd1 vssd1 vccd1 vccd1 _10905_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06124__A _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10193_ _09634_/A _10198_/B _10192_/X _07394_/X vssd1 vssd1 vccd1 vccd1 _10898_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_78_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06041__A1 _08105_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10428__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput13 io_wbs_m2s_addr[7] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_6
Xinput24 io_wbs_m2s_data[17] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_4
XFILLER_174_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput35 io_wbs_m2s_data[27] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput46 io_wbs_m2s_data[8] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10529_ _10529_/A vssd1 vssd1 vccd1 vccd1 _10529_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_155_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07740_ _07740_/A _07740_/B vssd1 vssd1 vccd1 vccd1 _07741_/B sky130_fd_sc_hd__xnor2_2
XFILLER_96_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07671_ _07671_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07673_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09410_ _10966_/Q _10965_/Q _09443_/B _09411_/A vssd1 vssd1 vccd1 vccd1 _09494_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06622_ _06663_/A _06622_/B _06692_/A _06692_/B vssd1 vssd1 vccd1 vccd1 _06650_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10419__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09341_ _10893_/Q _10909_/Q vssd1 vssd1 vccd1 vccd1 _09343_/A sky130_fd_sc_hd__and2b_1
X_06553_ _06346_/A _06346_/B _10497_/A vssd1 vssd1 vccd1 vccd1 _06555_/A sky130_fd_sc_hd__a21o_1
XFILLER_34_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05504_ _05363_/X _05503_/X _05495_/X _07871_/A vssd1 vssd1 vccd1 vccd1 _10556_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09272_ _09289_/A _09272_/B vssd1 vssd1 vccd1 vccd1 _09273_/A sky130_fd_sc_hd__and2_2
XFILLER_61_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06484_ _06458_/A _06458_/B _06647_/A _06453_/A vssd1 vssd1 vccd1 vccd1 _06486_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__06209__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05435_ _10639_/Q _05340_/X _05434_/X vssd1 vssd1 vccd1 vccd1 _05435_/X sky130_fd_sc_hd__o21a_1
XFILLER_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08223_ _08157_/X _08219_/X _08221_/Y _08222_/X vssd1 vssd1 vccd1 vccd1 _10696_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08245__C1 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ input47/X _08123_/X _08109_/X _08150_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08155_/B sky130_fd_sc_hd__o221a_1
X_05366_ _08198_/A _05369_/A vssd1 vssd1 vccd1 vccd1 _05366_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_147_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ _10985_/Q _07394_/A vssd1 vssd1 vccd1 vccd1 _07137_/C sky130_fd_sc_hd__nand2_1
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08085_ _05279_/A _08043_/A _08080_/Y _06117_/C _08084_/X vssd1 vssd1 vccd1 vccd1
+ _08090_/A sky130_fd_sc_hd__a221o_1
X_05297_ _10658_/Q _06039_/A _05383_/A vssd1 vssd1 vccd1 vccd1 _05373_/B sky130_fd_sc_hd__or3_1
XFILLER_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07036_ _07555_/B _07037_/B vssd1 vssd1 vccd1 vccd1 _07428_/B sky130_fd_sc_hd__or2_1
XFILLER_162_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09255__A _09255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08987_ _09211_/B vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_87_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07938_ _09154_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07939_/A sky130_fd_sc_hd__or2_1
XFILLER_169_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07869_ _10577_/Q _07910_/A vssd1 vssd1 vccd1 vccd1 _07906_/A sky130_fd_sc_hd__and2b_2
XFILLER_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06326__A2 _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09608_ _09608_/A _09608_/B vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__xnor2_4
XFILLER_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10880_ _10881_/CLK _10880_/D vssd1 vssd1 vccd1 vccd1 _10880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09539_ _09596_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__or2_1
XANTENNA__08318__B _08352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06119__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05958__A _10531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08787__B1 _08786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10314_ _10944_/Q _10960_/Q vssd1 vssd1 vccd1 vccd1 _10316_/A sky130_fd_sc_hd__and2b_1
XFILLER_125_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10245_ _10245_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10252_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09200__B2 _10727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10176_ _07061_/A _10174_/X _10170_/X _10888_/Q vssd1 vssd1 vccd1 vccd1 _10888_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_51_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09503__A2 _09879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08509__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10282__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09019__A1 _08998_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_155_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08910_ _09153_/A _08910_/B vssd1 vssd1 vccd1 vccd1 _10827_/D sky130_fd_sc_hd__nor2_1
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09889_/B _09890_/B vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__and2b_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08841_/A _08841_/B _08841_/C vssd1 vssd1 vccd1 vccd1 _08871_/A sky130_fd_sc_hd__and3_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08772_ _10811_/Q _08796_/B vssd1 vssd1 vccd1 vccd1 _08773_/B sky130_fd_sc_hd__or2_1
X_05984_ _05482_/X _05975_/X _05982_/Y _05983_/X vssd1 vssd1 vccd1 vccd1 _10574_/D
+ sky130_fd_sc_hd__a211o_1
X_07723_ _07555_/B _07556_/A _07418_/Y vssd1 vssd1 vccd1 vccd1 _07724_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07654_ _07654_/A _07654_/B vssd1 vssd1 vccd1 vccd1 _09483_/A sky130_fd_sc_hd__nand2_2
XFILLER_93_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06605_ _06607_/C _06605_/B vssd1 vssd1 vccd1 vccd1 _06680_/B sky130_fd_sc_hd__or2_1
X_07585_ _07585_/A _07721_/A vssd1 vssd1 vccd1 vccd1 _07586_/B sky130_fd_sc_hd__xor2_2
XFILLER_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09324_ _09402_/A _09324_/B vssd1 vssd1 vccd1 vccd1 _09326_/B sky130_fd_sc_hd__nand2_1
X_06536_ _06536_/A _06536_/B vssd1 vssd1 vccd1 vccd1 _06663_/A sky130_fd_sc_hd__nor2_2
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09255_ _09255_/A vssd1 vssd1 vccd1 vccd1 _10857_/D sky130_fd_sc_hd__clkbuf_1
X_06467_ _06456_/A _06460_/B _06917_/A vssd1 vssd1 vccd1 vccd1 _06468_/B sky130_fd_sc_hd__a21boi_1
XFILLER_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08206_ _08206_/A vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__buf_2
XFILLER_154_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05418_ _10624_/Q _05383_/X _05385_/Y _05462_/A _05417_/X vssd1 vssd1 vccd1 vccd1
+ _05418_/X sky130_fd_sc_hd__o221a_1
XFILLER_166_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06398_ _06456_/A vssd1 vssd1 vccd1 vccd1 _06626_/A sky130_fd_sc_hd__clkbuf_2
X_09186_ _10945_/Q _09143_/Y _09185_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09186_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_147_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05349_ _10635_/Q vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10834__D _10834_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08137_ _08150_/B _08136_/Y _08062_/A vssd1 vssd1 vccd1 vccd1 _08137_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07993__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08068_ _08075_/B _08072_/B _08067_/X _06033_/X vssd1 vssd1 vccd1 vccd1 _08068_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_162_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07019_ _07472_/A _07434_/A _07416_/A vssd1 vssd1 vccd1 vccd1 _07035_/A sky130_fd_sc_hd__and3b_1
X_10030_ _10031_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10030_/X sky130_fd_sc_hd__and2_1
XFILLER_89_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10932_ _10935_/CLK _10932_/D vssd1 vssd1 vccd1 vccd1 _10932_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10863_ _10863_/CLK _10863_/D vssd1 vssd1 vccd1 vccd1 _10863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _10798_/CLK _10794_/D vssd1 vssd1 vccd1 vccd1 _10794_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06235__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06015__C input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10228_ _10228_/A vssd1 vssd1 vccd1 vccd1 _10228_/Y sky130_fd_sc_hd__inv_2
XFILLER_95_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__xnor2_4
XFILLER_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08696__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07370_ _07412_/C _07370_/B vssd1 vssd1 vccd1 vccd1 _07374_/A sky130_fd_sc_hd__nor2_2
XANTENNA__06982__A _07747_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06321_ _06321_/A _06320_/Y vssd1 vssd1 vccd1 vccd1 _06735_/A sky130_fd_sc_hd__or2b_2
X_06252_ input39/X _06145_/B _06251_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10614_/D
+ sky130_fd_sc_hd__o211a_1
X_09040_ _05279_/A _08995_/X _09039_/X _08981_/A vssd1 vssd1 vccd1 vccd1 _09040_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_164_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06183_ _06204_/B vssd1 vssd1 vccd1 vccd1 _06183_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _09943_/A _09943_/B _09943_/C vssd1 vssd1 vccd1 vccd1 _10012_/A sky130_fd_sc_hd__o21a_1
XFILLER_86_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09874_/B sky130_fd_sc_hd__and2_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08824_ hold3/A _08856_/B vssd1 vssd1 vccd1 vccd1 _08825_/B sky130_fd_sc_hd__or2_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09533__A _10967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08755_ _08688_/X _08753_/Y _08754_/X vssd1 vssd1 vccd1 vccd1 _10808_/D sky130_fd_sc_hd__o21a_1
X_05967_ input15/X input6/X input5/X vssd1 vssd1 vccd1 vccd1 _08414_/A sky130_fd_sc_hd__or3_2
XFILLER_54_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07706_ _07610_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _07706_/X sky130_fd_sc_hd__and2b_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _08686_/A _08819_/A vssd1 vssd1 vccd1 vccd1 _08808_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_32_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10666_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05898_ _06038_/A _05906_/A vssd1 vssd1 vccd1 vccd1 _05904_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07053__A _10985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07637_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__xnor2_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07988__A _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07568_ _07726_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__nand2_1
XFILLER_167_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09307_ _09387_/A vssd1 vssd1 vccd1 vccd1 _09443_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_47_clock clkbuf_opt_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _10862_/CLK sky130_fd_sc_hd__clkbuf_16
X_06519_ _06519_/A _06519_/B vssd1 vssd1 vccd1 vccd1 _06523_/C sky130_fd_sc_hd__nor2_1
XFILLER_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07499_ _07499_/A _07499_/B vssd1 vssd1 vccd1 vccd1 _07504_/A sky130_fd_sc_hd__xnor2_1
XFILLER_166_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09238_ _08268_/A _09237_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09238_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09169_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06217__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08612__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10013_ _10081_/B _10013_/B vssd1 vssd1 vccd1 vccd1 _10015_/B sky130_fd_sc_hd__or2_1
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09443__A _10967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input22_A io_wbs_m2s_data[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08142__A1 _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10915_ _10981_/CLK _10915_/D vssd1 vssd1 vccd1 vccd1 _10915_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10846_ _10848_/CLK _10846_/D vssd1 vssd1 vccd1 vccd1 _10846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10777_ _10782_/CLK _10777_/D vssd1 vssd1 vccd1 vccd1 _10777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06870_ _07761_/A _07761_/B vssd1 vssd1 vccd1 vccd1 _06871_/B sky130_fd_sc_hd__xnor2_2
XFILLER_68_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05821_ _05906_/A vssd1 vssd1 vccd1 vccd1 _05886_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08540_ _08543_/B _08580_/B _08540_/C vssd1 vssd1 vccd1 vccd1 _08541_/A sky130_fd_sc_hd__and3b_1
XFILLER_48_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05752_ _10560_/Q vssd1 vssd1 vccd1 vccd1 _05752_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08133__B2 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08471_ _08477_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _08472_/A sky130_fd_sc_hd__or2_1
X_05683_ _08317_/A _05583_/Y _05684_/B _08327_/A vssd1 vssd1 vccd1 vccd1 _05683_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ _07421_/Y _07043_/A _07417_/A _07044_/A vssd1 vssd1 vccd1 vccd1 _07424_/B
+ sky130_fd_sc_hd__o211a_1
X_07353_ _07369_/B _07353_/B vssd1 vssd1 vccd1 vccd1 _07461_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06304_ _06304_/A _06304_/B vssd1 vssd1 vccd1 vccd1 _06374_/B sky130_fd_sc_hd__nand2_2
XFILLER_109_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07284_ _07284_/A _07284_/B vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__and2_1
XFILLER_148_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09023_ _10578_/Q _08972_/X _08974_/X _09022_/X vssd1 vssd1 vccd1 vccd1 _09023_/X
+ sky130_fd_sc_hd__o211a_1
X_06235_ input31/X _06225_/X _06233_/X _06234_/X vssd1 vssd1 vccd1 vccd1 _10607_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06166_ _06163_/X _06158_/X _06165_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10590_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07947__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06097_ _10686_/Q _08117_/B vssd1 vssd1 vccd1 vccd1 _08132_/B sky130_fd_sc_hd__or2_1
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09925_ _09925_/A _09925_/B vssd1 vssd1 vccd1 vccd1 _10141_/B sky130_fd_sc_hd__xnor2_4
XFILLER_120_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _10484_/A _09930_/C _09856_/C vssd1 vssd1 vccd1 vccd1 _10076_/A sky130_fd_sc_hd__nand3_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09263__A _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08807_ _08801_/X _08802_/Y _08804_/Y _08806_/Y vssd1 vssd1 vccd1 vccd1 _08810_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09787_/A _09787_/B _09787_/C vssd1 vssd1 vccd1 vccd1 _09848_/B sky130_fd_sc_hd__or3_1
XFILLER_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06999_ _07007_/A _07570_/C vssd1 vssd1 vccd1 vccd1 _07000_/B sky130_fd_sc_hd__nand2_1
XFILLER_74_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _10537_/A _08694_/X _08695_/X _10806_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08738_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10202__A _10933_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _10799_/Q _08669_/B _08669_/C vssd1 vssd1 vccd1 vccd1 _08670_/C sky130_fd_sc_hd__nand3_1
XFILLER_82_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ _10703_/CLK _10700_/D vssd1 vssd1 vccd1 vccd1 _10700_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10631_ _10814_/CLK _10631_/D vssd1 vssd1 vccd1 vccd1 _10631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10562_ _10562_/CLK _10562_/D vssd1 vssd1 vccd1 vccd1 _10562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06127__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10493_ _10493_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10493_/X sky130_fd_sc_hd__or2_1
XFILLER_6_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08342__A _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_3_0_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_0_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_92_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08517__A _10177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10829_ _10830_/CLK _10829_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09076__C1 _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06020_ _08258_/A vssd1 vssd1 vccd1 vccd1 _06020_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_133_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07971_ _10517_/A _09263_/A vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09710_ _09710_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09711_/B sky130_fd_sc_hd__and2_1
X_06922_ _06922_/A _06922_/B vssd1 vssd1 vccd1 vccd1 _06926_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08354__A1 _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08354__B2 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09641_ _09641_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__xor2_2
X_06853_ _06853_/A _06853_/B vssd1 vssd1 vccd1 vccd1 _07780_/B sky130_fd_sc_hd__nor2_1
XFILLER_56_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05804_ _08321_/A _05769_/A _10566_/Q _05781_/Y vssd1 vssd1 vccd1 vccd1 _05804_/X
+ sky130_fd_sc_hd__a22o_1
X_09572_ _10115_/A vssd1 vssd1 vccd1 vccd1 _09572_/X sky130_fd_sc_hd__clkbuf_2
X_06784_ _06828_/A _06828_/B vssd1 vssd1 vccd1 vccd1 _06882_/A sky130_fd_sc_hd__or2_1
X_08523_ _08935_/A _10762_/Q vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__and2_1
XANTENNA__09811__A _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05735_ _08093_/A _05547_/A _05536_/B _05733_/X _05734_/X vssd1 vssd1 vccd1 vccd1
+ _05788_/B sky130_fd_sc_hd__o221ai_2
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08454_ _08454_/A vssd1 vssd1 vccd1 vccd1 _10735_/D sky130_fd_sc_hd__clkbuf_1
X_05666_ _10693_/Q _05664_/Y _05615_/Y _05877_/A vssd1 vssd1 vccd1 vccd1 _05666_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07405_ _07405_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _07540_/A sky130_fd_sc_hd__or2_1
XFILLER_51_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08409__A2 _10744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08385_ _10198_/A vssd1 vssd1 vccd1 vccd1 _08395_/A sky130_fd_sc_hd__clkbuf_1
X_05597_ _10700_/Q vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07336_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07522_/B sky130_fd_sc_hd__and2_1
XFILLER_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07267_ _07268_/A _07268_/B vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__or2_1
XANTENNA__07985__B _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09006_ _10069_/A vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__buf_2
X_06218_ hold6/A _06223_/B vssd1 vssd1 vccd1 vccd1 _06218_/X sky130_fd_sc_hd__or2_1
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07198_ _07193_/A _07193_/B _07194_/B _07210_/A _07260_/A vssd1 vssd1 vccd1 vccd1
+ _07277_/B sky130_fd_sc_hd__a32o_1
XFILLER_117_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10842__D _10842_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06149_ _06149_/A vssd1 vssd1 vccd1 vccd1 _06238_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_133_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09908_ _09908_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _10049_/C sky130_fd_sc_hd__nand2_2
XFILLER_59_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08345__A1 input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08345__B2 _05570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09839_ _09974_/A _09839_/B _09839_/C vssd1 vssd1 vccd1 vccd1 _09841_/A sky130_fd_sc_hd__and3_1
XFILLER_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10614_ _10864_/CLK _10614_/D vssd1 vssd1 vccd1 vccd1 _10614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ _10545_/CLK _10545_/D vssd1 vssd1 vccd1 vccd1 _10545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10476_ _10517_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10493_/B sky130_fd_sc_hd__nor2_1
XFILLER_108_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10391__A1 _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07416__A _07416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05520_ _05329_/X _05517_/X _05513_/X _07914_/A vssd1 vssd1 vccd1 vccd1 _10568_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05451_ _10620_/Q vssd1 vssd1 vccd1 vccd1 _05453_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_46_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08170_ _08180_/B vssd1 vssd1 vccd1 vccd1 _08181_/B sky130_fd_sc_hd__inv_2
XFILLER_174_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05382_ _10656_/Q _05382_/B vssd1 vssd1 vccd1 vccd1 _05383_/B sky130_fd_sc_hd__nand2_1
X_07121_ _07145_/A _07145_/B vssd1 vssd1 vccd1 vccd1 _07136_/A sky130_fd_sc_hd__and2b_1
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07052_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07373_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09078__A _09078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06003_ _06003_/A vssd1 vssd1 vccd1 vccd1 _10577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07954_ input43/X _06038_/X _07983_/A vssd1 vssd1 vccd1 vccd1 _07955_/B sky130_fd_sc_hd__mux2_1
XFILLER_101_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06905_ _06567_/B _06368_/B _06895_/B vssd1 vssd1 vccd1 vccd1 _06922_/B sky130_fd_sc_hd__a21oi_2
XFILLER_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07885_ _07885_/A vssd1 vssd1 vccd1 vccd1 _07885_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09624_ _09624_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__and2_1
XFILLER_83_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06836_ _06836_/A vssd1 vssd1 vccd1 vccd1 _06836_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09555_ _09555_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__nand2_1
X_06767_ _06775_/A vssd1 vssd1 vccd1 vccd1 _06900_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08506_ _08514_/A vssd1 vssd1 vccd1 vccd1 _08506_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05718_ _05718_/A vssd1 vssd1 vccd1 vccd1 _08082_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _09486_/A _09486_/B vssd1 vssd1 vccd1 vccd1 _09562_/A sky130_fd_sc_hd__xnor2_1
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06698_ _06697_/B _06698_/B vssd1 vssd1 vccd1 vccd1 _06698_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08157__A _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07061__A _07061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10837__D _10837_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _08437_/A vssd1 vssd1 vccd1 vccd1 _10730_/D sky130_fd_sc_hd__clkbuf_1
X_05649_ _05719_/A _05641_/Y _05648_/X vssd1 vssd1 vccd1 vccd1 _05649_/X sky130_fd_sc_hd__a21o_1
XFILLER_12_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07996__A _08209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08368_ _10729_/Q vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07319_ _07319_/A _07319_/B vssd1 vssd1 vccd1 vccd1 _07341_/B sky130_fd_sc_hd__or2_1
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08299_ _08305_/B _08253_/X _08297_/Y _08298_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08299_/X sky130_fd_sc_hd__a311o_1
XFILLER_20_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10330_ _10330_/A _10330_/B vssd1 vssd1 vccd1 vccd1 _10330_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10261_ _10261_/A _10261_/B vssd1 vssd1 vccd1 vccd1 _10261_/X sky130_fd_sc_hd__xor2_2
XFILLER_133_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10192_ _10192_/A vssd1 vssd1 vccd1 vccd1 _10192_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_106_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06041__A2 _06038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08067__A _08092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 io_wbs_m2s_addr[8] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
XFILLER_122_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08254__B1 _05598_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput25 io_wbs_m2s_data[18] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_4
Xinput36 io_wbs_m2s_data[28] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_4
Xinput47 io_wbs_m2s_data[9] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_4
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10528_ _10528_/A _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10528_/X sky130_fd_sc_hd__or3_1
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10459_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10459_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_130_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10116__A1 _10109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07670_ _07670_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07671_/B sky130_fd_sc_hd__nand2_1
XFILLER_93_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06621_ _06621_/A _06621_/B vssd1 vssd1 vccd1 vccd1 _06692_/B sky130_fd_sc_hd__nor2_2
XFILLER_92_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09340_ _06993_/A _10894_/Q vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__and2b_1
X_06552_ _10971_/Q vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__clkinv_2
XFILLER_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05503_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05503_/X sky130_fd_sc_hd__clkbuf_1
X_09271_ _10825_/Q _09243_/X _09244_/X _09269_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09272_/B sky130_fd_sc_hd__a32o_1
XFILLER_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06483_ _06646_/A _06646_/B vssd1 vssd1 vccd1 vccd1 _06647_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08222_ input23/X _08164_/X _08165_/X _08216_/X _08394_/A vssd1 vssd1 vccd1 vccd1
+ _08222_/X sky130_fd_sc_hd__o221a_1
X_05434_ _07896_/A _05343_/Y _05431_/X _05433_/X vssd1 vssd1 vccd1 vccd1 _05434_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08153_ _07976_/A _08043_/A _08152_/X _08038_/A _08096_/A vssd1 vssd1 vccd1 vccd1
+ _08155_/A sky130_fd_sc_hd__a221o_1
XFILLER_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05365_ _10662_/Q vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_147_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07104_ _07142_/B vssd1 vssd1 vccd1 vccd1 _07394_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08084_ _08113_/A _08081_/X _08083_/Y _06024_/A vssd1 vssd1 vccd1 vccd1 _08084_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06225__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05296_ _10656_/Q _05382_/B vssd1 vssd1 vccd1 vccd1 _05383_/A sky130_fd_sc_hd__or2_1
XFILLER_162_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07035_ _07035_/A _07415_/C vssd1 vssd1 vccd1 vccd1 _07037_/B sky130_fd_sc_hd__xor2_1
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09536__A _10969_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__and2_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07937_ input16/X _05475_/X _07964_/A vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__mux2_1
XFILLER_130_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07868_ _07848_/X _05460_/B _07865_/X _07867_/Y vssd1 vssd1 vccd1 vccd1 _10630_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09607_ _09607_/A _09676_/D vssd1 vssd1 vccd1 vccd1 _09608_/B sky130_fd_sc_hd__xor2_4
XFILLER_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06819_ _10502_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _07779_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07799_ _07799_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _07799_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09538_ _09538_/A _09638_/C vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__and2_1
XFILLER_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09469_ _09534_/C _09469_/B vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08787__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10313_ _09920_/B _10283_/X _10312_/X _10293_/X vssd1 vssd1 vccd1 vccd1 _10910_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10244_ _10953_/Q _10937_/Q vssd1 vssd1 vccd1 vccd1 _10245_/B sky130_fd_sc_hd__and2b_1
XFILLER_152_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10175_ _07066_/A _10174_/X _10170_/X _10887_/Q vssd1 vssd1 vccd1 vccd1 _10887_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08711__A1 _10533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09019__A2 _09001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08244__B _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09356__A _09356_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _10819_/Q _08840_/B vssd1 vssd1 vccd1 vccd1 _08844_/A sky130_fd_sc_hd__xnor2_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08771_ _08771_/A _08796_/B vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__nand2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05983_ _08445_/A vssd1 vssd1 vccd1 vccd1 _05983_/X sky130_fd_sc_hd__clkbuf_8
XFILLER_111_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07722_ _07585_/A _07721_/Y _07584_/A vssd1 vssd1 vccd1 vccd1 _07741_/A sky130_fd_sc_hd__a21oi_1
XFILLER_84_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07653_ _07653_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07654_/B sky130_fd_sc_hd__nand2_1
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06604_ _06593_/A _06593_/B _06593_/C vssd1 vssd1 vccd1 vccd1 _06605_/B sky130_fd_sc_hd__a21oi_1
X_07584_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07721_/A sky130_fd_sc_hd__or2_1
XFILLER_53_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09323_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09324_/B sky130_fd_sc_hd__or2_1
X_06535_ _06534_/B _06535_/B vssd1 vssd1 vccd1 vccd1 _06536_/B sky130_fd_sc_hd__and2b_1
XFILLER_34_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09254_ _09259_/A _09254_/B vssd1 vssd1 vccd1 vccd1 _09255_/A sky130_fd_sc_hd__and2_4
XFILLER_139_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06466_ _06480_/C _06466_/B vssd1 vssd1 vccd1 vccd1 _06688_/A sky130_fd_sc_hd__or2_1
X_08205_ _08206_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08224_/C sky130_fd_sc_hd__and2_1
XFILLER_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05417_ _05462_/B _05389_/Y _05385_/Y _10623_/Q _05416_/X vssd1 vssd1 vccd1 vccd1
+ _05417_/X sky130_fd_sc_hd__a221o_1
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09185_ _10961_/Q _09194_/B vssd1 vssd1 vccd1 vccd1 _09185_/Y sky130_fd_sc_hd__nor2_1
X_06397_ _10977_/Q vssd1 vssd1 vccd1 vccd1 _06456_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_135_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08136_ _08132_/A _08132_/B _06035_/A vssd1 vssd1 vccd1 vccd1 _08136_/Y sky130_fd_sc_hd__o21ai_1
X_05348_ _05854_/A _05348_/B vssd1 vssd1 vccd1 vccd1 _05348_/X sky130_fd_sc_hd__and2_1
XFILLER_174_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08067_ _08092_/A vssd1 vssd1 vccd1 vccd1 _08067_/X sky130_fd_sc_hd__buf_2
X_05279_ _05279_/A vssd1 vssd1 vccd1 vccd1 _05818_/A sky130_fd_sc_hd__inv_2
X_07018_ _07229_/A vssd1 vssd1 vccd1 vccd1 _07416_/A sky130_fd_sc_hd__buf_2
XFILLER_122_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08969_ _09142_/B _09142_/C _08965_/B _08968_/X vssd1 vssd1 vccd1 vccd1 _08969_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_29_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09205__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10931_ _10935_/CLK _10931_/D vssd1 vssd1 vccd1 vccd1 _10931_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10862_ _10862_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _10862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ _10798_/CLK _10793_/D vssd1 vssd1 vccd1 vccd1 _10793_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10227_ _10226_/B _10217_/X _10214_/A vssd1 vssd1 vccd1 vccd1 _10228_/A sky130_fd_sc_hd__a21o_1
XFILLER_95_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10115__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10158_ _10158_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__xnor2_2
XFILLER_95_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_94_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10089_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10090_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06171__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06320_ _10924_/Q _10907_/Q vssd1 vssd1 vccd1 vccd1 _06320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_149_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06251_ _10614_/Q _06253_/B vssd1 vssd1 vccd1 vccd1 _06251_/X sky130_fd_sc_hd__or2_1
XFILLER_129_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09948__B1 _10493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06182_ input17/X vssd1 vssd1 vccd1 vccd1 _06182_/X sky130_fd_sc_hd__buf_4
XFILLER_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09941_ _10009_/B _09941_/B vssd1 vssd1 vccd1 vccd1 _09943_/C sky130_fd_sc_hd__and2_1
XFILLER_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10025__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09943_/A sky130_fd_sc_hd__nor2_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10682__CLK _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08823_ hold3/X _08865_/B vssd1 vssd1 vccd1 vccd1 _08825_/A sky130_fd_sc_hd__nand2_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08754_ _06178_/X _08694_/X _08695_/X _10808_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08754_/X sky130_fd_sc_hd__o221a_1
X_05966_ _09016_/A _09126_/A vssd1 vssd1 vccd1 vccd1 _08965_/A sky130_fd_sc_hd__or2_2
X_07705_ _07616_/X _09899_/B _07704_/Y vssd1 vssd1 vccd1 vccd1 _09969_/B sky130_fd_sc_hd__a21bo_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08683_/X _08684_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10801_/D sky130_fd_sc_hd__o21a_1
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05897_ _10656_/Q _05900_/A vssd1 vssd1 vccd1 vccd1 _05897_/X sky130_fd_sc_hd__xor2_1
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _07636_/A _07636_/B vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__xor2_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07567_ _07567_/A vssd1 vssd1 vccd1 vccd1 _07726_/A sky130_fd_sc_hd__buf_2
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09306_ _09306_/A _09316_/A vssd1 vssd1 vccd1 vccd1 _09387_/A sky130_fd_sc_hd__or2_1
X_06518_ _06521_/A _06521_/B _06612_/A _06503_/Y vssd1 vssd1 vccd1 vccd1 _06519_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_167_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07498_ _07534_/B _07534_/C _07534_/A vssd1 vssd1 vccd1 vccd1 _07535_/A sky130_fd_sc_hd__o21a_1
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08165__A _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _08267_/A _07893_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09237_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10845__D _10845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06449_ _06472_/A _06470_/A _06426_/A _06568_/B vssd1 vssd1 vccd1 vccd1 _06450_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_21_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09168_ _09168_/A vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08119_ _08119_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08119_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _10493_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _09114_/A sky130_fd_sc_hd__nor2_2
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10580__D _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10012_ _10012_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input15_A io_wbs_m2s_addr[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08059__B _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10914_ _10914_/CLK _10914_/D vssd1 vssd1 vccd1 vccd1 _10914_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10845_ _10847_/CLK _10845_/D vssd1 vssd1 vccd1 vccd1 _10845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10776_ _10776_/CLK _10776_/D vssd1 vssd1 vccd1 vccd1 _10776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09634__A _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05820_ _05905_/A _05905_/B vssd1 vssd1 vccd1 vccd1 _05906_/A sky130_fd_sc_hd__or2_2
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05751_ _10700_/Q vssd1 vssd1 vccd1 vccd1 _05751_/Y sky130_fd_sc_hd__clkinv_2
X_08470_ _10777_/Q _10740_/Q _08473_/S vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__mux2_1
X_05682_ _10707_/Q vssd1 vssd1 vccd1 vccd1 _08327_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__06993__A _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07421_ _07421_/A vssd1 vssd1 vccd1 vccd1 _07421_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07352_ _07366_/B _07291_/B _07291_/C vssd1 vssd1 vccd1 vccd1 _07353_/B sky130_fd_sc_hd__a21oi_1
XFILLER_149_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06303_ _06303_/A _06305_/C vssd1 vssd1 vccd1 vccd1 _06730_/B sky130_fd_sc_hd__or2_1
XFILLER_31_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07283_ _07357_/C _07283_/B vssd1 vssd1 vccd1 vccd1 _07284_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09022_ _06065_/X _08976_/X _09020_/X _09021_/Y _09078_/B vssd1 vssd1 vccd1 vccd1
+ _09022_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06234_ _07977_/A vssd1 vssd1 vccd1 vccd1 _06234_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06165_ _06165_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06096_ _10685_/Q _10684_/Q _08098_/B vssd1 vssd1 vccd1 vccd1 _08117_/B sky130_fd_sc_hd__or3_1
XFILLER_172_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09149__B2 _08160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06080__B1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09924_ _10131_/A _09924_/B vssd1 vssd1 vccd1 vccd1 _09925_/B sky130_fd_sc_hd__nand2_2
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input7_A io_wbs_m2s_addr[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _09855_/A _09855_/B vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__xor2_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08806_ _08806_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _08806_/Y sky130_fd_sc_hd__nor2_1
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09787_/C sky130_fd_sc_hd__xnor2_1
XFILLER_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06998_ _07028_/A _07008_/A _07007_/B vssd1 vssd1 vccd1 vccd1 _07570_/C sky130_fd_sc_hd__or3_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05949_ _08350_/A _05829_/X _05826_/X _05528_/X _05948_/X vssd1 vssd1 vccd1 vccd1
+ _05949_/X sky130_fd_sc_hd__o221a_1
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08737_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08737_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _08669_/B _08669_/C _10799_/Q vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__a21o_1
XFILLER_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07619_ _07625_/A _07624_/B _07624_/A vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__a21oi_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08599_ _09403_/B _08624_/B vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__or2_2
XFILLER_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10630_ _10814_/CLK _10630_/D vssd1 vssd1 vccd1 vccd1 _10630_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05312__A _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10561_ _10671_/CLK _10561_/D vssd1 vssd1 vccd1 vccd1 _10561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10492_ _06163_/X _10489_/B _10491_/X _10485_/X vssd1 vssd1 vccd1 vccd1 _10969_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06143__A _10526_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05949__B2 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05982__A _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08899__B1 _08786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10828_ _10864_/CLK _10828_/D vssd1 vssd1 vccd1 vccd1 _10828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10759_ _10935_/CLK _10759_/D vssd1 vssd1 vccd1 vccd1 _10759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09629__A _09629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08533__A _08881_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_31_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10814_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_141_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06062__B1 _05388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09263_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__06988__A _07563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06921_ _06921_/A _06921_/B vssd1 vssd1 vccd1 vccd1 _06922_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_46_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10859_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_42_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09640_ _09640_/A _09640_/B vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06852_ _06852_/A _06852_/B vssd1 vssd1 vccd1 vccd1 _06855_/A sky130_fd_sc_hd__xor2_2
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05803_ _05803_/A vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__inv_2
X_09571_ _10872_/Q _09408_/X _09570_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10872_/D
+ sky130_fd_sc_hd__a22o_1
X_06783_ _06902_/A _06892_/B _06782_/A vssd1 vssd1 vccd1 vccd1 _06828_/B sky130_fd_sc_hd__a21oi_2
XFILLER_36_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08522_ _08522_/A vssd1 vssd1 vccd1 vccd1 _10762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05734_ _05726_/A _05549_/A _05729_/Y _05728_/X vssd1 vssd1 vccd1 vccd1 _05734_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_24_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08453_ _08460_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08454_/A sky130_fd_sc_hd__or2_1
X_05665_ _05885_/A _05619_/X _05664_/Y _10693_/Q vssd1 vssd1 vccd1 vccd1 _05665_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07404_ _07404_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _07405_/B sky130_fd_sc_hd__and2_1
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08384_ _10251_/S vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__clkbuf_4
X_05596_ _05596_/A _05596_/B vssd1 vssd1 vccd1 vccd1 _05596_/X sky130_fd_sc_hd__and2_1
X_07335_ _07335_/A _07335_/B vssd1 vssd1 vccd1 vccd1 _07511_/B sky130_fd_sc_hd__and2_1
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07266_ _07266_/A _07270_/A vssd1 vssd1 vccd1 vccd1 _07268_/B sky130_fd_sc_hd__xnor2_1
XFILLER_118_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08443__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ _09931_/A vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_118_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06217_ input23/X _06207_/X _06216_/X _06200_/X vssd1 vssd1 vccd1 vccd1 _10600_/D
+ sky130_fd_sc_hd__o211a_1
X_07197_ _07197_/A _07197_/B _07197_/C vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__and3_1
XANTENNA__07059__A _07560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06148_ _10587_/Q vssd1 vssd1 vccd1 vccd1 _06151_/A sky130_fd_sc_hd__inv_2
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06079_ _06113_/A _08342_/A _06038_/X _08105_/A _06078_/X vssd1 vssd1 vccd1 vccd1
+ _06082_/C sky130_fd_sc_hd__a221o_1
XFILLER_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09274__A _09274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ _09907_/A _09907_/B vssd1 vssd1 vccd1 vccd1 _09910_/A sky130_fd_sc_hd__xnor2_1
XFILLER_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08345__A2 _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ _09906_/A _09838_/B vssd1 vssd1 vccd1 vccd1 _09839_/C sky130_fd_sc_hd__and2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09769_ _09769_/A _09769_/B _09769_/C vssd1 vssd1 vccd1 vccd1 _09771_/C sky130_fd_sc_hd__and3_1
XFILLER_74_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10613_ _10864_/CLK _10613_/D vssd1 vssd1 vccd1 vccd1 _10613_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05977__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ _10545_/CLK _10544_/D vssd1 vssd1 vccd1 vccd1 _10544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08281__B2 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10475_ _10489_/B vssd1 vssd1 vccd1 vccd1 _10475_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08033__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06044__B1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10123__A _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09297__A0 _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07432__A _07563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05450_ _05490_/A vssd1 vssd1 vccd1 vccd1 _05470_/A sky130_fd_sc_hd__inv_2
XFILLER_162_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05381_ _10625_/Q vssd1 vssd1 vccd1 vccd1 _05461_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07120_ _07135_/A _07511_/A _07149_/C _07235_/B vssd1 vssd1 vccd1 vccd1 _07145_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08263__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07051_ _07051_/A _07414_/A vssd1 vssd1 vccd1 vccd1 _07371_/B sky130_fd_sc_hd__xnor2_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09509__D _09599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06002_ _08483_/A _06002_/B vssd1 vssd1 vccd1 vccd1 _06003_/A sky130_fd_sc_hd__and2_1
XFILLER_115_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08024__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A0 _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07953_ _07953_/A vssd1 vssd1 vccd1 vccd1 _10652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06904_ _06921_/A _06921_/B vssd1 vssd1 vccd1 vccd1 _06904_/X sky130_fd_sc_hd__or2_1
X_07884_ _07898_/A _07884_/B vssd1 vssd1 vccd1 vccd1 _10634_/D sky130_fd_sc_hd__nor2_1
XFILLER_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ _09623_/A _09623_/B _09623_/C vssd1 vssd1 vccd1 vccd1 _09624_/B sky130_fd_sc_hd__or3_1
X_06835_ _06835_/A _06835_/B vssd1 vssd1 vccd1 vccd1 _06839_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09554_ _09805_/A _09692_/A _09554_/C vssd1 vssd1 vccd1 vccd1 _09652_/A sky130_fd_sc_hd__and3_1
X_06766_ _06766_/A _06766_/B vssd1 vssd1 vccd1 vccd1 _06828_/A sky130_fd_sc_hd__or2_1
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05717_ _05798_/A _05717_/B _05717_/C _05717_/D vssd1 vssd1 vccd1 vccd1 _05717_/X
+ sky130_fd_sc_hd__or4_2
X_08505_ _10788_/Q _08496_/X _08502_/X _10751_/Q vssd1 vssd1 vccd1 vccd1 _10751_/D
+ sky130_fd_sc_hd__a22o_1
X_09485_ _09904_/A _09744_/A vssd1 vssd1 vccd1 vccd1 _09486_/B sky130_fd_sc_hd__nand2_1
X_06697_ _06698_/B _06697_/B vssd1 vssd1 vccd1 vccd1 _06912_/B sky130_fd_sc_hd__xnor2_2
X_05648_ _05719_/A _05641_/Y _05644_/Y _08082_/C _05647_/X vssd1 vssd1 vccd1 vccd1
+ _05648_/X sky130_fd_sc_hd__o221a_1
X_08436_ _08443_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08437_/A sky130_fd_sc_hd__or2_1
XFILLER_169_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08367_ _08419_/A vssd1 vssd1 vccd1 vccd1 _08367_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05579_ _10566_/Q _05588_/A vssd1 vssd1 vccd1 vccd1 _05580_/B sky130_fd_sc_hd__nand2_1
XFILLER_149_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07318_ _07318_/A _07318_/B _07324_/A vssd1 vssd1 vccd1 vccd1 _07319_/B sky130_fd_sc_hd__and3_1
XFILLER_20_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08298_ _08298_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08298_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07926__A2_N _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07249_ _07517_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _07250_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10853__D _10853_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10323__A_N _10945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ _10258_/Y _10259_/X _10291_/S vssd1 vssd1 vccd1 vccd1 _10261_/B sky130_fd_sc_hd__mux2_1
XFILLER_105_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08901__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ _10197_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10198_/B sky130_fd_sc_hd__and2b_1
XFILLER_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06140__B _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08348__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08254__A1 _08242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput15 io_wbs_m2s_addr[9] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_2
XFILLER_128_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput26 io_wbs_m2s_data[19] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_4
Xinput37 io_wbs_m2s_data[29] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_8
Xinput48 io_wbs_m2s_sel[0] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_6
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10527_ _07726_/A _10522_/X _10526_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10981_/D
+ sky130_fd_sc_hd__o211a_2
XANTENNA__06315__B _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ _06178_/X _10446_/X _10456_/X _10457_/X vssd1 vssd1 vccd1 vccd1 _10956_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_171_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10389_ _10408_/A vssd1 vssd1 vccd1 vccd1 _10389_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10521__C1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06620_ _06620_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _06621_/B sky130_fd_sc_hd__and2_1
XFILLER_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06551_ _06561_/B _06561_/C _06587_/B vssd1 vssd1 vccd1 vccd1 _06564_/A sky130_fd_sc_hd__and3_1
XFILLER_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05502_ _05366_/Y _05497_/X _05490_/A _05460_/B vssd1 vssd1 vccd1 vccd1 _10555_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09270_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09270_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06482_ _06658_/A _06657_/B _06657_/A vssd1 vssd1 vccd1 vccd1 _06646_/B sky130_fd_sc_hd__o21ba_1
X_08221_ _08216_/X _08224_/C _08220_/Y vssd1 vssd1 vccd1 vccd1 _08221_/Y sky130_fd_sc_hd__a21oi_1
X_05433_ _10638_/Q _05343_/Y _05348_/X _07893_/A vssd1 vssd1 vccd1 vccd1 _05433_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08152_ _08065_/B _08147_/X _08149_/Y _08151_/Y _08074_/A vssd1 vssd1 vccd1 vccd1
+ _08152_/X sky130_fd_sc_hd__a32o_1
X_05364_ _10630_/Q vssd1 vssd1 vccd1 vccd1 _05460_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_146_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07103_ _07382_/A vssd1 vssd1 vccd1 vccd1 _07142_/B sky130_fd_sc_hd__clkbuf_2
X_08083_ _08095_/B vssd1 vssd1 vccd1 vccd1 _08083_/Y sky130_fd_sc_hd__inv_2
X_05295_ _05295_/A _05389_/A vssd1 vssd1 vccd1 vccd1 _05382_/B sky130_fd_sc_hd__nand2_1
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07034_ _07043_/A _07034_/B vssd1 vssd1 vccd1 vccd1 _07415_/C sky130_fd_sc_hd__xnor2_1
XFILLER_161_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08985_ _09168_/A vssd1 vssd1 vccd1 vccd1 _08985_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07936_ _07950_/A vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__buf_2
XFILLER_68_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07867_ _06204_/A _07849_/X _07850_/X _07866_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ _07867_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_44_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09606_ _09369_/X _09606_/B vssd1 vssd1 vccd1 vccd1 _09676_/D sky130_fd_sc_hd__and2b_1
X_06818_ _06818_/A _06818_/B vssd1 vssd1 vccd1 vccd1 _07767_/B sky130_fd_sc_hd__xnor2_4
XFILLER_28_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07798_ _07798_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _07802_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10848__D _10848_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09537_ _09538_/A _09638_/C vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06749_ _06769_/A _06758_/C vssd1 vssd1 vccd1 vccd1 _06772_/A sky130_fd_sc_hd__and2_1
XFILLER_71_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09468_ _09534_/C _09469_/B vssd1 vssd1 vccd1 vccd1 _09520_/A sky130_fd_sc_hd__or2_1
XFILLER_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08419_ _08419_/A _08419_/B vssd1 vssd1 vccd1 vccd1 _08419_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09399_ _09400_/B _09399_/B vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__and2b_1
XFILLER_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08787__A2 _08785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10312_ _10312_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10312_/X sky130_fd_sc_hd__xor2_1
XFILLER_164_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10243_ _10243_/A vssd1 vssd1 vccd1 vccd1 _10245_/A sky130_fd_sc_hd__inv_2
XFILLER_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10174_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10174_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input45_A io_wbs_m2s_data[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05990__A _08462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05289__A1 _05279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10282__A1 _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08525__B _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06061__A _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05982_ _05982_/A _05993_/S vssd1 vssd1 vccd1 vccd1 _05982_/Y sky130_fd_sc_hd__nor2_1
X_08770_ _10811_/Q vssd1 vssd1 vccd1 vccd1 _08771_/A sky130_fd_sc_hd__clkbuf_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07721_ _07721_/A vssd1 vssd1 vccd1 vccd1 _07721_/Y sky130_fd_sc_hd__inv_2
XFILLER_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07652_ _07653_/A _07653_/B vssd1 vssd1 vccd1 vccd1 _07654_/A sky130_fd_sc_hd__or2_1
XFILLER_92_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06603_ _06616_/A _06616_/B vssd1 vssd1 vccd1 vccd1 _06672_/A sky130_fd_sc_hd__xor2_1
XANTENNA__05405__A _05405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07583_ _07582_/B _07583_/B vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__and2b_1
XFILLER_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09322_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__nand2_1
X_06534_ _06535_/B _06534_/B vssd1 vssd1 vccd1 vccd1 _06536_/A sky130_fd_sc_hd__and2b_1
XFILLER_22_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09253_ _10822_/Q _09243_/X _09244_/X _09252_/X _09239_/X vssd1 vssd1 vccd1 vccd1
+ _09254_/B sky130_fd_sc_hd__a32o_1
X_06465_ _06465_/A _06465_/B vssd1 vssd1 vccd1 vccd1 _06466_/B sky130_fd_sc_hd__nor2_1
X_05416_ _10622_/Q _05389_/Y _05393_/X _05415_/X vssd1 vssd1 vccd1 vccd1 _05416_/X
+ sky130_fd_sc_hd__o22a_1
X_08204_ _08204_/A vssd1 vssd1 vccd1 vccd1 _10694_/D sky130_fd_sc_hd__clkbuf_1
X_09184_ _09202_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _10847_/D sky130_fd_sc_hd__nor2_4
X_06396_ _06396_/A vssd1 vssd1 vccd1 vccd1 _06871_/A sky130_fd_sc_hd__clkinv_2
XFILLER_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08135_ _08131_/X _08133_/X _08134_/X vssd1 vssd1 vccd1 vccd1 _10687_/D sky130_fd_sc_hd__o21a_1
X_05347_ _10669_/Q _05347_/B vssd1 vssd1 vccd1 vccd1 _05348_/B sky130_fd_sc_hd__nand2_1
XFILLER_135_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08066_ _08113_/A vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__buf_2
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05278_ _10651_/Q vssd1 vssd1 vccd1 vccd1 _05279_/A sky130_fd_sc_hd__buf_4
XANTENNA__05988__C1 _05977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ _07186_/A vssd1 vssd1 vccd1 vccd1 _07229_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_150_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08968_ _08968_/A vssd1 vssd1 vccd1 vccd1 _08968_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07919_ _07919_/A vssd1 vssd1 vccd1 vccd1 _07919_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08899_ input35/X _08785_/X _08786_/X hold12/A _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08899_/X sky130_fd_sc_hd__o221a_1
XFILLER_1_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10930_ _10930_/CLK _10930_/D vssd1 vssd1 vccd1 vccd1 _10930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05315__A _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10861_ _10862_/CLK _10861_/D vssd1 vssd1 vccd1 vccd1 _10861_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _10792_/CLK _10792_/D vssd1 vssd1 vccd1 vccd1 _10792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09221__S _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05985__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10226_ _10226_/A _10226_/B _10226_/C vssd1 vssd1 vccd1 vccd1 _10226_/X sky130_fd_sc_hd__and3_1
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10157_ _10157_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10088_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__or2_1
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08696__A1 _06147_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08536__A _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06250_ input37/X _06238_/X _06249_/X _06247_/X vssd1 vssd1 vccd1 vccd1 _10613_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_31_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06056__A _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06181_ _06178_/X _06158_/X _06180_/Y _06176_/X vssd1 vssd1 vccd1 vccd1 _10593_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09940_ _09940_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09941_/B sky130_fd_sc_hd__nand2_1
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10827__CLK _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _09933_/A _09871_/B vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__nand2_1
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08822_ _08814_/X _08817_/X _08818_/Y _08821_/X vssd1 vssd1 vccd1 vccd1 _10816_/D
+ sky130_fd_sc_hd__o31a_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08753_ _08759_/B _08753_/B vssd1 vssd1 vccd1 vccd1 _08753_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_73_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05965_ input8/X _09142_/C vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__or2_2
XANTENNA__10977__CLK _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08136__B1 _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07704_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _07704_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _10526_/A _08672_/X _08674_/X _10801_/Q vssd1 vssd1 vccd1 vccd1 _08684_/X
+ sky130_fd_sc_hd__a22o_1
X_05896_ _05896_/A vssd1 vssd1 vccd1 vccd1 _06035_/A sky130_fd_sc_hd__buf_2
XFILLER_93_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10494__A1 _06168_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07635_ _07635_/A _07635_/B vssd1 vssd1 vccd1 vccd1 _07636_/B sky130_fd_sc_hd__nand2_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09305_ _10898_/Q _10882_/Q vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__and2b_2
X_06517_ _06517_/A _06517_/B _06517_/C vssd1 vssd1 vccd1 vccd1 _06612_/A sky130_fd_sc_hd__and3_1
XFILLER_16_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07497_ _07497_/A _07497_/B vssd1 vssd1 vccd1 vccd1 _07534_/A sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_37_clock_A _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09236_ _09236_/A vssd1 vssd1 vccd1 vccd1 _10854_/D sky130_fd_sc_hd__buf_2
X_06448_ _06469_/B _06448_/B vssd1 vssd1 vccd1 vccd1 _06470_/A sky130_fd_sc_hd__and2b_1
XFILLER_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06379_ _06408_/B _06409_/C _06393_/A vssd1 vssd1 vccd1 vccd1 _06381_/C sky130_fd_sc_hd__a21oi_1
X_09167_ _09113_/X _09166_/X _08943_/X vssd1 vssd1 vccd1 vccd1 _09167_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08118_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__buf_2
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09098_ _09098_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__or2_1
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08049_ input8/X _09124_/C vssd1 vssd1 vccd1 vccd1 _08416_/A sky130_fd_sc_hd__nor2_1
XFILLER_135_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10011_ _10012_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10081_/B sky130_fd_sc_hd__and2_1
XFILLER_89_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08375__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10913_ _10980_/CLK _10913_/D vssd1 vssd1 vccd1 vccd1 _10913_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06015__D_N input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10844_ _10847_/CLK _10844_/D vssd1 vssd1 vccd1 vccd1 _10844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10775_ _10782_/CLK _10775_/D vssd1 vssd1 vccd1 vccd1 _10775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10209_ _10202_/X _10203_/X _10208_/X vssd1 vssd1 vccd1 vccd1 _10209_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07435__A _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05750_ _05744_/Y _10557_/Q _05747_/X _05749_/X vssd1 vssd1 vccd1 vccd1 _05750_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_76_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05681_ _10568_/Q _05681_/B vssd1 vssd1 vccd1 vccd1 _05684_/B sky130_fd_sc_hd__xnor2_1
XFILLER_62_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07420_ _07555_/B _07418_/Y _07419_/X vssd1 vssd1 vccd1 vccd1 _07426_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08266__A _08267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07351_ _07470_/B _07482_/A _07470_/A vssd1 vssd1 vccd1 vccd1 _07471_/A sky130_fd_sc_hd__o21a_1
XFILLER_149_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06302_ _06386_/A _06302_/B _06416_/A vssd1 vssd1 vccd1 vccd1 _06305_/C sky130_fd_sc_hd__or3b_1
X_07282_ _07282_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _07291_/B sky130_fd_sc_hd__or2_1
XFILLER_149_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06233_ _10607_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06233_/X sky130_fd_sc_hd__or2_1
X_09021_ _06066_/Y _06212_/B _08995_/X vssd1 vssd1 vccd1 vccd1 _09021_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_164_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06164_ _10590_/Q vssd1 vssd1 vccd1 vccd1 _06165_/A sky130_fd_sc_hd__inv_2
XFILLER_116_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10400__A1 _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06095_ _10683_/Q _10682_/Q _08075_/B vssd1 vssd1 vccd1 vccd1 _08098_/B sky130_fd_sc_hd__or3_2
XFILLER_116_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09923_ _09923_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09924_/B sky130_fd_sc_hd__or2_1
XFILLER_160_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09854_ _09795_/A _09795_/B _09853_/Y vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__a21bo_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _10814_/Q _10813_/Q _10812_/Q _08771_/A _08801_/B vssd1 vssd1 vccd1 vccd1
+ _08806_/B sky130_fd_sc_hd__o41a_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09785_ _09661_/X _09724_/A _09723_/Y vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__o21ai_1
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ _07013_/A _06997_/B _06997_/C vssd1 vssd1 vccd1 vccd1 _07007_/B sky130_fd_sc_hd__or3_1
XFILLER_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08736_ _08740_/C _08736_/B vssd1 vssd1 vccd1 vccd1 _08736_/X sky130_fd_sc_hd__xor2_1
X_05948_ _08350_/A _05829_/X _05946_/X _05947_/X vssd1 vssd1 vccd1 vccd1 _05948_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _10800_/Q _08678_/A vssd1 vssd1 vccd1 vccd1 _08669_/C sky130_fd_sc_hd__or2_1
XFILLER_82_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05879_ _10661_/Q vssd1 vssd1 vccd1 vccd1 _07988_/A sky130_fd_sc_hd__buf_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _07618_/A _07618_/B vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__xor2_4
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09609__B1 _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08598_ _10283_/A vssd1 vssd1 vccd1 vccd1 _08649_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05894__A1 _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ _07549_/A _07549_/B vssd1 vssd1 vccd1 vccd1 _07550_/B sky130_fd_sc_hd__and2_1
XANTENNA__09085__A1 _10937_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08832__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ _10562_/CLK _10560_/D vssd1 vssd1 vccd1 vccd1 _10560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09245_/S sky130_fd_sc_hd__clkbuf_2
X_10491_ _10491_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _10491_/X sky130_fd_sc_hd__or2_1
XFILLER_136_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07399__B2 _07560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08899__A1 input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10458__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08520__B1 _08517_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07702__B _07702_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05503__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10827_ _10856_/CLK _10827_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09076__B2 _08117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10758_ _10935_/CLK _10758_/D vssd1 vssd1 vccd1 vccd1 _10758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10689_ _10693_/CLK _10689_/D vssd1 vssd1 vccd1 vccd1 _10689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06053__B _08268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06920_ _06939_/A _06939_/B vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__nor2_2
XFILLER_68_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06851_ _06851_/A _06851_/B vssd1 vssd1 vccd1 vccd1 _06852_/B sky130_fd_sc_hd__nand2_1
XFILLER_68_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05802_ _05802_/A _05802_/B vssd1 vssd1 vccd1 vccd1 _05802_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09570_ _09570_/A _09574_/B vssd1 vssd1 vccd1 vccd1 _09570_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06782_ _06782_/A _06782_/B vssd1 vssd1 vccd1 vccd1 _06892_/B sky130_fd_sc_hd__nor2_2
X_08521_ _08935_/A input3/X vssd1 vssd1 vccd1 vccd1 _08522_/A sky130_fd_sc_hd__and2_1
XFILLER_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10449__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05733_ _08082_/A vssd1 vssd1 vccd1 vccd1 _05733_/X sky130_fd_sc_hd__buf_2
XFILLER_64_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08452_ _10772_/Q _10735_/Q _08455_/S vssd1 vssd1 vccd1 vccd1 _08453_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05664_ _05664_/A _05664_/B vssd1 vssd1 vccd1 vccd1 _05664_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07403_ _07404_/A _07404_/B vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__nor2_1
X_05595_ _10561_/Q _05602_/A _10562_/Q vssd1 vssd1 vccd1 vccd1 _05596_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09067__A1 _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08383_ _08419_/A vssd1 vssd1 vccd1 vccd1 _08383_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07334_ _07334_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07335_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07265_ _07269_/A _07514_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__a21oi_1
XFILLER_164_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09004_ _09867_/A vssd1 vssd1 vccd1 vccd1 _09931_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06216_ hold7/A _06223_/B vssd1 vssd1 vccd1 vccd1 _06216_/X sky130_fd_sc_hd__or2_1
XFILLER_164_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07196_ _07196_/A _07196_/B vssd1 vssd1 vccd1 vccd1 _07197_/C sky130_fd_sc_hd__xor2_1
XFILLER_145_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clock_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06147_ _10528_/A vssd1 vssd1 vccd1 vccd1 _06147_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06078_ _08251_/B _08244_/A vssd1 vssd1 vccd1 vccd1 _06078_/X sky130_fd_sc_hd__xor2_1
XFILLER_105_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09906_ _09906_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09837_ _09837_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09838_/B sky130_fd_sc_hd__or2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09768_ _09773_/A _09773_/B vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__nor2_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09290__A _09290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _08865_/B vssd1 vssd1 vccd1 vccd1 _08840_/B sky130_fd_sc_hd__buf_2
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _09769_/A _09764_/A _09810_/B _09769_/B vssd1 vssd1 vccd1 vccd1 _09844_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05867__A1 _08233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10612_ _10864_/CLK _10612_/D vssd1 vssd1 vccd1 vccd1 _10612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10543_ _10545_/CLK _10543_/D vssd1 vssd1 vccd1 vccd1 _10543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10474_ _10495_/A _10474_/B vssd1 vssd1 vccd1 vccd1 _10489_/B sky130_fd_sc_hd__nand2_2
XFILLER_124_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08033__A2 _07985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06044__B2 _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_6_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07713__A _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_92_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05380_ _05380_/A _05380_/B vssd1 vssd1 vccd1 vccd1 _05380_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07050_ _07048_/A _07048_/B _07464_/A vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__a21oi_1
XFILLER_146_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06001_ _10528_/A _07849_/A _06120_/S vssd1 vssd1 vccd1 vccd1 _06002_/B sky130_fd_sc_hd__mux2_1
XFILLER_161_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07952_ _07955_/A _07952_/B vssd1 vssd1 vccd1 vccd1 _07953_/A sky130_fd_sc_hd__or2_1
XFILLER_87_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06903_ _06903_/A _06903_/B vssd1 vssd1 vccd1 vccd1 _06921_/B sky130_fd_sc_hd__xor2_2
XFILLER_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07883_ hold5/X _07870_/X _07874_/X _07882_/Y vssd1 vssd1 vccd1 vccd1 _07884_/B sky130_fd_sc_hd__o2bb2a_1
X_09622_ _09623_/A _09623_/B _09623_/C vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__o21ai_1
XFILLER_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06834_ _06834_/A _06834_/B vssd1 vssd1 vccd1 vccd1 _06835_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09553_ _09553_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09554_/C sky130_fd_sc_hd__xnor2_1
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06765_ _06834_/A _06765_/B vssd1 vssd1 vccd1 vccd1 _06766_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08504_ _10787_/Q _08496_/X _08502_/X _10750_/Q vssd1 vssd1 vccd1 vccd1 _10750_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05716_ _08196_/A _10555_/Q _05663_/A _05704_/Y vssd1 vssd1 vccd1 vccd1 _05717_/D
+ sky130_fd_sc_hd__a22o_1
X_09484_ _10967_/Q _09579_/A vssd1 vssd1 vccd1 vccd1 _09486_/A sky130_fd_sc_hd__and2_1
XANTENNA__06239__A _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06696_ _06693_/A _06693_/B _06691_/A vssd1 vssd1 vccd1 vccd1 _06697_/B sky130_fd_sc_hd__o21a_1
XFILLER_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08435_ _10767_/Q _10730_/Q _08486_/S vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__mux2_1
XFILLER_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05647_ _05912_/B _05539_/Y _05540_/X _05646_/X vssd1 vssd1 vccd1 vccd1 _05647_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08366_ _08531_/A vssd1 vssd1 vccd1 vccd1 _08419_/A sky130_fd_sc_hd__clkbuf_2
X_05578_ _08315_/B vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08799__B1 _08786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07317_ _07317_/A _07317_/B vssd1 vssd1 vccd1 vccd1 _07341_/A sky130_fd_sc_hd__or2_1
XFILLER_109_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08297_/Y sky130_fd_sc_hd__nand2_1
XFILLER_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07248_ _07248_/A _07382_/A vssd1 vssd1 vccd1 vccd1 _07517_/A sky130_fd_sc_hd__and2_1
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07179_ _07188_/B vssd1 vssd1 vccd1 vccd1 _07587_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__A _09285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ _10947_/Q _10931_/Q vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__or2b_1
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08420__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_30_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10942_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_43_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_45_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10728_/CLK sky130_fd_sc_hd__clkbuf_16
Xinput16 io_wbs_m2s_data[0] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_6
XANTENNA_clkbuf_leaf_85_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput27 io_wbs_m2s_data[1] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_6
XFILLER_7_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 io_wbs_m2s_data[2] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_4
Xinput49 io_wbs_m2s_stb vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_6
X_10526_ _10526_/A _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10526_/X sky130_fd_sc_hd__or3_1
XFILLER_116_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10457_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10457_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07708__A _07708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ _10365_/X _10716_/Q _10386_/X _10387_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10935_/D sky130_fd_sc_hd__o221a_1
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07765__A1 _10504_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06550_ _10971_/Q _06550_/B _06550_/C vssd1 vssd1 vccd1 vccd1 _06587_/B sky130_fd_sc_hd__and3_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05501_ _05369_/Y _05497_/X _05495_/X _05460_/C vssd1 vssd1 vccd1 vccd1 _10554_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_21_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06481_ _06480_/B _06480_/C _06480_/A vssd1 vssd1 vccd1 vccd1 _06657_/A sky130_fd_sc_hd__o21a_1
X_08220_ _08216_/X _08224_/C _08067_/X vssd1 vssd1 vccd1 vccd1 _08220_/Y sky130_fd_sc_hd__o21ai_1
X_05432_ _10637_/Q vssd1 vssd1 vccd1 vccd1 _07893_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08274__A input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _08160_/B _08151_/B vssd1 vssd1 vccd1 vccd1 _08151_/Y sky130_fd_sc_hd__nand2_1
X_05363_ _05363_/A _05363_/B vssd1 vssd1 vccd1 vccd1 _05363_/X sky130_fd_sc_hd__and2_1
XANTENNA__08245__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07102_ _07102_/A vssd1 vssd1 vccd1 vccd1 _07382_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05294_ _05388_/A _05392_/A vssd1 vssd1 vccd1 vccd1 _05389_/A sky130_fd_sc_hd__and2_1
X_08082_ _08082_/A _08082_/B _08082_/C _08082_/D vssd1 vssd1 vccd1 vccd1 _08095_/B
+ sky130_fd_sc_hd__and4_1
X_07033_ _07044_/A _07421_/A _07417_/A vssd1 vssd1 vccd1 vccd1 _07034_/B sky130_fd_sc_hd__and3_1
XFILLER_134_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08984_ _09035_/B vssd1 vssd1 vccd1 vccd1 _09168_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_102_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07935_ _10432_/B _07935_/B vssd1 vssd1 vccd1 vccd1 _07950_/A sky130_fd_sc_hd__nand2_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05519__B1 _05474_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07866_ _10880_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07866_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09605_ _09549_/A _09549_/B _09678_/A vssd1 vssd1 vccd1 vccd1 _09608_/A sky130_fd_sc_hd__o21ai_2
X_06817_ _07670_/A _06817_/B vssd1 vssd1 vccd1 vccd1 _06818_/B sky130_fd_sc_hd__nand2_2
XFILLER_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07797_ _07797_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__xnor2_1
XFILLER_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09536_ _10969_/Q _09536_/B vssd1 vssd1 vccd1 vccd1 _09638_/C sky130_fd_sc_hd__nand2_1
XFILLER_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06748_ _06758_/B _06774_/B vssd1 vssd1 vccd1 vccd1 _06748_/X sky130_fd_sc_hd__and2_1
XFILLER_25_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09467_ _09516_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__or2_1
X_06679_ _06678_/A _06678_/C _06678_/B vssd1 vssd1 vccd1 vccd1 _06945_/B sky130_fd_sc_hd__a21oi_1
XFILLER_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08418_ _10394_/B _08418_/B vssd1 vssd1 vccd1 vccd1 _08419_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09398_ _09433_/A _09398_/B vssd1 vssd1 vccd1 vccd1 _09399_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ _08351_/A _08350_/B vssd1 vssd1 vccd1 vccd1 _08349_/X sky130_fd_sc_hd__and2_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10311_ _10310_/X _10309_/A _10329_/S vssd1 vssd1 vccd1 vccd1 _10312_/B sky130_fd_sc_hd__mux2_1
XFILLER_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10242_ _10937_/Q _10953_/Q vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__or2b_1
XFILLER_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10173_ _07056_/A _10167_/X _10170_/X _10886_/Q vssd1 vssd1 vccd1 vccd1 _10886_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_121_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input38_A io_wbs_m2s_data[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_5_0_clock _10856_/CLK vssd1 vssd1 vccd1 vccd1 _10836_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08094__A _08098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07986__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10509_ _05958_/X _10496_/X _10508_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10975_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_171_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07438__A _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06061__B _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05981_ _10533_/A vssd1 vssd1 vccd1 vccd1 _05982_/A sky130_fd_sc_hd__clkbuf_4
X_07720_ _07720_/A _07720_/B vssd1 vssd1 vccd1 vccd1 _07745_/A sky130_fd_sc_hd__xnor2_1
XFILLER_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07651_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _07653_/B sky130_fd_sc_hd__xnor2_1
XFILLER_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06602_ _06602_/A _06602_/B vssd1 vssd1 vccd1 vccd1 _06616_/B sky130_fd_sc_hd__or2_1
X_07582_ _07583_/B _07582_/B vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__and2b_1
XFILLER_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09321_ _09396_/B _09396_/C vssd1 vssd1 vccd1 vccd1 _09323_/B sky130_fd_sc_hd__xor2_1
X_06533_ _06533_/A _06538_/B vssd1 vssd1 vccd1 vccd1 _06534_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09252_ _08289_/A _09251_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09252_/X sky130_fd_sc_hd__mux2_1
X_06464_ _06465_/A _06465_/B vssd1 vssd1 vccd1 vccd1 _06480_/C sky130_fd_sc_hd__and2_1
XFILLER_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ _08200_/X _08203_/B vssd1 vssd1 vccd1 vccd1 _08204_/A sky130_fd_sc_hd__and2b_1
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05415_ _05462_/C _05393_/B _05414_/X vssd1 vssd1 vccd1 vccd1 _05415_/X sky130_fd_sc_hd__o21a_1
XFILLER_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09183_ _09112_/A _09178_/Y _09182_/X vssd1 vssd1 vccd1 vccd1 _09184_/B sky130_fd_sc_hd__a21oi_1
X_06395_ _06874_/A _06395_/B vssd1 vssd1 vccd1 vccd1 _06396_/A sky130_fd_sc_hd__xnor2_1
X_08134_ _06168_/X _08047_/X _08052_/X _08132_/A _08054_/X vssd1 vssd1 vccd1 vccd1
+ _08134_/X sky130_fd_sc_hd__o221a_1
X_05346_ _05347_/B _05346_/B vssd1 vssd1 vccd1 vccd1 _05346_/X sky130_fd_sc_hd__and2_1
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08732__A _10806_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08065_ _10580_/Q _08065_/B vssd1 vssd1 vccd1 vccd1 _08113_/A sky130_fd_sc_hd__and2_2
XFILLER_161_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05277_ _05291_/A _05818_/B vssd1 vssd1 vccd1 vccd1 _05277_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07016_ _07235_/C vssd1 vssd1 vccd1 vccd1 _07186_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08967_ _08962_/Y _10495_/B _08966_/Y vssd1 vssd1 vccd1 vccd1 _08967_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_33_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07918_ _09154_/A vssd1 vssd1 vccd1 vccd1 _08284_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_112_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08898_ _08889_/A _08892_/Y _08896_/X _08688_/A vssd1 vssd1 vccd1 vccd1 _08898_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10502__A _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08154__A1 input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08154__B2 _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07849_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07849_/X sky130_fd_sc_hd__buf_4
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10860_ _10860_/CLK _10860_/D vssd1 vssd1 vccd1 vccd1 _10860_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09519_ _09562_/B _09562_/C _09562_/A vssd1 vssd1 vccd1 vccd1 _09520_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__07811__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _10792_/CLK _10791_/D vssd1 vssd1 vccd1 vccd1 _10791_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08626__B _08649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05985__B input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06162__A input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10225_ _10225_/A _10225_/B vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__nor2_1
XFILLER_106_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10156_ _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _10157_/B sky130_fd_sc_hd__xnor2_1
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10087_ _10087_/A _10087_/B vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10412__A _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05506__A _05513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09920__B _09920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06180_ _06180_/A _06193_/B vssd1 vssd1 vccd1 vccd1 _06180_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08081__B1 _05733_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10204__B_N _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _09870_/A _09870_/B _09870_/C vssd1 vssd1 vccd1 vccd1 _09871_/B sky130_fd_sc_hd__or3_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09377__B_N _06993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08821_ input24/X _08819_/X _08820_/X _10816_/Q _08310_/X vssd1 vssd1 vccd1 vccd1
+ _08821_/X sky130_fd_sc_hd__o221a_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08748_/X _08815_/B _08759_/A vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__a21oi_1
X_05964_ input7/X input4/X input9/X vssd1 vssd1 vccd1 vccd1 _09142_/C sky130_fd_sc_hd__or3_2
X_07703_ _09824_/A _09824_/B _07702_/X vssd1 vssd1 vccd1 vccd1 _09899_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08683_ _08778_/A _08683_/B _08692_/B vssd1 vssd1 vccd1 vccd1 _08683_/X sky130_fd_sc_hd__and3_1
X_05895_ _05895_/A _05895_/B vssd1 vssd1 vccd1 vccd1 _05895_/X sky130_fd_sc_hd__and2_1
XFILLER_26_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07634_ _07670_/A vssd1 vssd1 vccd1 vccd1 _07635_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07565_ _07563_/X _07565_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__and2b_1
XFILLER_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09304_ _09304_/A _10882_/Q vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06516_ _06517_/A _06517_/B _06680_/A vssd1 vssd1 vccd1 vccd1 _06521_/B sky130_fd_sc_hd__and3_1
X_07496_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07534_/C sky130_fd_sc_hd__nor2_1
XFILLER_10_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09235_ _09259_/A _09235_/B vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__and2_2
X_06447_ _06472_/A _06472_/B _06675_/A _06675_/B vssd1 vssd1 vccd1 vccd1 _06448_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_10_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _09114_/X _09165_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__o21a_1
X_06378_ _06872_/A _06409_/C vssd1 vssd1 vccd1 vccd1 _06393_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08462__A _08462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08117_ _08117_/A _08117_/B vssd1 vssd1 vccd1 vccd1 _08117_/Y sky130_fd_sc_hd__nand2_1
X_05329_ _05329_/A _05329_/B vssd1 vssd1 vccd1 vccd1 _05329_/X sky130_fd_sc_hd__and2_1
XFILLER_135_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09097_ _10129_/A vssd1 vssd1 vccd1 vccd1 _10493_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08048_ _08048_/A vssd1 vssd1 vccd1 vccd1 _09124_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_150_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10010_ _10081_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10182__A1 _07008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _09999_/A vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__inv_2
XFILLER_62_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05326__A _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10912_ _10925_/CLK _10912_/D vssd1 vssd1 vccd1 vccd1 _10912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10843_ _10987_/CLK _10843_/D vssd1 vssd1 vccd1 vccd1 _10843_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10774_ _10776_/CLK _10774_/D vssd1 vssd1 vccd1 vccd1 _10774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05996__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08063__B1 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10208_ _10226_/A _10206_/Y _10279_/S vssd1 vssd1 vccd1 vccd1 _10208_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07435__B _07713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10139_ _10138_/B _10138_/Y _10139_/S vssd1 vssd1 vccd1 vccd1 _10143_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09866__B2 _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05680_ _05803_/A vssd1 vssd1 vccd1 vccd1 _08317_/A sky130_fd_sc_hd__buf_2
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07350_ _07461_/B _07350_/B vssd1 vssd1 vccd1 vccd1 _07470_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06301_ _10921_/Q _10904_/Q vssd1 vssd1 vccd1 vccd1 _06386_/A sky130_fd_sc_hd__xnor2_4
X_07281_ _07282_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _07366_/B sky130_fd_sc_hd__nand2_1
X_09020_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _09020_/X sky130_fd_sc_hd__or2_1
X_06232_ input30/X _06225_/X _06231_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10606_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06163_ _10535_/A vssd1 vssd1 vccd1 vccd1 _06163_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_129_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06094_ _10681_/Q _10680_/Q vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__or2_2
XFILLER_171_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09922_ _10065_/D _09922_/B vssd1 vssd1 vccd1 vccd1 _09925_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__06080__A2 _07998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09853_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09853_/Y sky130_fd_sc_hd__nand2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08804_ _08804_/A _08804_/B _08804_/C _08804_/D vssd1 vssd1 vccd1 vccd1 _08804_/Y
+ sky130_fd_sc_hd__nand4_1
X_09784_ _09784_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__or2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _10907_/Q vssd1 vssd1 vccd1 vccd1 _07013_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _10805_/Q _08815_/B _08726_/Y vssd1 vssd1 vccd1 vccd1 _08736_/B sky130_fd_sc_hd__a21bo_1
X_05947_ _08339_/A _05947_/B vssd1 vssd1 vccd1 vccd1 _05947_/X sky130_fd_sc_hd__or2_1
XFILLER_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__B1 _07865_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _10800_/Q _08678_/A vssd1 vssd1 vccd1 vccd1 _08669_/B sky130_fd_sc_hd__nand2_1
X_05878_ _07991_/A _05878_/B vssd1 vssd1 vccd1 vccd1 _05878_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07617_ _07622_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07618_/A sky130_fd_sc_hd__nand2_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ _08661_/A _08597_/B vssd1 vssd1 vccd1 vccd1 _08617_/B sky130_fd_sc_hd__and2_1
XFILLER_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07548_ _07549_/A _07549_/B vssd1 vssd1 vccd1 vccd1 _07743_/B sky130_fd_sc_hd__nor2_1
XFILLER_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07479_ _07497_/A _07497_/B vssd1 vssd1 vccd1 vccd1 _07504_/B sky130_fd_sc_hd__and2_1
XFILLER_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09218_ _09218_/A vssd1 vssd1 vccd1 vccd1 _10851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _05982_/A _10489_/B _10489_/Y _10485_/X vssd1 vssd1 vccd1 vccd1 _10968_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08045__B1 _06033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ _05461_/B _09136_/X _09148_/X _08160_/A _07935_/B vssd1 vssd1 vccd1 vccd1
+ _09149_/X sky130_fd_sc_hd__a221o_1
XFILLER_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_2_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08899__A2 _08785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input20_A io_wbs_m2s_data[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10826_ _10830_/CLK _10826_/D vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_158_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_2_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10757_ _10792_/CLK _10757_/D vssd1 vssd1 vccd1 vccd1 _10757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10688_ _10693_/CLK _10688_/D vssd1 vssd1 vccd1 vccd1 _10688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06062__A2 _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06850_ _06850_/A _06288_/X vssd1 vssd1 vccd1 vccd1 _06852_/A sky130_fd_sc_hd__or2b_1
X_05801_ _05717_/X _05742_/C _05796_/X _05800_/X _05702_/X vssd1 vssd1 vccd1 vccd1
+ _05802_/B sky130_fd_sc_hd__o32a_1
X_06781_ _06781_/A _06781_/B vssd1 vssd1 vccd1 vccd1 _06782_/B sky130_fd_sc_hd__nor2_1
XFILLER_110_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08520_ _10798_/Q _08514_/X _08517_/X _10761_/Q vssd1 vssd1 vccd1 vccd1 _10761_/D
+ sky130_fd_sc_hd__a22o_1
X_05732_ _05794_/A _05732_/B _05732_/C _05732_/D vssd1 vssd1 vccd1 vccd1 _05788_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_36_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08451_ _08451_/A vssd1 vssd1 vccd1 vccd1 _10734_/D sky130_fd_sc_hd__clkbuf_1
X_05663_ _05663_/A _05663_/B vssd1 vssd1 vccd1 vccd1 _05664_/B sky130_fd_sc_hd__and2_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07402_ _07402_/A _07402_/B vssd1 vssd1 vccd1 vccd1 _07404_/B sky130_fd_sc_hd__xnor2_1
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08382_ _08367_/X _10734_/Q _08380_/X _08381_/X vssd1 vssd1 vccd1 vccd1 _10716_/D
+ sky130_fd_sc_hd__o211a_1
X_05594_ _10701_/Q vssd1 vssd1 vccd1 vccd1 _08277_/B sky130_fd_sc_hd__clkbuf_2
X_07333_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07522_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07264_ _07264_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07266_/A sky130_fd_sc_hd__xor2_1
XFILLER_137_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09003_ _09610_/A vssd1 vssd1 vccd1 vccd1 _09867_/A sky130_fd_sc_hd__clkbuf_2
X_06215_ _06206_/X _06207_/X _06214_/X _06200_/X vssd1 vssd1 vccd1 vccd1 _10599_/D
+ sky130_fd_sc_hd__o211a_1
X_07195_ _07195_/A _07334_/A vssd1 vssd1 vccd1 vccd1 _07196_/B sky130_fd_sc_hd__or2b_1
XFILLER_3_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06146_ _06143_/X _06131_/X _06145_/Y _06137_/X vssd1 vssd1 vccd1 vccd1 _10586_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06077_ _08355_/A _08352_/A _08029_/A _10709_/Q _06076_/X vssd1 vssd1 vccd1 vccd1
+ _06082_/B sky130_fd_sc_hd__a221o_1
XFILLER_160_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07356__A _07560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _09971_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__nor2_1
XFILLER_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _09837_/A _09837_/B vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09767_ _09767_/A _09767_/B vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__and2_1
X_06979_ _10900_/Q vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _08856_/B vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _09767_/A _09767_/B vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10510__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _08649_/A _08649_/B _08649_/C vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__and3_1
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _10643_/CLK _10611_/D vssd1 vssd1 vccd1 vccd1 _10611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10542_ _10545_/CLK _10542_/D vssd1 vssd1 vccd1 vccd1 _10542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ _06206_/X _10459_/A _10472_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10962_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08741__A1 _10806_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06201__C1 _06200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10809_ _10942_/CLK _10809_/D vssd1 vssd1 vccd1 vccd1 _10809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06000_ _10577_/Q vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_161_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09375__B _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08980__A1 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07951_ input42/X _05905_/A _07983_/A vssd1 vssd1 vccd1 vccd1 _07952_/B sky130_fd_sc_hd__mux2_1
XFILLER_96_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06902_ _06902_/A _06902_/B vssd1 vssd1 vccd1 vccd1 _06921_/A sky130_fd_sc_hd__nor2_1
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07882_ _07882_/A vssd1 vssd1 vccd1 vccd1 _07882_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08193__C1 _08175_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _09621_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09623_/C sky130_fd_sc_hd__xor2_1
X_06833_ _06833_/A _06833_/B vssd1 vssd1 vccd1 vccd1 _06835_/A sky130_fd_sc_hd__nand2_1
X_09552_ _09610_/A _09552_/B _09599_/B vssd1 vssd1 vccd1 vccd1 _09604_/B sky130_fd_sc_hd__and3_1
X_06764_ _06834_/A _06765_/B vssd1 vssd1 vccd1 vccd1 _06766_/A sky130_fd_sc_hd__and2_1
XFILLER_55_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08503_ _10786_/Q _08496_/X _08502_/X _10749_/Q vssd1 vssd1 vccd1 vccd1 _10749_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05715_ _08139_/A _10549_/Q _05702_/X _05708_/Y _05714_/X vssd1 vssd1 vccd1 vccd1
+ _05717_/C sky130_fd_sc_hd__a2111o_1
XFILLER_36_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09483_ _09483_/A _09483_/B vssd1 vssd1 vccd1 vccd1 _09527_/A sky130_fd_sc_hd__xor2_4
XFILLER_70_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06695_ _06695_/A _06695_/B vssd1 vssd1 vccd1 vccd1 _06698_/B sky130_fd_sc_hd__xor2_2
XFILLER_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08434_ _08476_/S vssd1 vssd1 vccd1 vccd1 _08486_/S sky130_fd_sc_hd__buf_2
XFILLER_169_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05646_ _10681_/Q _05644_/Y _05541_/X vssd1 vssd1 vccd1 vccd1 _05646_/X sky130_fd_sc_hd__a21bo_1
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08365_ _10729_/Q vssd1 vssd1 vccd1 vccd1 _08531_/A sky130_fd_sc_hd__inv_2
X_05577_ _10705_/Q vssd1 vssd1 vccd1 vccd1 _08315_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08799__A1 _06206_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _07309_/A _07152_/B _07322_/A vssd1 vssd1 vccd1 vccd1 _07317_/B sky130_fd_sc_hd__a21oi_1
XFILLER_164_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08296_ _08297_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08296_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06255__A _07848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07247_ _07269_/A _07247_/B vssd1 vssd1 vccd1 vccd1 _07513_/A sky130_fd_sc_hd__nand2_1
XFILLER_164_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07178_ _07178_/A vssd1 vssd1 vccd1 vccd1 _07398_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06129_ _10432_/B _06129_/B vssd1 vssd1 vccd1 vccd1 _06149_/A sky130_fd_sc_hd__nand2_1
XFILLER_106_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10224__B _10935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09819_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09820_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10530__A1 _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08239__B1 _08124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_opt_1_0_clock clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _10835_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_28_clock_A _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput17 io_wbs_m2s_data[10] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_6
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 io_wbs_m2s_data[20] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_6
XFILLER_10_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 io_wbs_m2s_data[30] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_4
XFILLER_156_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ _07442_/X _10522_/X _10524_/X _10511_/X vssd1 vssd1 vccd1 vccd1 _10980_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10456_ _10956_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10456_/X sky130_fd_sc_hd__or2_1
XFILLER_136_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10349__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08380__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08411__B1 _08992_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _10935_/Q _10379_/B _10376_/X vssd1 vssd1 vccd1 vccd1 _10387_/X sky130_fd_sc_hd__a21bo_1
XFILLER_112_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05776__A1 _08297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05776__B2 _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05500_ _05371_/Y _05497_/X _05495_/X _05460_/D vssd1 vssd1 vccd1 vccd1 _10553_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_06480_ _06480_/A _06480_/B _06480_/C vssd1 vssd1 vccd1 vccd1 _06657_/B sky130_fd_sc_hd__nor3_1
XFILLER_33_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05431_ _07889_/A _05346_/X _05348_/X _10637_/Q _05430_/X vssd1 vssd1 vccd1 vccd1
+ _05431_/X sky130_fd_sc_hd__a221o_1
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__nand2_1
X_05362_ _10663_/Q _05362_/B vssd1 vssd1 vccd1 vccd1 _05363_/B sky130_fd_sc_hd__nand2_1
XFILLER_146_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07101_ _10986_/Q _07327_/A vssd1 vssd1 vccd1 vccd1 _07384_/A sky130_fd_sc_hd__nand2_1
X_08081_ _08075_/A _08059_/A _08082_/D _05733_/X vssd1 vssd1 vccd1 vccd1 _08081_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_146_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05293_ _10653_/Q _05391_/B vssd1 vssd1 vccd1 vccd1 _05392_/A sky130_fd_sc_hd__nor2_1
XFILLER_134_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07032_ _07042_/A _07042_/B vssd1 vssd1 vccd1 vccd1 _07043_/A sky130_fd_sc_hd__and2_1
XFILLER_106_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10325__A _10944_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08953__A1 _10931_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ _06019_/A _08972_/X _08974_/X _08982_/X vssd1 vssd1 vccd1 vccd1 _08983_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07934_ _08995_/A vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07634__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07865_ _08557_/A vssd1 vssd1 vccd1 vccd1 _07865_/X sky130_fd_sc_hd__buf_2
XANTENNA__09552__C _09599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10512__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08159__B1_N _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _09655_/A _09604_/B vssd1 vssd1 vccd1 vccd1 _09613_/B sky130_fd_sc_hd__and2_1
XANTENNA__10060__A _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06816_ _06856_/A vssd1 vssd1 vccd1 vccd1 _10502_/A sky130_fd_sc_hd__buf_2
X_07796_ _07796_/A _07796_/B _07795_/X vssd1 vssd1 vccd1 vccd1 _07797_/B sky130_fd_sc_hd__or3b_1
XFILLER_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09535_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__xnor2_1
X_06747_ _06785_/A _06747_/B _06776_/A vssd1 vssd1 vccd1 vccd1 _06763_/A sky130_fd_sc_hd__and3_1
XFILLER_25_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09466_ _09552_/B _09466_/B vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__and2_1
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06678_ _06678_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__and3_1
XFILLER_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05629_ _10548_/Q _05629_/B vssd1 vssd1 vccd1 vccd1 _05630_/B sky130_fd_sc_hd__nand2_1
X_08417_ _09037_/A vssd1 vssd1 vccd1 vccd1 _08418_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09397_ _10131_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09398_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08348_ input39/X vssd1 vssd1 vccd1 vccd1 _08348_/Y sky130_fd_sc_hd__inv_2
XFILLER_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08279_ _08278_/A _08278_/B _08255_/A vssd1 vssd1 vccd1 vccd1 _08279_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08912__B _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10310_ _10292_/A _10289_/A _10298_/B _10309_/Y vssd1 vssd1 vccd1 vccd1 _10310_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_137_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10241_ _07066_/A _10192_/X _10240_/Y vssd1 vssd1 vccd1 vccd1 _10903_/D sky130_fd_sc_hd__a21o_1
XFILLER_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10172_ _07113_/A _10167_/X _10170_/X _10885_/Q vssd1 vssd1 vccd1 vccd1 _10885_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10503__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05999__A input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10508_ _10508_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10508_/X sky130_fd_sc_hd__or2_1
XFILLER_7_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10439_ _10949_/Q _10431_/X _10438_/X vssd1 vssd1 vccd1 vccd1 _10949_/D sky130_fd_sc_hd__a21o_1
XFILLER_152_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05980_ input43/X vssd1 vssd1 vccd1 vccd1 _10533_/A sky130_fd_sc_hd__buf_6
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09186__A1_N _10945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07650_ _07659_/A _07658_/B _07635_/A vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__o21a_1
XFILLER_26_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06601_ _06775_/A _06409_/B _06522_/C vssd1 vssd1 vccd1 vccd1 _06602_/B sky130_fd_sc_hd__a21oi_1
XFILLER_81_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07581_ _07581_/A _07581_/B vssd1 vssd1 vccd1 vccd1 _07582_/B sky130_fd_sc_hd__xor2_1
XFILLER_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09320_ _10069_/A _09744_/A vssd1 vssd1 vccd1 vccd1 _09396_/C sky130_fd_sc_hd__nand2_1
X_06532_ _06532_/A _06532_/B vssd1 vssd1 vccd1 vccd1 _06538_/B sky130_fd_sc_hd__xor2_1
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09251_ _08287_/A _07900_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09251_/X sky130_fd_sc_hd__mux2_1
X_06463_ _06479_/A _06479_/B vssd1 vssd1 vccd1 vccd1 _06465_/B sky130_fd_sc_hd__xor2_1
X_08202_ input21/X _08123_/X _08124_/X _05877_/X _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08203_/B sky130_fd_sc_hd__o221a_1
XFILLER_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05414_ _10620_/Q _05487_/A _05413_/X vssd1 vssd1 vccd1 vccd1 _05414_/X sky130_fd_sc_hd__a21o_1
X_09182_ _10812_/Q _09168_/X _09079_/X _10725_/Q _09181_/X vssd1 vssd1 vccd1 vccd1
+ _09182_/X sky130_fd_sc_hd__a221o_1
X_06394_ _06394_/A _06394_/B vssd1 vssd1 vccd1 vccd1 _06395_/B sky130_fd_sc_hd__xnor2_1
X_08133_ _08038_/X _08074_/X _08132_/Y _08044_/X _06050_/X vssd1 vssd1 vccd1 vccd1
+ _08133_/X sky130_fd_sc_hd__a32o_1
X_05345_ _10667_/Q _05350_/B _10668_/Q vssd1 vssd1 vccd1 vccd1 _05346_/B sky130_fd_sc_hd__o21ai_1
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08064_ _05813_/A _08058_/X _08063_/X vssd1 vssd1 vccd1 vccd1 _08064_/X sky130_fd_sc_hd__o21ba_1
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05276_ _10576_/Q vssd1 vssd1 vccd1 vccd1 _05818_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05988__A1 _09078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07015_ _10982_/Q vssd1 vssd1 vccd1 vccd1 _07235_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_115_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08966_ _07780_/C _08964_/A _08965_/Y vssd1 vssd1 vccd1 vccd1 _08966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07917_ _08462_/A vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_44_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10855_/CLK sky130_fd_sc_hd__clkbuf_16
X_08897_ _08889_/A _08892_/Y _08896_/X vssd1 vssd1 vccd1 vccd1 _08897_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07848_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07848_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_84_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07779_ _07779_/A _07779_/B vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09518_ _09562_/A _09562_/B _09562_/C vssd1 vssd1 vccd1 vccd1 _09520_/B sky130_fd_sc_hd__and3_1
XFILLER_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _10790_/CLK _10790_/D vssd1 vssd1 vccd1 vccd1 _10790_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_59_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10665_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08311__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09449_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09552_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05979__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input50_A io_wbs_m2s_we vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09754__A _09754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _10224_/A _10935_/Q vssd1 vssd1 vccd1 vccd1 _10225_/B sky130_fd_sc_hd__and2_1
XFILLER_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10156_/B sky130_fd_sc_hd__xnor2_1
XFILLER_121_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10086_ _09998_/A _10138_/B _09997_/B _10017_/A vssd1 vssd1 vccd1 vccd1 _10087_/B
+ sky130_fd_sc_hd__a31oi_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08853__B1 _08786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08908__A1 input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08820_ _08820_/A vssd1 vssd1 vccd1 vccd1 _08820_/X sky130_fd_sc_hd__clkbuf_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05963_ _07967_/A vssd1 vssd1 vccd1 vccd1 _09016_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_08751_ _10808_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08759_/B sky130_fd_sc_hd__xor2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10322__B _10945_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07702_ _07621_/A _07702_/B vssd1 vssd1 vccd1 vccd1 _07702_/X sky130_fd_sc_hd__and2b_1
XFILLER_65_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05894_ _07974_/A _05900_/A _06039_/A vssd1 vssd1 vccd1 vccd1 _05895_/B sky130_fd_sc_hd__o21ai_1
X_08682_ _08669_/B _08670_/C _08679_/X _08680_/Y vssd1 vssd1 vccd1 vccd1 _08692_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07633_ _07633_/A _07633_/B vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__xor2_2
XFILLER_26_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07564_ _07563_/A _07727_/B _07563_/C vssd1 vssd1 vccd1 vccd1 _07565_/B sky130_fd_sc_hd__a21o_1
XFILLER_94_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09303_ _09303_/A _09303_/B vssd1 vssd1 vccd1 vccd1 _09310_/C sky130_fd_sc_hd__nor2_2
X_06515_ _06758_/B _06515_/B vssd1 vssd1 vccd1 vccd1 _06680_/A sky130_fd_sc_hd__nand2_1
X_07495_ _07495_/A _07495_/B vssd1 vssd1 vccd1 vccd1 _07506_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09234_ _08847_/X _09210_/X _09212_/X _09233_/X _09203_/X vssd1 vssd1 vccd1 vccd1
+ _09235_/B sky130_fd_sc_hd__a32o_1
XFILLER_10_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06446_ _06461_/B _06459_/B vssd1 vssd1 vccd1 vccd1 _06675_/B sky130_fd_sc_hd__nand2_1
XFILLER_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09165_ _10943_/Q _09008_/X _09164_/Y _08948_/X vssd1 vssd1 vccd1 vccd1 _09165_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06377_ _06436_/A _06513_/D vssd1 vssd1 vccd1 vccd1 _06409_/C sky130_fd_sc_hd__and2_1
X_08116_ _08117_/A _08116_/B vssd1 vssd1 vccd1 vccd1 _08116_/Y sky130_fd_sc_hd__nor2_1
X_05328_ _10675_/Q _05834_/A vssd1 vssd1 vccd1 vccd1 _05329_/B sky130_fd_sc_hd__nand2_1
X_09096_ _09977_/A vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06083__B1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08047_ _08248_/A vssd1 vssd1 vccd1 vccd1 _08047_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10513__A _10513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _09998_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09999_/A sky130_fd_sc_hd__xnor2_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08949_ input10/X vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__inv_2
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10911_ _10925_/CLK _10911_/D vssd1 vssd1 vccd1 vccd1 _10911_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09088__A0 _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _10847_/CLK _10842_/D vssd1 vssd1 vccd1 vccd1 _10842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10773_ _10782_/CLK _10773_/D vssd1 vssd1 vccd1 vccd1 _10773_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06074__B1 _07979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09484__A _10967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09012__A0 _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10207_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10279_/S sky130_fd_sc_hd__buf_2
XFILLER_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05517__A _05517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _10487_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10138_/Y sky130_fd_sc_hd__nand2_1
XFILLER_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10069_ _10069_/A _10069_/B _10140_/B vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__and3_1
XFILLER_63_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07732__A _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06300_ _06262_/A _06304_/A _06304_/B vssd1 vssd1 vccd1 vccd1 _06303_/A sky130_fd_sc_hd__a21bo_1
X_07280_ _07280_/A _07280_/B _07280_/C _07289_/A vssd1 vssd1 vccd1 vccd1 _07282_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__08563__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06231_ _10606_/Q _06236_/B vssd1 vssd1 vccd1 vccd1 _06231_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_76_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08282__B _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09251__A0 _08287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06162_ input44/X vssd1 vssd1 vccd1 vccd1 _10535_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_129_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06093_ _08236_/A vssd1 vssd1 vccd1 vccd1 _08062_/A sky130_fd_sc_hd__buf_2
XFILLER_160_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09921_ _09921_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _10065_/D sky130_fd_sc_hd__nor2_2
XFILLER_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09852_ _09852_/A _09852_/B vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__nor2_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08762__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08803_ _08777_/A _08803_/B _08803_/C _08803_/D vssd1 vssd1 vccd1 vccd1 _08804_/D
+ sky130_fd_sc_hd__and4b_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _09713_/B _09718_/Y _09781_/Y _09780_/X vssd1 vssd1 vccd1 vccd1 _09784_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _09344_/B vssd1 vssd1 vccd1 vccd1 _07008_/A sky130_fd_sc_hd__buf_2
XFILLER_100_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08734_ _08928_/B vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__buf_2
X_05946_ _08339_/A _05947_/B _05836_/X _08332_/A _05945_/X vssd1 vssd1 vccd1 vccd1
+ _05946_/X sky130_fd_sc_hd__a221o_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _10832_/Q _10764_/Q vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__xnor2_1
X_05877_ _05877_/A vssd1 vssd1 vccd1 vccd1 _05877_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_53_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07616_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _07616_/X sky130_fd_sc_hd__or2_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09609__A2 _09610_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08596_ _08623_/C vssd1 vssd1 vccd1 vccd1 _08597_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07547_ _07743_/A _07547_/B vssd1 vssd1 vccd1 vccd1 _07549_/B sky130_fd_sc_hd__or2_1
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07478_ _07477_/A _07477_/B _07480_/A _07480_/B vssd1 vssd1 vccd1 vccd1 _07497_/B
+ sky130_fd_sc_hd__o2bb2ai_1
XANTENNA__09349__A_N _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09217_ _09228_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09218_/A sky130_fd_sc_hd__and2_2
XFILLER_155_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06429_ _06630_/A _06407_/B _06425_/Y _06656_/A vssd1 vssd1 vccd1 vccd1 _06430_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__10508__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08045__A1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09148_ _09148_/A vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09079_ _09079_/A vssd1 vssd1 vccd1 vccd1 _09079_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input13_A io_wbs_m2s_addr[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06168__A _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10825_ _10830_/CLK _10825_/D vssd1 vssd1 vccd1 vccd1 _10825_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09481__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _10792_/CLK _10756_/D vssd1 vssd1 vccd1 vccd1 _10756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10687_ _10987_/CLK _10687_/D vssd1 vssd1 vccd1 vccd1 _10687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09233__A0 _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output81_A _10837_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07727__A _07727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05800_ _05717_/D _05799_/X _05708_/B vssd1 vssd1 vccd1 vccd1 _05800_/X sky130_fd_sc_hd__o21a_1
X_06780_ _06781_/A _06781_/B vssd1 vssd1 vccd1 vccd1 _06782_/A sky130_fd_sc_hd__and2_1
XFILLER_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05731_ _05728_/X _05729_/Y _05547_/A _08093_/A vssd1 vssd1 vccd1 vccd1 _05732_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05662_ _08169_/A _05617_/X _05619_/X _05885_/A _05661_/X vssd1 vssd1 vccd1 vccd1
+ _05662_/X sky130_fd_sc_hd__a221o_1
X_08450_ _08460_/A _08450_/B vssd1 vssd1 vccd1 vccd1 _08451_/A sky130_fd_sc_hd__or2_1
XFILLER_91_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07401_ _07070_/A _07359_/A _07398_/B _07562_/A vssd1 vssd1 vccd1 vccd1 _07402_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08381_ _08381_/A _10750_/Q vssd1 vssd1 vccd1 vccd1 _08381_/X sky130_fd_sc_hd__or2_1
X_05593_ _05593_/A _05593_/B vssd1 vssd1 vccd1 vccd1 _05593_/X sky130_fd_sc_hd__and2_1
XFILLER_91_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07332_ _07333_/A _07333_/B vssd1 vssd1 vccd1 vccd1 _07525_/A sky130_fd_sc_hd__or2b_1
XFILLER_52_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07263_ _07334_/A _07195_/A _07262_/X vssd1 vssd1 vccd1 vccd1 _07268_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10973__D _10973_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09002_ _10964_/Q vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_06214_ _10599_/Q _06223_/B vssd1 vssd1 vccd1 vccd1 _06214_/X sky130_fd_sc_hd__or2_1
X_07194_ _07194_/A _07194_/B vssd1 vssd1 vccd1 vccd1 _07210_/A sky130_fd_sc_hd__xnor2_1
XFILLER_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06145_ _06145_/A _06145_/B vssd1 vssd1 vccd1 vccd1 _06145_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06076_ _05781_/Y _05844_/A _08256_/A _05751_/Y vssd1 vssd1 vccd1 vccd1 _06076_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_160_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _09904_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _09905_/B sky130_fd_sc_hd__nand2_1
XFILLER_99_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _09837_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input5_A io_wbs_m2s_addr[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09766_ _09842_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__or2_1
XFILLER_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06978_ _10902_/Q vssd1 vssd1 vccd1 vccd1 _07056_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08717_ _08801_/B vssd1 vssd1 vccd1 vccd1 _08856_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05929_ _05877_/X _05878_/Y _05876_/X _08206_/A _05928_/X vssd1 vssd1 vccd1 vccd1
+ _05929_/X sky130_fd_sc_hd__a221o_1
X_09697_ _09588_/A _09640_/A _09639_/B _09769_/B vssd1 vssd1 vccd1 vccd1 _09767_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_26_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08648_ _10797_/Q _08648_/B vssd1 vssd1 vccd1 vccd1 _08649_/C sky130_fd_sc_hd__nand2_1
XFILLER_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08579_ _10778_/Q _08578_/C _08578_/D _10779_/Q vssd1 vssd1 vccd1 vccd1 _08580_/C
+ sky130_fd_sc_hd__a31o_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09299__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10610_ _10643_/CLK _10610_/D vssd1 vssd1 vccd1 vccd1 _10610_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08634__C _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10541_ _10654_/CLK _10541_/D vssd1 vssd1 vccd1 vccd1 _10541_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09215__A0 _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10472_ _10962_/Q _10472_/B vssd1 vssd1 vccd1 vccd1 _10472_/X sky130_fd_sc_hd__or2_1
XFILLER_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06029__B1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10808_ _10942_/CLK _10808_/D vssd1 vssd1 vccd1 vccd1 _10808_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10739_ _10788_/CLK _10739_/D vssd1 vssd1 vccd1 vccd1 _10739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08980__A2 _06212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _07950_/A vssd1 vssd1 vccd1 vccd1 _07983_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_114_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06901_ _10504_/A _07776_/B _06773_/C vssd1 vssd1 vccd1 vccd1 _06902_/B sky130_fd_sc_hd__a21oi_1
X_07881_ _07899_/A vssd1 vssd1 vccd1 vccd1 _07898_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_110_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__xnor2_1
XFILLER_110_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06832_ _06832_/A _06794_/B vssd1 vssd1 vccd1 vccd1 _06833_/B sky130_fd_sc_hd__or2b_1
XFILLER_96_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09551_ _09867_/B _09760_/B vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06763_ _06763_/A _06763_/B vssd1 vssd1 vccd1 vccd1 _06765_/B sky130_fd_sc_hd__xor2_1
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08502_ _10177_/A vssd1 vssd1 vccd1 vccd1 _08502_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05714_ _05709_/Y _10551_/Q _10550_/Q _05711_/Y _05713_/X vssd1 vssd1 vccd1 vccd1
+ _05714_/X sky130_fd_sc_hd__a221o_1
X_09482_ _09479_/Y _09481_/X _10870_/Q _09406_/X vssd1 vssd1 vccd1 vccd1 _10870_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06694_ _06915_/B _06942_/A _06915_/A vssd1 vssd1 vccd1 vccd1 _06916_/A sky130_fd_sc_hd__o21a_2
XFILLER_24_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _10218_/A _08661_/A _08432_/Y vssd1 vssd1 vccd1 vccd1 _08476_/S sky130_fd_sc_hd__a21oi_2
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05645_ _10681_/Q vssd1 vssd1 vccd1 vccd1 _08082_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05576_ _05576_/A _05576_/B vssd1 vssd1 vccd1 vccd1 _05576_/X sky130_fd_sc_hd__and2_1
X_08364_ _08364_/A vssd1 vssd1 vccd1 vccd1 _10711_/D sky130_fd_sc_hd__clkbuf_1
X_07315_ _07347_/A _07347_/B vssd1 vssd1 vccd1 vccd1 _07470_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09996__A1 _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08799__A2 _08785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09996__B2 _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08295_ _10704_/Q _10703_/Q _08295_/C vssd1 vssd1 vccd1 vccd1 _08315_/C sky130_fd_sc_hd__and3_1
X_07246_ _07246_/A _07246_/B vssd1 vssd1 vccd1 vccd1 _07247_/B sky130_fd_sc_hd__or2_1
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07177_ _07200_/A _07200_/B _07176_/A vssd1 vssd1 vccd1 vccd1 _07183_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06128_ _09250_/A vssd1 vssd1 vccd1 vccd1 _06129_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__08420__A1 _06143_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06059_ _08232_/A _08235_/A _07991_/A _05877_/X vssd1 vssd1 vccd1 vccd1 _06059_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_132_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09818_ _09819_/A _09819_/B vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__and2_1
XANTENNA__08198__A _08198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09749_ _09749_/A _09749_/B vssd1 vssd1 vccd1 vccd1 _09750_/B sky130_fd_sc_hd__and2_1
XFILLER_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08926__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10294__A1 _07008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07830__A _10577_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08239__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08239__B2 _08233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput18 io_wbs_m2s_data[11] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_2
XFILLER_156_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput29 io_wbs_m2s_data[21] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09757__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10524_ input27/X _10531_/B _10533_/C vssd1 vssd1 vccd1 vccd1 _10524_/X sky130_fd_sc_hd__or3_1
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08661__A _08661_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ _06172_/X _10446_/X _10454_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10955_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _10531_/A _10394_/B _10394_/C vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__and3_1
XFILLER_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05430_ _07885_/A _05350_/X _05346_/X _10636_/Q _05429_/X vssd1 vssd1 vccd1 vccd1
+ _05430_/X sky130_fd_sc_hd__o221a_1
XFILLER_159_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05361_ _10631_/Q vssd1 vssd1 vccd1 vccd1 _07871_/A sky130_fd_sc_hd__buf_2
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07100_ _07235_/B vssd1 vssd1 vccd1 vccd1 _07327_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _08098_/B _08079_/Y _06117_/D vssd1 vssd1 vccd1 vccd1 _08080_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05292_ _05277_/Y _05398_/A _05397_/B vssd1 vssd1 vccd1 vccd1 _05391_/B sky130_fd_sc_hd__a21o_1
XFILLER_146_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07031_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07042_/B sky130_fd_sc_hd__nor2_1
XFILLER_146_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08982_ _05475_/X _08976_/X _08979_/X _08980_/Y _09078_/B vssd1 vssd1 vccd1 vccd1
+ _08982_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07933_ _09124_/B _09092_/A vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07864_ _07848_/X _05460_/C _07844_/X _07863_/Y vssd1 vssd1 vccd1 vccd1 _10629_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__05519__A2 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09603_ _09610_/B _09610_/C vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__and2_1
X_06815_ _07780_/C _07766_/B vssd1 vssd1 vccd1 vccd1 _07779_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07795_ _06719_/B _06718_/A _06718_/B _07791_/A vssd1 vssd1 vccd1 vccd1 _07795_/X
+ sky130_fd_sc_hd__a31o_1
X_09534_ _10968_/Q _09579_/A _09534_/C vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__and3_1
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06746_ _06746_/A _06746_/B vssd1 vssd1 vccd1 vccd1 _06776_/A sky130_fd_sc_hd__xnor2_2
XFILLER_25_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09465_ _09552_/B _09466_/B vssd1 vssd1 vccd1 vccd1 _09516_/A sky130_fd_sc_hd__nor2_1
X_06677_ _06678_/A _06678_/B _06678_/C vssd1 vssd1 vccd1 vccd1 _06943_/B sky130_fd_sc_hd__nand3_1
XFILLER_25_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08416_ _08416_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__and2_1
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05628_ _10549_/Q _05630_/A vssd1 vssd1 vccd1 vccd1 _05628_/X sky130_fd_sc_hd__xor2_1
X_09396_ _09396_/A _09396_/B _09396_/C vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__nand3_1
X_08347_ _08347_/A vssd1 vssd1 vccd1 vccd1 _10709_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05559_ _10563_/Q _05596_/A vssd1 vssd1 vccd1 vccd1 _05593_/A sky130_fd_sc_hd__or2_1
XFILLER_137_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08278_ _08278_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08278_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07229_ _07229_/A _07229_/B _07244_/A vssd1 vssd1 vccd1 vccd1 _07231_/B sky130_fd_sc_hd__and3_1
XFILLER_164_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10240_ _10246_/C _10238_/X _10239_/Y vssd1 vssd1 vccd1 vccd1 _10240_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10171_ _07747_/A _10167_/X _10170_/X _10884_/Q vssd1 vssd1 vccd1 vccd1 _10884_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08656__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A _07560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06176__A _10343_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10507_ _06147_/X _10496_/X _10506_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10974_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10438_ _06143_/X _10440_/B _05977_/X vssd1 vssd1 vccd1 vccd1 _10438_/X sky130_fd_sc_hd__a21o_1
XFILLER_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10369_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__and2_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06600_ _06600_/A vssd1 vssd1 vccd1 vccd1 _06775_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07580_ _07580_/A _07580_/B vssd1 vssd1 vccd1 vccd1 _07581_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06531_ _06521_/A _06519_/A _06507_/A vssd1 vssd1 vccd1 vccd1 _06532_/B sky130_fd_sc_hd__o21bai_2
X_09250_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09276_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_33_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06462_ _06470_/A _06462_/B vssd1 vssd1 vccd1 vccd1 _06479_/B sky130_fd_sc_hd__xor2_1
XFILLER_167_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08201_ _08201_/A vssd1 vssd1 vccd1 vccd1 _08201_/X sky130_fd_sc_hd__clkbuf_2
X_05413_ _10620_/Q _05487_/A _05485_/A _10619_/Q _05412_/X vssd1 vssd1 vccd1 vccd1
+ _05413_/X sky130_fd_sc_hd__o221a_1
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06393_ _06393_/A _06393_/B vssd1 vssd1 vccd1 vccd1 _06394_/B sky130_fd_sc_hd__xor2_1
X_09181_ _07988_/A _09226_/S _09203_/A _09180_/X vssd1 vssd1 vccd1 vccd1 _09181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05344_ _10636_/Q vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08132_ _08132_/A _08132_/B vssd1 vssd1 vccd1 vccd1 _08132_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_147_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10981__D _10981_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05275_ _10652_/Q vssd1 vssd1 vccd1 vccd1 _05291_/A sky130_fd_sc_hd__clkinv_2
XFILLER_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08063_ _08075_/B _08072_/B _08306_/B _08062_/X vssd1 vssd1 vccd1 vccd1 _08063_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07014_ _07039_/C vssd1 vssd1 vccd1 vccd1 _07434_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_89_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08965_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08965_/Y sky130_fd_sc_hd__nor2_4
XFILLER_25_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07916_ _07916_/A _07916_/B vssd1 vssd1 vccd1 vccd1 _10643_/D sky130_fd_sc_hd__nor2_1
XANTENNA__10071__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08896_ hold12/A _08902_/B vssd1 vssd1 vccd1 vccd1 _08896_/X sky130_fd_sc_hd__xor2_1
XFILLER_29_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07847_ _07827_/X _05461_/C _07844_/X _07846_/Y vssd1 vssd1 vccd1 vccd1 _10625_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07778_ _07778_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07787_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09517_ _09516_/B _09516_/C _09516_/A vssd1 vssd1 vccd1 vccd1 _09562_/C sky130_fd_sc_hd__a21o_1
X_06729_ _06729_/A _06729_/B vssd1 vssd1 vccd1 vccd1 _06752_/A sky130_fd_sc_hd__xnor2_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08311__B1 _08088_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09448_/A _09448_/B vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__xnor2_4
XFILLER_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08862__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09379_ _10896_/Q _09379_/B vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__and2b_1
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10223_ _10224_/A _10935_/Q vssd1 vssd1 vccd1 vccd1 _10225_/A sky130_fd_sc_hd__nor2_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10185__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07555__A _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A io_wbs_m2s_data[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10154_ _10154_/A _10154_/B vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__xnor2_1
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__nand2_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10488__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10987_ _10987_/CLK _10987_/D vssd1 vssd1 vccd1 vccd1 _10987_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_128_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08853__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09030__B2 _10933_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08747_/X _08749_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10807_/D sky130_fd_sc_hd__o21a_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05962_ input10/X _09142_/B vssd1 vssd1 vccd1 vccd1 _07967_/A sky130_fd_sc_hd__or2_2
XFILLER_39_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07701_ _09759_/A _09759_/B _07700_/Y vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08681_ _08679_/X _08680_/Y _08669_/B _08670_/C vssd1 vssd1 vccd1 vccd1 _08683_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_39_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05893_ _10656_/Q vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_26_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07632_ _07715_/D _07632_/B vssd1 vssd1 vccd1 vccd1 _07633_/B sky130_fd_sc_hd__nand2_1
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08296__A _08297_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06809__A _10911_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10976__D _10976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07563_ _07563_/A _07727_/B _07563_/C vssd1 vssd1 vccd1 vccd1 _07563_/X sky130_fd_sc_hd__and3_1
XFILLER_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09302_ _10497_/A _09302_/B vssd1 vssd1 vccd1 vccd1 _09303_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06514_ _06527_/A _06522_/B _06517_/B _06567_/A vssd1 vssd1 vccd1 vccd1 _06523_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07494_ _07508_/B _07508_/A vssd1 vssd1 vccd1 vccd1 _07506_/A sky130_fd_sc_hd__or2b_1
X_09233_ _08256_/A _09231_/X _09257_/S vssd1 vssd1 vccd1 vccd1 _09233_/X sky130_fd_sc_hd__mux2_1
X_06445_ _10975_/Q _06576_/B vssd1 vssd1 vccd1 vccd1 _06675_/A sky130_fd_sc_hd__nand2_1
XFILLER_148_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _10959_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09164_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06376_ _06517_/B vssd1 vssd1 vccd1 vccd1 _06513_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08115_ _08115_/A _08115_/B vssd1 vssd1 vccd1 vccd1 _08130_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10403__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05327_ _10643_/Q vssd1 vssd1 vccd1 vccd1 _07914_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09095_ _09769_/A vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08046_ _08212_/A vssd1 vssd1 vccd1 vccd1 _08248_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09021__A1 _06066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09997_ _10138_/B _09997_/B vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08948_ _08968_/A vssd1 vssd1 vccd1 vccd1 _08948_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_103_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08879_ input32/X _08830_/X _08831_/X _08876_/A vssd1 vssd1 vccd1 vccd1 _08879_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10255__A_N _10938_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08918__B _08918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10910_ _10925_/CLK _10910_/D vssd1 vssd1 vccd1 vccd1 _10910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _10856_/CLK _10841_/D vssd1 vssd1 vccd1 vccd1 _10841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10772_ _10807_/CLK _10772_/D vssd1 vssd1 vccd1 vccd1 _10772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _10197_/A _10196_/B _10204_/X vssd1 vssd1 vccd1 vccd1 _10206_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_95_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ _10137_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10144_/A sky130_fd_sc_hd__xnor2_1
XFILLER_67_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10068_ _10068_/A _10068_/B vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06230_ input29/X _06225_/X _06229_/X _06221_/X vssd1 vssd1 vccd1 vccd1 _10605_/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_43_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10674_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_157_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06161_ _05982_/A _06158_/X _06160_/Y _06153_/X vssd1 vssd1 vccd1 vccd1 _10589_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06092_ _08037_/A vssd1 vssd1 vccd1 vccd1 _06117_/C sky130_fd_sc_hd__buf_2
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09920_ _10894_/Q _09920_/B vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__and2b_1
XFILLER_131_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10554_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09851_ _09851_/A _09851_/B _09851_/C vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__nor3_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08211__C1 _06020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10333__B _10946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _10815_/Q _08856_/B vssd1 vssd1 vccd1 vccd1 _08802_/Y sky130_fd_sc_hd__nor2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09782_ _09780_/X _09781_/Y _09718_/Y _09713_/B vssd1 vssd1 vccd1 vccd1 _09784_/A
+ sky130_fd_sc_hd__a211oi_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06994_ _10909_/Q vssd1 vssd1 vccd1 vccd1 _07028_/A sky130_fd_sc_hd__buf_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10840__CLK _10840_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08733_ _08918_/B vssd1 vssd1 vccd1 vccd1 _08928_/B sky130_fd_sc_hd__buf_2
XFILLER_67_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05945_ _08324_/A _05839_/X _05836_/X _08339_/B _05944_/X vssd1 vssd1 vccd1 vccd1
+ _05945_/X sky130_fd_sc_hd__o221a_1
XFILLER_22_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _08778_/A vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05876_ _05848_/B _05823_/A _05875_/Y vssd1 vssd1 vccd1 vccd1 _05876_/X sky130_fd_sc_hd__o21a_1
XFILLER_26_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07615_ _07615_/A _07615_/B vssd1 vssd1 vccd1 vccd1 _09898_/B sky130_fd_sc_hd__xnor2_4
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08595_ _10784_/Q _10783_/Q vssd1 vssd1 vccd1 vccd1 _08623_/C sky130_fd_sc_hd__and2_1
XFILLER_54_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07546_ _07545_/B _07546_/B vssd1 vssd1 vccd1 vccd1 _07547_/B sky130_fd_sc_hd__and2b_1
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07477_ _07477_/A _07477_/B vssd1 vssd1 vccd1 vccd1 _07480_/B sky130_fd_sc_hd__xnor2_1
X_09216_ _10816_/Q _09210_/X _09212_/X _09203_/X _09215_/X vssd1 vssd1 vccd1 vccd1
+ _09217_/B sky130_fd_sc_hd__a32o_1
XFILLER_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06428_ _06800_/A _06428_/B _06690_/A vssd1 vssd1 vccd1 vccd1 _06656_/A sky130_fd_sc_hd__and3_1
X_09147_ _09113_/X _09146_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09147_/Y sky130_fd_sc_hd__o21ai_1
X_06359_ _09302_/B _06736_/A vssd1 vssd1 vccd1 vccd1 _06359_/Y sky130_fd_sc_hd__nor2_1
XFILLER_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09078_ _09078_/A _09078_/B vssd1 vssd1 vccd1 vccd1 _09078_/Y sky130_fd_sc_hd__nand2_1
X_08029_ _08029_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10524__A input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10824_ _10830_/CLK _10824_/D vssd1 vssd1 vccd1 vccd1 _10824_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10755_ _10784_/CLK _10755_/D vssd1 vssd1 vccd1 vccd1 _10755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_20_clock_A _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10686_ _10987_/CLK _10686_/D vssd1 vssd1 vccd1 vccd1 _10686_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_173_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05528__A _05528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05730_ _08095_/A vssd1 vssd1 vccd1 vccd1 _08093_/A sky130_fd_sc_hd__buf_2
XFILLER_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05661_ _08169_/B _05623_/X _05617_/X _08169_/A _05660_/X vssd1 vssd1 vccd1 vccd1
+ _05661_/X sky130_fd_sc_hd__o221a_1
XFILLER_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ _07406_/A _07753_/A _07399_/X vssd1 vssd1 vccd1 vccd1 _07404_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08380_ _08394_/A vssd1 vssd1 vccd1 vccd1 _08380_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05592_ _10563_/Q _05596_/A vssd1 vssd1 vccd1 vccd1 _05593_/B sky130_fd_sc_hd__nand2_1
XFILLER_32_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07331_ _07331_/A _07331_/B vssd1 vssd1 vccd1 vccd1 _07333_/B sky130_fd_sc_hd__and2_1
XFILLER_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07262_ _07169_/A _07197_/B _07186_/B _07166_/A vssd1 vssd1 vccd1 vccd1 _07262_/X
+ sky130_fd_sc_hd__a22o_1
X_09001_ _10713_/Q _08990_/C _09000_/X vssd1 vssd1 vccd1 vccd1 _09001_/X sky130_fd_sc_hd__o21a_2
X_06213_ _06253_/B vssd1 vssd1 vccd1 vccd1 _06223_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07193_ _07193_/A _07193_/B vssd1 vssd1 vccd1 vccd1 _07194_/A sky130_fd_sc_hd__nand2_1
XFILLER_118_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07918__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06144_ _10586_/Q vssd1 vssd1 vccd1 vccd1 _06145_/A sky130_fd_sc_hd__inv_2
XFILLER_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06075_ _10677_/Q vssd1 vssd1 vccd1 vccd1 _08029_/A sky130_fd_sc_hd__inv_2
XFILLER_116_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09903_ _09903_/A vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_99_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09834_ _09834_/A _09834_/B _09977_/B _09903_/A vssd1 vssd1 vccd1 vccd1 _09835_/B
+ sky130_fd_sc_hd__and4_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09765_ _09763_/C _09829_/A vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__and2b_1
X_06977_ _10903_/Q vssd1 vssd1 vccd1 vccd1 _07066_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08716_ _08789_/B vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_27_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05928_ _08188_/A _05884_/Y _05878_/Y _05877_/A _05927_/X vssd1 vssd1 vccd1 vccd1
+ _05928_/X sky130_fd_sc_hd__o221a_1
X_09696_ _09696_/A vssd1 vssd1 vccd1 vccd1 _09769_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__B1 _09127_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _10796_/Q _08600_/A _08643_/C _10797_/Q vssd1 vssd1 vccd1 vccd1 _08649_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05859_ _10668_/Q _05863_/B vssd1 vssd1 vccd1 vccd1 _05859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _10779_/Q _10778_/Q _08578_/C _08578_/D vssd1 vssd1 vccd1 vccd1 _08585_/C
+ sky130_fd_sc_hd__and4_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _07529_/A _07529_/B vssd1 vssd1 vccd1 vccd1 _07639_/A sky130_fd_sc_hd__or2_1
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _10728_/CLK _10540_/D vssd1 vssd1 vccd1 vccd1 _10540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ _06202_/X _10459_/X _10469_/X _10470_/X vssd1 vssd1 vccd1 vccd1 _10961_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_108_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06029__A1 _10412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06201__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A _07563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08394__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05811__A _05818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _10807_/CLK _10807_/D vssd1 vssd1 vccd1 vccd1 _10807_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10738_ _10776_/CLK _10738_/D vssd1 vssd1 vccd1 vccd1 _10738_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08662__C1 _09090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10669_ _10671_/CLK _10669_/D vssd1 vssd1 vccd1 vccd1 _10669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06900_ _06900_/A vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__buf_2
X_07880_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _10633_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08193__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08193__B2 _08191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06831_ _06875_/A _06875_/B vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__and2b_1
XFILLER_28_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09550_ _09610_/C vssd1 vssd1 vccd1 vccd1 _09760_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06762_ _06762_/A _06762_/B vssd1 vssd1 vccd1 vccd1 _06763_/B sky130_fd_sc_hd__xor2_2
XFILLER_37_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08501_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10177_/A sky130_fd_sc_hd__clkbuf_4
X_05713_ _10549_/Q _08139_/A _08146_/A _05712_/Y vssd1 vssd1 vccd1 vccd1 _05713_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_09481_ _09479_/A _09479_/B _09480_/X vssd1 vssd1 vccd1 vccd1 _09481_/X sky130_fd_sc_hd__a21o_1
X_06693_ _06693_/A _06693_/B vssd1 vssd1 vccd1 vccd1 _06915_/A sky130_fd_sc_hd__xor2_1
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08432_ _08432_/A _08432_/B _08578_/C vssd1 vssd1 vccd1 vccd1 _08432_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05644_ _05913_/A _05644_/B vssd1 vssd1 vccd1 vccd1 _05644_/Y sky130_fd_sc_hd__nand2_1
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06817__A _07670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10984__D _10984_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08363_ _08363_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08364_/A sky130_fd_sc_hd__and2_1
X_05575_ _10568_/Q _05769_/A _05582_/B _10569_/Q vssd1 vssd1 vccd1 vccd1 _05576_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07314_ _07344_/A _07344_/B _07345_/B _07313_/A vssd1 vssd1 vccd1 vccd1 _07347_/B
+ sky130_fd_sc_hd__a31o_1
X_08294_ _08294_/A vssd1 vssd1 vccd1 vccd1 _10703_/D sky130_fd_sc_hd__clkbuf_1
X_07245_ _07264_/A _07264_/B _07269_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07254_/A
+ sky130_fd_sc_hd__a211o_1
X_07176_ _07176_/A _07176_/B vssd1 vssd1 vccd1 vccd1 _07200_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06552__A _10971_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07759__A1 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06127_ input9/X _10432_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__and3_4
XFILLER_118_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06058_ _10666_/Q vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__buf_2
XFILLER_160_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08184__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08184__B2 _08180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__xnor2_1
XFILLER_86_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08198__B _08235_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ _09749_/A _09749_/B vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__nor2_2
XFILLER_74_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09679_/A _09679_/B vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__xor2_4
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput19 io_wbs_m2s_data[12] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_6
X_10523_ _10523_/A vssd1 vssd1 vccd1 vccd1 _10533_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10454_ _10955_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10454_/X sky130_fd_sc_hd__or2_1
XFILLER_109_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10385_ _10365_/X _10715_/Q _10383_/X _10384_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10934_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05360_ _06052_/A _05848_/B vssd1 vssd1 vccd1 vccd1 _05360_/X sky130_fd_sc_hd__xor2_2
XFILLER_158_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07989__A1 _06195_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05291_ _05291_/A _10576_/Q vssd1 vssd1 vccd1 vccd1 _05397_/B sky130_fd_sc_hd__nor2_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07030_ _07169_/A _07166_/A _07030_/C _07417_/A vssd1 vssd1 vccd1 vccd1 _07031_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_162_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08981_ _08981_/A vssd1 vssd1 vccd1 vccd1 _09078_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07932_ _09016_/A _09013_/A vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__or2_1
XFILLER_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10979__D _10979_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07863_ _06197_/A _07849_/X _07850_/X _07862_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ _07863_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_111_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09602_ _09780_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__nand2_1
X_06814_ _06814_/A _06853_/B vssd1 vssd1 vccd1 vccd1 _07766_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07794_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07796_/B sky130_fd_sc_hd__nor2_1
X_09533_ _10967_/Q _09533_/B _09533_/C vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__and3_1
X_06745_ _07675_/A _06745_/B vssd1 vssd1 vccd1 vccd1 _06746_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09464_ _09501_/A _09464_/B vssd1 vssd1 vccd1 vccd1 _09466_/B sky130_fd_sc_hd__or2_1
XFILLER_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06676_ _06674_/A _06674_/C _06681_/A vssd1 vssd1 vccd1 vccd1 _06678_/C sky130_fd_sc_hd__a21o_1
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08415_ input1/X input49/X input14/X _08415_/D vssd1 vssd1 vccd1 vccd1 _08989_/B
+ sky130_fd_sc_hd__and4_1
X_05627_ _10688_/Q vssd1 vssd1 vccd1 vccd1 _05896_/A sky130_fd_sc_hd__clkbuf_2
X_09395_ _09678_/A vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08346_ _08344_/X _08346_/B vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__and2b_1
X_05558_ _10562_/Q _10561_/Q _05602_/A vssd1 vssd1 vccd1 vccd1 _05596_/A sky130_fd_sc_hd__or3_1
X_08277_ _08277_/A _08277_/B _08277_/C vssd1 vssd1 vccd1 vccd1 _08295_/C sky130_fd_sc_hd__and3_1
XFILLER_138_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05489_ _05489_/A vssd1 vssd1 vccd1 vccd1 _05489_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_67_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07228_ _07232_/A _07232_/B _07225_/X vssd1 vssd1 vccd1 vccd1 _07231_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07378__A _07728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07159_ _07229_/A _07164_/B _07178_/A _07188_/A vssd1 vssd1 vccd1 vccd1 _07159_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_145_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10170_ _10177_/A vssd1 vssd1 vccd1 vccd1 _10170_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08002__A _08015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10506_ _10506_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10506_/X sky130_fd_sc_hd__or2_1
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10437_ _06008_/X _10431_/X _10436_/X _08563_/X vssd1 vssd1 vccd1 vccd1 _10948_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_152_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10931_/Q _10379_/B vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__and2_1
XFILLER_151_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10442__A _10498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10299_ _10301_/A _10289_/X _10300_/A vssd1 vssd1 vccd1 vccd1 _10299_/X sky130_fd_sc_hd__o21ba_1
XFILLER_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06530_ _06541_/C _06528_/Y _06529_/X vssd1 vssd1 vccd1 vccd1 _06533_/A sky130_fd_sc_hd__o21ai_1
XFILLER_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08320__A1 _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08320__B2 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06461_ _06472_/A _06461_/B _06547_/C vssd1 vssd1 vccd1 vccd1 _06462_/B sky130_fd_sc_hd__and3b_1
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08200_ _08114_/X _08207_/B _08196_/X _08199_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08200_/X sky130_fd_sc_hd__o311a_1
X_05412_ _10619_/Q _05485_/A _05402_/X _05411_/X vssd1 vssd1 vccd1 vccd1 _05412_/X
+ sky130_fd_sc_hd__a22o_1
X_09180_ _05460_/C _09136_/X _09148_/X _08191_/A _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09180_/X sky130_fd_sc_hd__a221o_1
X_06392_ _10515_/A _06627_/B vssd1 vssd1 vccd1 vccd1 _06393_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08131_ _08092_/X _08129_/X _08139_/B _08096_/X vssd1 vssd1 vccd1 vccd1 _08131_/X
+ sky130_fd_sc_hd__a31o_1
X_05343_ _08013_/A _05854_/A vssd1 vssd1 vccd1 vccd1 _05343_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08084__B1 _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08062_ _08062_/A vssd1 vssd1 vccd1 vccd1 _08062_/X sky130_fd_sc_hd__buf_4
XFILLER_119_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05274_ _10654_/Q vssd1 vssd1 vccd1 vccd1 _05388_/A sky130_fd_sc_hd__clkinv_2
XFILLER_146_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07013_ _07013_/A _07013_/B vssd1 vssd1 vccd1 vccd1 _07039_/C sky130_fd_sc_hd__xnor2_2
XFILLER_161_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08964_ _08964_/A vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07915_ _10611_/Q _07906_/X _07910_/X _07914_/Y vssd1 vssd1 vccd1 vccd1 _07916_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_57_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08895_ _08893_/X _08894_/X _08780_/X vssd1 vssd1 vccd1 vccd1 _10825_/D sky130_fd_sc_hd__o21a_1
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07846_ _06180_/A _07828_/X _07829_/X _07845_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07846_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_56_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07777_ _07777_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07778_/B sky130_fd_sc_hd__xnor2_1
XFILLER_84_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09516_ _09516_/A _09516_/B _09516_/C vssd1 vssd1 vccd1 vccd1 _09562_/B sky130_fd_sc_hd__nand3_1
X_06728_ _06734_/A _06734_/B _06320_/Y _06321_/A vssd1 vssd1 vccd1 vccd1 _06729_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06277__A _10898_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08311__A1 input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09447_ _09678_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09448_/B sky130_fd_sc_hd__nand2_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06659_ _06660_/A _06660_/B vssd1 vssd1 vccd1 vccd1 _06661_/A sky130_fd_sc_hd__and2_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09378_ _09921_/B _09922_/B _10065_/B _09377_/X vssd1 vssd1 vccd1 vccd1 _10063_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_149_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08492__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08329_ _08339_/C _08329_/B vssd1 vssd1 vccd1 vccd1 _08329_/Y sky130_fd_sc_hd__nor2_1
XFILLER_137_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07822__B1 _06257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10222_ _10951_/Q vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__inv_2
XFILLER_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10185__A1 _09920_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10153_ _10153_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10154_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input36_A io_wbs_m2s_data[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10084_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__or2_1
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07571__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10986_ _10986_/CLK _10986_/D vssd1 vssd1 vccd1 vccd1 _10986_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06187__A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08853__A2 _08785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07813__B1 _06257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08081__A3 _08082_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10176__A1 _07061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05961_ input11/X input13/X input12/X vssd1 vssd1 vccd1 vccd1 _09142_/B sky130_fd_sc_hd__or3_4
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07700_ _07700_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _07700_/Y sky130_fd_sc_hd__nor2_1
X_08680_ _10801_/Q _08698_/A vssd1 vssd1 vccd1 vccd1 _08680_/Y sky130_fd_sc_hd__nor2_1
X_05892_ _08169_/B _05892_/B vssd1 vssd1 vccd1 vccd1 _05892_/X sky130_fd_sc_hd__and2_1
X_07631_ _07698_/A _07698_/B vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__xnor2_4
XFILLER_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07562_ _07562_/A _07729_/B _07562_/C vssd1 vssd1 vccd1 vccd1 _07563_/C sky130_fd_sc_hd__and3_1
XFILLER_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08829__C1 _08670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09301_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10043_/A sky130_fd_sc_hd__buf_2
X_06513_ _06527_/A _06600_/A _06522_/B _06513_/D vssd1 vssd1 vccd1 vccd1 _06532_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07493_ _07493_/A _07493_/B vssd1 vssd1 vccd1 vccd1 _07508_/A sky130_fd_sc_hd__xor2_2
XFILLER_62_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09232_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09257_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06444_ _10976_/Q _06587_/A _06947_/A vssd1 vssd1 vccd1 vccd1 _06472_/B sky130_fd_sc_hd__and3_1
XFILLER_167_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09163_ _09202_/A _09163_/B vssd1 vssd1 vccd1 vccd1 _10845_/D sky130_fd_sc_hd__nor2_4
X_06375_ _06375_/A _06387_/B vssd1 vssd1 vccd1 vccd1 _06517_/B sky130_fd_sc_hd__xnor2_4
XFILLER_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ _08263_/A vssd1 vssd1 vccd1 vccd1 _08114_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_108_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05326_ _05830_/A _05831_/B vssd1 vssd1 vccd1 vccd1 _05326_/X sky130_fd_sc_hd__xor2_2
X_09094_ _10970_/Q vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_108_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08045_ _05475_/X _08044_/X _06033_/X vssd1 vssd1 vccd1 vccd1 _08045_/X sky130_fd_sc_hd__a21o_1
XFILLER_162_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09021__A2 _06212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09996_ _10123_/A _09919_/B _10122_/B _10487_/A vssd1 vssd1 vccd1 vccd1 _09997_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08947_ _08947_/A vssd1 vssd1 vccd1 vccd1 _10430_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08878_ _08883_/A _08876_/Y _08871_/Y _08873_/Y vssd1 vssd1 vccd1 vccd1 _08878_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07829_ _07850_/A vssd1 vssd1 vccd1 vccd1 _07829_/X sky130_fd_sc_hd__buf_4
XFILLER_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10840_ _10840_/CLK _10840_/D vssd1 vssd1 vccd1 vccd1 _10840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10771_ _10782_/CLK _10771_/D vssd1 vssd1 vccd1 vccd1 _10771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06846__A1 _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09111__A _09111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08063__A3 _08306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06074__A2 _08034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _10191_/B _10204_/X _10196_/B vssd1 vssd1 vccd1 vccd1 _10226_/A sky130_fd_sc_hd__a21o_1
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08220__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _10491_/A _10129_/B _10061_/A _10059_/A vssd1 vssd1 vccd1 vccd1 _10137_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10067_ _10131_/B _10067_/B vssd1 vssd1 vccd1 vccd1 _10068_/B sky130_fd_sc_hd__xnor2_2
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10969_ _10970_/CLK _10969_/D vssd1 vssd1 vccd1 vccd1 _10969_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08039__B1 _05736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10167__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06160_ _06160_/A _06170_/B vssd1 vssd1 vccd1 vccd1 _06160_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07262__A1 _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06091_ _10580_/Q vssd1 vssd1 vccd1 vccd1 _08037_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__07262__B2 _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08333__C_N _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09850_ _09851_/A _09851_/B _09851_/C vssd1 vssd1 vccd1 vccd1 _09852_/A sky130_fd_sc_hd__o21a_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _10815_/Q _08801_/B vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__and2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09781_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09781_/Y sky130_fd_sc_hd__nand2_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _06993_/A vssd1 vssd1 vccd1 vccd1 _09920_/B sky130_fd_sc_hd__buf_2
XFILLER_112_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05944_ _05939_/X _05940_/X _05942_/X _05943_/X vssd1 vssd1 vccd1 vccd1 _05944_/X
+ sky130_fd_sc_hd__a31o_1
X_08732_ _10806_/Q _08732_/B vssd1 vssd1 vccd1 vccd1 _08740_/C sky130_fd_sc_hd__xor2_1
XFILLER_85_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10987__D _10987_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _10799_/Q _08658_/X _08662_/X vssd1 vssd1 vccd1 vccd1 _10799_/D sky130_fd_sc_hd__a21boi_1
X_05875_ _08198_/A _05878_/B _10663_/Q vssd1 vssd1 vccd1 vccd1 _05875_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10321__A1 _07570_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07614_ _07620_/A _06962_/B _07624_/A vssd1 vssd1 vccd1 vccd1 _07615_/B sky130_fd_sc_hd__a21oi_2
XFILLER_121_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _10783_/Q _08550_/X _08593_/Y vssd1 vssd1 vccd1 vccd1 _10783_/D sky130_fd_sc_hd__o21a_1
XFILLER_42_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07545_ _07546_/B _07545_/B vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__and2b_1
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07476_ _07589_/A vssd1 vssd1 vccd1 vccd1 _07480_/A sky130_fd_sc_hd__inv_2
XFILLER_139_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06427_ _06690_/A _06630_/A _06425_/Y _06428_/B _06800_/A vssd1 vssd1 vccd1 vccd1
+ _06631_/A sky130_fd_sc_hd__o2111a_1
X_09215_ _08000_/A _09214_/X _09297_/S vssd1 vssd1 vccd1 vccd1 _09215_/X sky130_fd_sc_hd__mux2_1
XFILLER_167_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09146_ _09114_/X _09145_/X _09119_/X vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__o21a_1
X_06358_ _06558_/B _06558_/C vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__nand2_2
XFILLER_147_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05309_ _10672_/Q _05340_/A vssd1 vssd1 vccd1 vccd1 _05336_/A sky130_fd_sc_hd__or2_1
X_09077_ _08119_/A _08976_/X _09076_/X _09078_/B vssd1 vssd1 vccd1 vccd1 _09077_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06289_ _10928_/Q _10911_/Q vssd1 vssd1 vccd1 vccd1 _06851_/A sky130_fd_sc_hd__or2_1
XFILLER_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08028_ input36/X _07985_/B _08027_/X _08019_/X vssd1 vssd1 vccd1 vccd1 _10676_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08202__B1 _08124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09979_ _10049_/C _09976_/Y _09978_/X vssd1 vssd1 vccd1 vccd1 _09980_/B sky130_fd_sc_hd__o21a_1
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10823_ _10830_/CLK _10823_/D vssd1 vssd1 vccd1 vccd1 _10823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10754_ _10784_/CLK _10754_/D vssd1 vssd1 vccd1 vccd1 _10754_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ _10987_/CLK _10685_/D vssd1 vssd1 vccd1 vccd1 _10685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10119_ _10107_/A _10107_/B _10118_/X vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__a21oi_2
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05660_ _08148_/A _05626_/X _05623_/X _10690_/Q _05659_/X vssd1 vssd1 vccd1 vccd1
+ _05660_/X sky130_fd_sc_hd__a221o_1
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05591_ _10702_/Q vssd1 vssd1 vccd1 vccd1 _08277_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07330_ _07330_/A _07335_/A vssd1 vssd1 vccd1 vccd1 _07331_/B sky130_fd_sc_hd__nand2_1
XFILLER_91_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07483__A1 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07261_ _07273_/A _07273_/B vssd1 vssd1 vccd1 vccd1 _07318_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07483__B2 _07715_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ _10766_/Q _08418_/B _09168_/A _10800_/Q _08999_/X vssd1 vssd1 vccd1 vccd1
+ _09000_/X sky130_fd_sc_hd__a221o_1
X_06212_ _10517_/A _06212_/B vssd1 vssd1 vccd1 vccd1 _06253_/B sky130_fd_sc_hd__nor2_4
XFILLER_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07192_ _07192_/A _07192_/B vssd1 vssd1 vccd1 vccd1 _07194_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08590__A _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06143_ _10526_/A vssd1 vssd1 vccd1 vccd1 _06143_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_133_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08983__A1 _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06074_ _10711_/Q _08034_/A _07979_/A _05709_/Y _06073_/X vssd1 vssd1 vccd1 vccd1
+ _06082_/A sky130_fd_sc_hd__a221o_1
XFILLER_133_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05797__A1 _08160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09902_ _10023_/A _09829_/A vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__or2b_1
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09833_ _09834_/A _09977_/B _09903_/A _10057_/A vssd1 vssd1 vccd1 vccd1 _09835_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09764_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06976_ _10906_/Q vssd1 vssd1 vccd1 vccd1 _06997_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08715_ _08744_/B vssd1 vssd1 vccd1 vccd1 _08789_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08499__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05927_ _10693_/Q _05884_/Y _05888_/X _05926_/X vssd1 vssd1 vccd1 vccd1 _05927_/X
+ sky130_fd_sc_hd__a22o_1
X_09695_ _09646_/B _09695_/B vssd1 vssd1 vccd1 vccd1 _09707_/A sky130_fd_sc_hd__and2b_1
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09160__A1 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05858_ _05858_/A _05858_/B vssd1 vssd1 vccd1 vccd1 _05858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08646_ _08648_/B _08646_/B vssd1 vssd1 vccd1 vccd1 _10796_/D sky130_fd_sc_hd__nor2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08577_ _08583_/A _08577_/B vssd1 vssd1 vccd1 vccd1 _10778_/D sky130_fd_sc_hd__nor2_1
X_05789_ _05789_/A _05764_/A vssd1 vssd1 vccd1 vccd1 _05789_/X sky130_fd_sc_hd__or2b_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07528_ _07528_/A _07528_/B _07528_/C vssd1 vssd1 vccd1 vccd1 _07529_/B sky130_fd_sc_hd__and3_1
XFILLER_10_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ _09304_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07460_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10470_ _10498_/A vssd1 vssd1 vccd1 vccd1 _10470_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__06029__A2 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ _08748_/X _08985_/X _08988_/X _10720_/Q _09128_/X vssd1 vssd1 vccd1 vccd1
+ _09129_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10535__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07844__A _08557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06737__B1 _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10671_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09151__B2 _10722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10806_ _10942_/CLK _10806_/D vssd1 vssd1 vccd1 vccd1 _10806_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_57_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10654_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__06195__A input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10737_ _10776_/CLK _10737_/D vssd1 vssd1 vccd1 vccd1 _10737_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05476__B1 _05474_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10668_ _10671_/CLK _10668_/D vssd1 vssd1 vccd1 vccd1 _10668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _10814_/CLK _10599_/D vssd1 vssd1 vccd1 vccd1 _10599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05779__B2 _05778_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06830_ _06844_/C _06856_/C _06884_/A vssd1 vssd1 vccd1 vccd1 _06875_/B sky130_fd_sc_hd__o21bai_2
XFILLER_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06761_ _06772_/A _06786_/A _06856_/A vssd1 vssd1 vccd1 vccd1 _06762_/B sky130_fd_sc_hd__and3b_1
XFILLER_83_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08500_ _08633_/A vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__buf_2
X_05712_ _10550_/Q vssd1 vssd1 vccd1 vccd1 _05712_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09480_ _09757_/A vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_64_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06692_ _06692_/A _06692_/B vssd1 vssd1 vccd1 vccd1 _06693_/B sky130_fd_sc_hd__xnor2_1
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05643_ _05643_/A _10541_/Q vssd1 vssd1 vccd1 vccd1 _05644_/B sky130_fd_sc_hd__xor2_1
X_08431_ _10729_/Q _08565_/C vssd1 vssd1 vccd1 vccd1 _08578_/C sky130_fd_sc_hd__and2_1
XFILLER_51_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08362_ input40/X _08123_/X _08109_/X _05528_/X _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08363_/B sky130_fd_sc_hd__o221a_1
X_05574_ _08332_/A vssd1 vssd1 vccd1 vccd1 _05574_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07313_ _07313_/A _07313_/B vssd1 vssd1 vccd1 vccd1 _07345_/B sky130_fd_sc_hd__nor2_1
X_08293_ _08291_/X _08293_/B vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__and2b_1
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07244_ _07244_/A _07244_/B vssd1 vssd1 vccd1 vccd1 _07269_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07929__A _08284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07175_ _07193_/A _07175_/B vssd1 vssd1 vccd1 vccd1 _07176_/B sky130_fd_sc_hd__nand2_1
XFILLER_118_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10355__A _10355_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06126_ input7/X input4/X _07967_/A _06126_/D vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__nor4_4
XFILLER_105_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06057_ _10668_/Q vssd1 vssd1 vccd1 vccd1 _08256_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_133_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09816_ _09961_/A _09753_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__o21a_1
XFILLER_101_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_63_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09747_ _10478_/A _09672_/B _10129_/B _09670_/Y vssd1 vssd1 vccd1 vccd1 _09749_/B
+ sky130_fd_sc_hd__a31oi_2
X_06959_ _07636_/A _07635_/B vssd1 vssd1 vccd1 vccd1 _07629_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09678_/A _09923_/B vssd1 vssd1 vccd1 vccd1 _09679_/B sky130_fd_sc_hd__nand2_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _10792_/Q _08631_/C _08642_/D _08550_/X vssd1 vssd1 vccd1 vccd1 _08630_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _10522_/A vssd1 vssd1 vccd1 vccd1 _10522_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10453_ _06168_/X _10446_/X _10452_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10954_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10384_ _10528_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10384_/X sky130_fd_sc_hd__a21bo_1
XFILLER_136_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06186__A1 _06182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06918__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05290_ _05818_/A _05910_/B _05289_/Y vssd1 vssd1 vccd1 vccd1 _05398_/A sky130_fd_sc_hd__a21oi_2
XFILLER_158_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09964__A _09964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05269__A _10679_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08980_ _05736_/A _06212_/B _08976_/X vssd1 vssd1 vccd1 vccd1 _08980_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_102_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07931_ _08944_/A _09142_/C vssd1 vssd1 vccd1 vccd1 _09013_/A sky130_fd_sc_hd__or2_1
XFILLER_29_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07862_ _10879_/Q _07866_/B vssd1 vssd1 vccd1 vccd1 _07862_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06177__A1 _06172_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09601_ _09599_/A _09692_/A _09761_/C _09805_/A vssd1 vssd1 vccd1 vccd1 _09602_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_84_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06813_ _06813_/A _06813_/B vssd1 vssd1 vccd1 vccd1 _06853_/B sky130_fd_sc_hd__xor2_2
X_07793_ _06869_/A _06869_/B _06868_/A vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__a21oi_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09532_ _09532_/A _09532_/B vssd1 vssd1 vccd1 vccd1 _09567_/A sky130_fd_sc_hd__xor2_4
X_06744_ _06775_/A _06774_/B vssd1 vssd1 vccd1 vccd1 _06747_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09463_ _09462_/A _09462_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _09464_/B sky130_fd_sc_hd__a21oi_1
X_06675_ _06675_/A _06675_/B vssd1 vssd1 vccd1 vccd1 _06678_/B sky130_fd_sc_hd__xor2_2
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08414_ _08414_/A vssd1 vssd1 vccd1 vccd1 _08415_/D sky130_fd_sc_hd__inv_2
XFILLER_169_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05626_ _05626_/A _05626_/B vssd1 vssd1 vccd1 vccd1 _05626_/X sky130_fd_sc_hd__and2_1
X_09394_ _09424_/A vssd1 vssd1 vccd1 vccd1 _09678_/A sky130_fd_sc_hd__buf_2
XFILLER_145_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08345_ input37/X _08248_/A _08052_/A _05570_/X _08175_/A vssd1 vssd1 vccd1 vccd1
+ _08346_/B sky130_fd_sc_hd__o221a_1
X_05557_ _10560_/Q _05604_/A vssd1 vssd1 vccd1 vccd1 _05602_/A sky130_fd_sc_hd__or2_1
XFILLER_20_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08276_ _08278_/A _08276_/B vssd1 vssd1 vccd1 vccd1 _08276_/Y sky130_fd_sc_hd__nor2_1
X_05488_ _05818_/B _05470_/B _05495_/A _05453_/A _05487_/Y vssd1 vssd1 vccd1 vccd1
+ _10545_/D sky130_fd_sc_hd__a221o_1
X_07227_ _07225_/X _07227_/B vssd1 vssd1 vccd1 vccd1 _07232_/B sky130_fd_sc_hd__and2b_1
XFILLER_153_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07158_ _07186_/A _07188_/A _07164_/B _07178_/A vssd1 vssd1 vccd1 vccd1 _07280_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_3_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09051__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06109_ _10705_/Q _08305_/B vssd1 vssd1 vccd1 vccd1 _08317_/B sky130_fd_sc_hd__or2_1
XFILLER_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07089_ _07089_/A _07089_/B vssd1 vssd1 vccd1 vccd1 _07090_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05915__A1 _05408_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__B _10529_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09106__A1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07569__A _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10505_ _06143_/X _10496_/X _10504_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10973_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10436_ _10948_/Q _10440_/B vssd1 vssd1 vccd1 vccd1 _10436_/X sky130_fd_sc_hd__or2_1
XFILLER_98_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10367_ _10427_/B vssd1 vssd1 vccd1 vccd1 _10379_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10298_/A _10298_/B vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__nand2_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06460_ _10978_/Q _06460_/B _06670_/A vssd1 vssd1 vccd1 vccd1 _06479_/A sky130_fd_sc_hd__and3_1
XFILLER_61_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05411_ _10618_/Q _05483_/A _05407_/X _05410_/X vssd1 vssd1 vccd1 vccd1 _05411_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06391_ _06489_/B vssd1 vssd1 vccd1 vccd1 _06627_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08130_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08139_/B sky130_fd_sc_hd__nand2_1
XFILLER_159_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05342_ _10670_/Q vssd1 vssd1 vccd1 vccd1 _08013_/A sky130_fd_sc_hd__inv_2
XFILLER_30_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09281__A0 _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08061_ _08061_/A vssd1 vssd1 vccd1 vccd1 _08306_/B sky130_fd_sc_hd__buf_2
XFILLER_88_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05273_ _10655_/Q vssd1 vssd1 vccd1 vccd1 _05295_/A sky130_fd_sc_hd__inv_2
XFILLER_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ _06997_/B _06997_/C _07007_/A vssd1 vssd1 vccd1 vccd1 _07013_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09033__A0 _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ _09092_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07914_ _07914_/A vssd1 vssd1 vccd1 vccd1 _07914_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08894_ input34/X _08830_/X _08831_/X _10825_/Q vssd1 vssd1 vccd1 vccd1 _08894_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07845_ _10875_/Q _07845_/B vssd1 vssd1 vccd1 vccd1 _07845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07776_ _10515_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07777_/B sky130_fd_sc_hd__nand2_1
XFILLER_140_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09515_ _09514_/A _09514_/B _09514_/C vssd1 vssd1 vccd1 vccd1 _09516_/C sky130_fd_sc_hd__a21o_1
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06727_ _07794_/A _07794_/B vssd1 vssd1 vccd1 vccd1 _07761_/A sky130_fd_sc_hd__xnor2_1
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _09811_/B _09677_/B vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__or2_4
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ _06658_/A _06658_/B vssd1 vssd1 vccd1 vccd1 _06660_/B sky130_fd_sc_hd__xnor2_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05609_ _10557_/Q _05612_/A vssd1 vssd1 vccd1 vccd1 _05610_/B sky130_fd_sc_hd__nand2_1
X_09377_ _10894_/Q _06993_/A vssd1 vssd1 vccd1 vccd1 _09377_/X sky130_fd_sc_hd__or2b_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06589_ _06589_/A _06589_/B vssd1 vssd1 vccd1 vccd1 _06951_/B sky130_fd_sc_hd__or2_1
XANTENNA__08492__B _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08328_ _08324_/A _08327_/B _08067_/X vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__07389__A _07728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06086__B1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ _08114_/X _08277_/C _08252_/Y _08257_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08259_/X sky130_fd_sc_hd__o311a_1
XFILLER_119_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10221_ _07113_/A _10115_/X _10220_/Y _10043_/X vssd1 vssd1 vccd1 vccd1 _10901_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _10152_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10153_/B sky130_fd_sc_hd__xnor2_1
XFILLER_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10083_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_87_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input29_A io_wbs_m2s_data[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08838__B1 _08786_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10985_ _10985_/CLK _10985_/D vssd1 vssd1 vccd1 vccd1 _10985_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09015__A0 _10502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10419_ _06191_/X _10371_/A _10415_/X vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__a21bo_1
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05960_ _10369_/A vssd1 vssd1 vccd1 vccd1 _10432_/B sky130_fd_sc_hd__buf_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05891_ _05891_/A _05891_/B vssd1 vssd1 vccd1 vccd1 _05892_/B sky130_fd_sc_hd__and2_1
XANTENNA__06001__A0 _10528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07630_ _07630_/A _07630_/B vssd1 vssd1 vccd1 vccd1 _07698_/B sky130_fd_sc_hd__xnor2_4
XFILLER_93_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07561_ _07729_/A _07728_/B vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__nand2_1
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09300_ _09300_/A vssd1 vssd1 vccd1 vccd1 _10865_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06512_ _06541_/C _06512_/B vssd1 vssd1 vccd1 vccd1 _06620_/A sky130_fd_sc_hd__xnor2_1
XFILLER_80_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09689__A _09689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07492_ _07490_/A _07490_/B _07510_/A vssd1 vssd1 vccd1 vccd1 _07508_/B sky130_fd_sc_hd__o21ba_1
XFILLER_110_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09231_ _05598_/X _07889_/A _09245_/S vssd1 vssd1 vccd1 vccd1 _09231_/X sky130_fd_sc_hd__mux2_1
X_06443_ _10975_/Q _06575_/B vssd1 vssd1 vccd1 vccd1 _06947_/A sky130_fd_sc_hd__nand2_1
XFILLER_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06374_ _06374_/A _06374_/B vssd1 vssd1 vccd1 vccd1 _06387_/B sky130_fd_sc_hd__xnor2_4
X_09162_ _09112_/X _09158_/Y _09161_/X vssd1 vssd1 vccd1 vccd1 _09163_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06068__B1 _06065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05325_ _10644_/Q vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__clkbuf_2
X_08113_ _08113_/A vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__inv_2
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09093_ _10515_/A _09118_/A vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__nor2_1
XFILLER_174_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08044_ _08044_/A vssd1 vssd1 vccd1 vccd1 _08044_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09995_ _10489_/A _10056_/C _10122_/B vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__or3b_2
XFILLER_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09309__A1 _09313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ _09124_/A _08968_/A vssd1 vssd1 vccd1 vccd1 _08947_/A sky130_fd_sc_hd__nor2_1
XFILLER_103_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08877_ _08871_/Y _08873_/Y _08883_/A _08876_/Y vssd1 vssd1 vccd1 vccd1 _08891_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07828_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07828_/X sky130_fd_sc_hd__buf_4
XFILLER_151_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07759_ _07635_/A _06966_/A _06966_/B vssd1 vssd1 vccd1 vccd1 _07764_/A sky130_fd_sc_hd__a21oi_2
X_10770_ _10770_/CLK _10770_/D vssd1 vssd1 vccd1 vccd1 _10770_/Q sky130_fd_sc_hd__dfxtp_1
X_09429_ _09429_/A _09460_/B vssd1 vssd1 vccd1 vccd1 _09430_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05757__A1_N _08242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09245__A0 _08278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08008__A _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08950__B _09142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10204_ _10948_/Q _10932_/Q vssd1 vssd1 vccd1 vccd1 _10204_/X sky130_fd_sc_hd__or2b_1
XFILLER_133_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ _10049_/B _09880_/A _09976_/Y _09879_/B vssd1 vssd1 vccd1 vccd1 _10137_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10066_ _10066_/A _10131_/C vssd1 vssd1 vccd1 vccd1 _10067_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10968_ _10968_/CLK _10968_/D vssd1 vssd1 vccd1 vccd1 _10968_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05830__A _05830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09302__A _10497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ _10980_/CLK _10899_/D vssd1 vssd1 vccd1 vccd1 _10899_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__08039__A1 _08074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_117_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06090_ _06036_/X _06071_/X _06082_/X _06089_/X _10579_/Q vssd1 vssd1 vccd1 vccd1
+ _08065_/B sky130_fd_sc_hd__o41a_4
XFILLER_129_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05277__A _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08211__A1 _08114_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08688_/X _08798_/X _08799_/X vssd1 vssd1 vccd1 vccd1 _10814_/D sky130_fd_sc_hd__o21a_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09780_ _09780_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09780_/X sky130_fd_sc_hd__or2b_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _07021_/A vssd1 vssd1 vccd1 vccd1 _07574_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08731_ _08727_/X _08730_/X _08676_/X vssd1 vssd1 vccd1 vccd1 _10805_/D sky130_fd_sc_hd__o21a_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05943_ _08315_/A _05838_/B _05941_/Y _05839_/X _08327_/A vssd1 vssd1 vccd1 vccd1
+ _05943_/X sky130_fd_sc_hd__a32o_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08662_ _06124_/A _08819_/A _08820_/A _10799_/Q _09090_/A vssd1 vssd1 vccd1 vccd1
+ _08662_/X sky130_fd_sc_hd__o221a_1
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05874_ _10661_/Q _05883_/A _05886_/A _05886_/B vssd1 vssd1 vccd1 vccd1 _05878_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07613_ _07613_/A vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__inv_2
XFILLER_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08593_ _10783_/Q _08550_/X _08630_/A vssd1 vssd1 vccd1 vccd1 _08593_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07544_ _07544_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07545_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09212__A _09275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07475_ _07728_/A _07475_/B _07475_/C vssd1 vssd1 vccd1 vccd1 _07589_/A sky130_fd_sc_hd__and3_1
XFILLER_50_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09214_ _06061_/A _07878_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09214_/X sky130_fd_sc_hd__mux2_1
X_06426_ _06426_/A vssd1 vssd1 vccd1 vccd1 _06800_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_09145_ _10941_/Q _09143_/Y _09144_/Y _08968_/X vssd1 vssd1 vccd1 vccd1 _09145_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_06357_ _06436_/A vssd1 vssd1 vccd1 vccd1 _06719_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_148_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05308_ _10671_/Q _10670_/Q _05854_/A vssd1 vssd1 vccd1 vccd1 _05340_/A sky130_fd_sc_hd__or3_1
XANTENNA__07667__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06288_ _10929_/Q _10912_/Q vssd1 vssd1 vccd1 vccd1 _06288_/X sky130_fd_sc_hd__or2_1
X_09076_ _05462_/B _09020_/B _06129_/B _08117_/A _09297_/S vssd1 vssd1 vccd1 vccd1
+ _09076_/X sky130_fd_sc_hd__o221a_1
XFILLER_162_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08027_ _08027_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08027_/X sky130_fd_sc_hd__or2_1
XFILLER_2_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08202__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08202__B2 _05877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_opt_1_0_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09978_ _09908_/A _10049_/B _10095_/A vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__07961__A0 _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _08920_/A _08927_/X _08928_/X vssd1 vssd1 vccd1 vccd1 _08929_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_130_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10822_ _10822_/CLK _10822_/D vssd1 vssd1 vccd1 vccd1 _10822_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _10784_/CLK _10753_/D vssd1 vssd1 vccd1 vccd1 _10753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10684_ _10684_/CLK _10684_/D vssd1 vssd1 vccd1 vccd1 _10684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_58_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07401__C1 _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10118_ _10104_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10118_/X sky130_fd_sc_hd__and2b_1
XFILLER_49_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08201__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10049_ _10129_/A _10049_/B _10049_/C vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__and3_1
XFILLER_64_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05590_ _10564_/Q _05593_/A vssd1 vssd1 vccd1 vccd1 _05590_/X sky130_fd_sc_hd__xor2_1
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07260_ _07260_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _07273_/B sky130_fd_sc_hd__nor2_1
XFILLER_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06211_ _09148_/A vssd1 vssd1 vccd1 vccd1 _06212_/B sky130_fd_sc_hd__buf_2
XFILLER_118_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07191_ _07229_/A _07197_/B _07186_/B _07188_/A vssd1 vssd1 vccd1 vccd1 _07193_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06142_ input38/X vssd1 vssd1 vccd1 vccd1 _10526_/A sky130_fd_sc_hd__buf_6
XFILLER_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06073_ _05702_/A _08209_/A _05818_/A _08082_/A vssd1 vssd1 vccd1 vccd1 _06073_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_144_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ _09901_/A _09901_/B vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__nor2_1
XFILLER_99_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08217__B1_N _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09832_ _09647_/A _09971_/A _09834_/A _09761_/C vssd1 vssd1 vccd1 vccd1 _09837_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _09908_/A _09947_/B _09763_/C vssd1 vssd1 vccd1 vccd1 _09842_/A sky130_fd_sc_hd__and3_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06975_ _07086_/B vssd1 vssd1 vccd1 vccd1 _07563_/A sky130_fd_sc_hd__buf_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08714_ _10805_/Q _08744_/B vssd1 vssd1 vccd1 vccd1 _08740_/A sky130_fd_sc_hd__xor2_1
X_05926_ _05885_/A _05888_/B _05889_/X _05692_/A _05925_/X vssd1 vssd1 vccd1 vccd1
+ _05926_/X sky130_fd_sc_hd__a221o_1
X_09694_ _09904_/A _09828_/B _09647_/A _09693_/Y vssd1 vssd1 vccd1 vccd1 _09710_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _10796_/Q _08638_/X _10192_/A vssd1 vssd1 vccd1 vccd1 _08646_/B sky130_fd_sc_hd__o21ai_1
X_05857_ _08268_/A _05857_/B vssd1 vssd1 vccd1 vccd1 _05858_/A sky130_fd_sc_hd__and2_1
XFILLER_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08576_ _10778_/Q _08576_/B vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__xor2_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05788_ _05788_/A _05788_/B _05788_/C _05802_/A vssd1 vssd1 vccd1 vccd1 _05788_/X
+ sky130_fd_sc_hd__or4_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10058__A1 _10487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07527_ _07648_/B _07527_/B _07643_/A vssd1 vssd1 vccd1 vccd1 _07638_/B sky130_fd_sc_hd__or3b_1
XFILLER_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07458_ _07493_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07460_/A sky130_fd_sc_hd__xor2_1
XFILLER_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06409_ _06626_/A _06409_/B _06409_/C vssd1 vssd1 vccd1 vccd1 _06717_/A sky130_fd_sc_hd__and3_1
XFILLER_148_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07389_ _07728_/A vssd1 vssd1 vccd1 vccd1 _07592_/A sky130_fd_sc_hd__buf_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09128_ _07974_/A _09123_/X _09125_/X _09127_/X vssd1 vssd1 vccd1 vccd1 _09128_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09059_ _10057_/A vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input11_A io_wbs_m2s_addr[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09439__B1 _10351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10805_ _10821_/CLK _10805_/D vssd1 vssd1 vccd1 vccd1 _10805_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10736_ _10751_/CLK _10736_/D vssd1 vssd1 vccd1 vccd1 _10736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08662__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08662__B2 _10799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05476__B2 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10667_ _10671_/CLK _10667_/D vssd1 vssd1 vccd1 vccd1 _10667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10598_ _10968_/CLK _10598_/D vssd1 vssd1 vccd1 vccd1 _10598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_115_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10221__B2 _10043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06760_ _06779_/A _06779_/B vssd1 vssd1 vccd1 vccd1 _06762_/A sky130_fd_sc_hd__and2b_1
XFILLER_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05951__A2 _05788_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05711_ _08146_/A vssd1 vssd1 vccd1 vccd1 _05711_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06691_ _06691_/A _06691_/B vssd1 vssd1 vccd1 vccd1 _06693_/A sky130_fd_sc_hd__nand2_1
XFILLER_91_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08430_ _10774_/Q _10773_/Q _08559_/B vssd1 vssd1 vccd1 vccd1 _08565_/C sky130_fd_sc_hd__and3_1
XFILLER_52_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05642_ _10680_/Q vssd1 vssd1 vccd1 vccd1 _05913_/A sky130_fd_sc_hd__inv_2
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08361_ _10679_/Q _08044_/A _08359_/Y _08360_/X vssd1 vssd1 vccd1 vccd1 _08363_/A
+ sky130_fd_sc_hd__a211o_1
X_05573_ _08339_/B vssd1 vssd1 vccd1 vccd1 _08332_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__08102__B1 _05728_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ _07312_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07313_/B sky130_fd_sc_hd__and2_1
XFILLER_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ input31/X _08212_/X _08052_/A _08287_/A _08175_/A vssd1 vssd1 vccd1 vccd1
+ _08293_/B sky130_fd_sc_hd__o221a_1
X_07243_ _07246_/A _07246_/B vssd1 vssd1 vccd1 vccd1 _07269_/A sky130_fd_sc_hd__nand2_1
XFILLER_20_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07174_ _07193_/A _07175_/B vssd1 vssd1 vccd1 vccd1 _07176_/A sky130_fd_sc_hd__or2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06125_ input8/X vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__buf_2
XFILLER_127_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06056_ _08318_/A vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__clkinv_2
XFILLER_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input3_A io_qei_ch_b vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _09815_/A _09815_/B vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__xor2_2
XFILLER_87_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09749_/A sky130_fd_sc_hd__xnor2_1
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06958_ _07641_/A _07645_/A _07644_/B vssd1 vssd1 vccd1 vccd1 _07635_/B sky130_fd_sc_hd__nand3_1
XFILLER_55_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05909_ _05909_/A _05909_/B vssd1 vssd1 vccd1 vccd1 _05909_/Y sky130_fd_sc_hd__xnor2_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09811_/B _09677_/B _09676_/X vssd1 vssd1 vccd1 vccd1 _09923_/B sky130_fd_sc_hd__or3b_1
XFILLER_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06889_ _06886_/A _06886_/B _06891_/A _06891_/B vssd1 vssd1 vccd1 vccd1 _06890_/B
+ sky130_fd_sc_hd__a2bb2oi_2
XANTENNA__08341__B1 _05570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05912__B _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _10792_/Q _10791_/Q _08628_/C vssd1 vssd1 vccd1 vccd1 _08642_/D sky130_fd_sc_hd__and3_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08559_ _10773_/Q _08559_/B vssd1 vssd1 vccd1 vccd1 _08559_/X sky130_fd_sc_hd__and2_1
XFILLER_161_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10521_ _06124_/X _10522_/A _10520_/X _05983_/X vssd1 vssd1 vccd1 vccd1 _10979_/D
+ sky130_fd_sc_hd__a211o_2
XANTENNA__10451__A1 _06163_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10452_ _10954_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__or2_1
XFILLER_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08016__A _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10383_ _10934_/Q _10405_/B vssd1 vssd1 vccd1 vccd1 _10383_/X sky130_fd_sc_hd__and2_1
XFILLER_124_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08686__A _08686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09281__S _09296_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06918__B _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09310__A _09313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10719_ _10935_/CLK _10719_/D vssd1 vssd1 vccd1 vccd1 _10719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09060__A1 _10935_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07930_ input8/X vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__inv_2
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07861_ _07848_/X _05460_/D _07844_/X _07860_/Y vssd1 vssd1 vccd1 vccd1 _10628_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_69_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09600_ _09600_/A _09653_/A vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__or2_1
XFILLER_110_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06812_ _06805_/A _06805_/B _06293_/A vssd1 vssd1 vccd1 vccd1 _06813_/B sky130_fd_sc_hd__a21oi_1
XFILLER_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07792_ _07792_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__xnor2_1
X_09531_ _10871_/Q _09408_/X _09529_/Y _09530_/X vssd1 vssd1 vccd1 vccd1 _10871_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06743_ _06752_/B _06743_/B vssd1 vssd1 vccd1 vccd1 _06774_/B sky130_fd_sc_hd__xnor2_2
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09462_ _09462_/A _09462_/B _09462_/C vssd1 vssd1 vccd1 vccd1 _09501_/A sky130_fd_sc_hd__and3_1
XFILLER_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06674_ _06674_/A _06681_/A _06674_/C vssd1 vssd1 vccd1 vccd1 _06678_/A sky130_fd_sc_hd__nand3_1
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05688__A1 _05570_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08413_ _10495_/A vssd1 vssd1 vccd1 vccd1 _10394_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05625_ _10549_/Q _05630_/A _10550_/Q vssd1 vssd1 vccd1 vccd1 _05626_/B sky130_fd_sc_hd__o21ai_1
X_09393_ _09430_/A _09393_/B vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10069__C _10140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08344_ _08263_/X _08350_/B _08340_/Y _08343_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08344_/X sky130_fd_sc_hd__o311a_1
X_05556_ _10559_/Q _10558_/Q _05610_/A vssd1 vssd1 vccd1 vccd1 _05604_/A sky130_fd_sc_hd__or3_1
XFILLER_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06844__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08275_ _08277_/A vssd1 vssd1 vccd1 vccd1 _08278_/A sky130_fd_sc_hd__buf_2
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05487_ _05487_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05487_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10366__A _10495_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07226_ _07235_/C _07142_/B _07224_/X _07223_/X _07217_/Y vssd1 vssd1 vccd1 vccd1
+ _07227_/B sky130_fd_sc_hd__a311o_1
XFILLER_20_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_41_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10640_/CLK sky130_fd_sc_hd__clkbuf_16
X_07157_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07282_/A sky130_fd_sc_hd__xor2_1
XFILLER_3_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06108_ _10704_/Q _08297_/B vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__or2_1
XFILLER_133_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07675__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07088_ _07089_/A _07089_/B vssd1 vssd1 vccd1 vccd1 _07359_/A sky130_fd_sc_hd__and2_1
XFILLER_161_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06039_ _06039_/A vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05915__A2 _05912_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _09647_/A _09647_/B _09728_/X vssd1 vssd1 vccd1 vccd1 _09730_/B sky130_fd_sc_hd__a21oi_2
XFILLER_43_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10504_ _10504_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10504_/X sky130_fd_sc_hd__or2_1
XFILLER_156_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10435_ _06124_/X _10431_/X _10434_/X _08563_/X vssd1 vssd1 vccd1 vccd1 _10947_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10188__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09042__A1 _07732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_7_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 _10709_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10366_ _10495_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10427_/B sky130_fd_sc_hd__nand2_1
XFILLER_98_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10297_ _10297_/A vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__inv_2
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05833__A _10675_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05410_ _05408_/Y hold10/A _05480_/A _08994_/A vssd1 vssd1 vccd1 vccd1 _05410_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06390_ _06502_/C vssd1 vssd1 vccd1 vccd1 _06489_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_159_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05341_ _10638_/Q vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08060_ _08352_/B vssd1 vssd1 vccd1 vccd1 _08061_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_135_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05272_ _10657_/Q vssd1 vssd1 vccd1 vccd1 _06039_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07011_ _07567_/A _07433_/A vssd1 vssd1 vccd1 vccd1 _07472_/A sky130_fd_sc_hd__and2_1
XFILLER_161_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08962_ _10947_/Q _10430_/B _08961_/X vssd1 vssd1 vccd1 vccd1 _08962_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_88_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07913_ _07916_/A _07913_/B vssd1 vssd1 vccd1 vccd1 _10642_/D sky130_fd_sc_hd__nor2_1
XANTENNA__09573__A_N _09567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08893_ _08889_/X _08890_/X _08891_/X _08892_/Y _08670_/A vssd1 vssd1 vccd1 vccd1
+ _08893_/X sky130_fd_sc_hd__o311a_1
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07844_ _08557_/A vssd1 vssd1 vccd1 vccd1 _07844_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07775_ _07773_/Y _07773_/B _07775_/S vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _09514_/A _09514_/B _09514_/C vssd1 vssd1 vccd1 vccd1 _09516_/B sky130_fd_sc_hd__nand3_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06726_ _07796_/A _06726_/B vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__or2_1
XFILLER_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09445_ _09676_/B _09445_/B vssd1 vssd1 vccd1 vccd1 _09448_/A sky130_fd_sc_hd__xor2_4
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06657_ _06657_/A _06657_/B vssd1 vssd1 vccd1 vccd1 _06658_/B sky130_fd_sc_hd__nor2_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05608_ _10696_/Q vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__clkbuf_2
X_09376_ _09376_/A vssd1 vssd1 vccd1 vccd1 _10065_/B sky130_fd_sc_hd__inv_2
XFILLER_40_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06588_ _06576_/B _06587_/C _06587_/B vssd1 vssd1 vccd1 vccd1 _06589_/B sky130_fd_sc_hd__a21oi_1
XFILLER_71_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10406__A1 _06178_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ _08327_/A _08327_/B vssd1 vssd1 vccd1 vccd1 _08339_/C sky130_fd_sc_hd__and2_1
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05539_ _10541_/Q vssd1 vssd1 vccd1 vccd1 _05539_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10096__A _10097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06086__B2 _06066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ _08258_/A vssd1 vssd1 vccd1 vccd1 _08258_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07209_ _07280_/C _07209_/B vssd1 vssd1 vccd1 vccd1 _07279_/B sky130_fd_sc_hd__or2_1
XFILLER_106_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09024__A1 _10198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08189_ _08191_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08189_/X sky130_fd_sc_hd__or2_1
X_10220_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10220_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10151_ _10151_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _10126_/A _10082_/B vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__and2_1
XFILLER_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10342__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06749__A _06769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08838__A1 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ _10984_/CLK _10984_/D vssd1 vssd1 vccd1 vccd1 _10984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05521__B1 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10418_ _10943_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10418_/X sky130_fd_sc_hd__and2_1
XFILLER_125_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _09312_/X _06371_/C _10346_/X _10918_/Q vssd1 vssd1 vccd1 vccd1 _10918_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_140_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07329__A1 _07562_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05890_ _10658_/Q _05895_/A vssd1 vssd1 vccd1 vccd1 _05891_/B sky130_fd_sc_hd__nand2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07560_ _07560_/A vssd1 vssd1 vccd1 vccd1 _07729_/A sky130_fd_sc_hd__buf_2
XFILLER_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06511_ _06511_/A _06511_/B vssd1 vssd1 vccd1 vccd1 _06512_/B sky130_fd_sc_hd__nand2_1
XFILLER_62_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07491_ _07509_/A _07509_/B vssd1 vssd1 vccd1 vccd1 _07510_/A sky130_fd_sc_hd__nor2_1
XFILLER_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09230_ _10441_/A vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06442_ _06442_/A _06442_/B vssd1 vssd1 vccd1 vccd1 _06469_/B sky130_fd_sc_hd__nand2_1
XFILLER_142_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ _10810_/Q _08985_/X _08988_/X _10723_/Q _09160_/X vssd1 vssd1 vccd1 vccd1
+ _09161_/X sky130_fd_sc_hd__a221o_1
X_06373_ _06305_/A _06274_/B _06262_/A vssd1 vssd1 vccd1 vccd1 _06374_/A sky130_fd_sc_hd__o21ai_2
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08112_ _08112_/A vssd1 vssd1 vccd1 vccd1 _10685_/D sky130_fd_sc_hd__clkbuf_1
X_05324_ _05827_/A _05324_/B vssd1 vssd1 vccd1 vccd1 _05324_/X sky130_fd_sc_hd__and2_1
XANTENNA__06068__B2 _06066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ _09092_/A _09098_/B vssd1 vssd1 vccd1 vccd1 _09118_/A sky130_fd_sc_hd__or2_1
XFILLER_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05815__A1 _05405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08043_ _08043_/A vssd1 vssd1 vccd1 vccd1 _08044_/A sky130_fd_sc_hd__buf_2
XFILLER_135_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08114__A _08263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09994_ _10123_/A vssd1 vssd1 vccd1 vccd1 _10489_/A sky130_fd_sc_hd__inv_2
XANTENNA__09309__A2 _09310_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08945_ _09124_/C _09142_/D vssd1 vssd1 vccd1 vccd1 _08968_/A sky130_fd_sc_hd__or2_1
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08876_ _08876_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _08876_/Y sky130_fd_sc_hd__nor2_1
XFILLER_97_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07827_ _07848_/A vssd1 vssd1 vccd1 vccd1 _07827_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06288__B _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07758_ _07758_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _10117_/A sky130_fd_sc_hd__xnor2_4
XFILLER_71_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06709_ _06717_/A _06717_/B vssd1 vssd1 vccd1 vccd1 _06711_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09599__B _09599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _07689_/A _09441_/A vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__or2b_1
XFILLER_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _09454_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09460_/B sky130_fd_sc_hd__xor2_1
XFILLER_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09359_ _09359_/A vssd1 vssd1 vccd1 vccd1 _09361_/A sky130_fd_sc_hd__inv_2
XFILLER_166_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06059__B2 _05877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10203_ _10949_/Q _10933_/Q vssd1 vssd1 vccd1 vccd1 _10203_/X sky130_fd_sc_hd__or2b_1
XFILLER_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08959__A _09736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input41_A io_wbs_m2s_data[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _10134_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__xnor2_1
XFILLER_48_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10065_ _09924_/B _10065_/B _10065_/C _10065_/D vssd1 vssd1 vccd1 vccd1 _10131_/C
+ sky130_fd_sc_hd__and4b_1
XFILLER_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_54_clock_A _10682_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10967_ _10967_/CLK _10967_/D vssd1 vssd1 vccd1 vccd1 _10967_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10898_ _10926_/CLK _10898_/D vssd1 vssd1 vccd1 vccd1 _10898_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_15_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06222__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07773__A _10508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06991_ _07166_/A vssd1 vssd1 vccd1 vccd1 _07021_/A sky130_fd_sc_hd__clkbuf_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08730_ _06163_/X _08728_/X _08729_/X _10805_/Q vssd1 vssd1 vccd1 vccd1 _08730_/X
+ sky130_fd_sc_hd__a22o_1
X_05942_ _05838_/B _05941_/Y _05803_/A vssd1 vssd1 vccd1 vccd1 _05942_/X sky130_fd_sc_hd__a21o_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08661_ _08661_/A _08671_/A vssd1 vssd1 vccd1 vccd1 _08820_/A sky130_fd_sc_hd__or2_2
XFILLER_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05873_ _10660_/Q vssd1 vssd1 vccd1 vccd1 _05883_/A sky130_fd_sc_hd__buf_2
X_07612_ _07539_/A _07505_/A _07505_/B _07536_/X _07611_/Y vssd1 vssd1 vccd1 vccd1
+ _07613_/A sky130_fd_sc_hd__a41o_1
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08592_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ _07543_/A _07753_/A vssd1 vssd1 vccd1 vccd1 _07544_/B sky130_fd_sc_hd__nor2_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07474_ _07747_/B _07474_/B vssd1 vssd1 vccd1 vccd1 _07475_/C sky130_fd_sc_hd__nand2_1
XFILLER_61_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08109__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09213_ _09250_/A vssd1 vssd1 vccd1 vccd1 _09296_/S sky130_fd_sc_hd__buf_2
XANTENNA__07013__A _07013_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06425_ _06425_/A _06425_/B vssd1 vssd1 vccd1 vccd1 _06425_/Y sky130_fd_sc_hd__nor2_1
XFILLER_148_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09144_ _10957_/Q _09164_/B vssd1 vssd1 vccd1 vccd1 _09144_/Y sky130_fd_sc_hd__nor2_1
X_06356_ _10978_/Q _06554_/B _06554_/C vssd1 vssd1 vccd1 vccd1 _06451_/C sky130_fd_sc_hd__and3_1
XFILLER_148_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05307_ _10669_/Q _05347_/B vssd1 vssd1 vccd1 vccd1 _05854_/A sky130_fd_sc_hd__or2_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09075_ _09179_/A vssd1 vssd1 vccd1 vccd1 _09297_/S sky130_fd_sc_hd__clkbuf_4
X_06287_ _06287_/A _06287_/B vssd1 vssd1 vccd1 vccd1 _06371_/C sky130_fd_sc_hd__nor2_2
XFILLER_163_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08026_ input35/X _08015_/X _08025_/X _08019_/X vssd1 vssd1 vccd1 vccd1 _10675_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_107_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09882__B _09882_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ _09977_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _10095_/A sky130_fd_sc_hd__nand2_1
XFILLER_104_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07961__A1 _06050_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ hold11/A _08928_/B vssd1 vssd1 vccd1 vccd1 _08928_/X sky130_fd_sc_hd__xor2_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_opt_5_0_clock_A _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08859_ _08845_/Y _08870_/B _08858_/X vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__a21o_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _10821_/CLK _10821_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10752_ _10784_/CLK _10752_/D vssd1 vssd1 vccd1 vccd1 _10752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08019__A _08563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10683_ _10987_/CLK _10683_/D vssd1 vssd1 vccd1 vccd1 _10683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10117_ _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__xor2_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10048_ _09980_/A _09980_/B _09975_/A vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06002__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06210_ _09104_/B vssd1 vssd1 vccd1 vccd1 _09148_/A sky130_fd_sc_hd__clkbuf_2
X_07190_ _07190_/A _07190_/B vssd1 vssd1 vccd1 vccd1 _07277_/A sky130_fd_sc_hd__or2_1
XFILLER_118_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06141_ _06008_/X _06131_/X _06140_/Y _06137_/X vssd1 vssd1 vccd1 vccd1 _10585_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06072_ _10658_/Q vssd1 vssd1 vccd1 vccd1 _07979_/A sky130_fd_sc_hd__buf_2
XFILLER_144_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09900_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09915_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08599__A _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09831_ _09908_/A _09828_/B _09830_/X vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__a21o_1
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09971_/A _09762_/B vssd1 vssd1 vccd1 vccd1 _09763_/C sky130_fd_sc_hd__xor2_1
X_06974_ _10983_/Q vssd1 vssd1 vccd1 vccd1 _07086_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08732_/B vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__07008__A _07008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05925_ _05892_/X _05924_/X _05889_/X _08169_/A vssd1 vssd1 vccd1 vccd1 _05925_/X
+ sky130_fd_sc_hd__o22a_1
X_09693_ _09904_/A _09947_/B _09828_/B _10057_/A vssd1 vssd1 vccd1 vccd1 _09693_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08644_ _10283_/A vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__buf_4
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05856_ _10669_/Q vssd1 vssd1 vccd1 vccd1 _08268_/A sky130_fd_sc_hd__buf_2
XFILLER_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08575_ _08575_/A vssd1 vssd1 vccd1 vccd1 _10777_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05787_ _05787_/A _05787_/B vssd1 vssd1 vccd1 vccd1 _05802_/A sky130_fd_sc_hd__nand2_2
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10369__A _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07526_ _07526_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__xor2_4
XFILLER_81_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07457_ _07394_/X _07327_/X _07378_/Y vssd1 vssd1 vccd1 vccd1 _07493_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07678__A _07678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ _06626_/A _06408_/B _06408_/C vssd1 vssd1 vccd1 vccd1 _06645_/A sky130_fd_sc_hd__and3_1
X_07388_ _07456_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07454_/C sky130_fd_sc_hd__nor2_1
XFILLER_148_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09127_ _09270_/A vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__buf_2
XFILLER_136_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06339_ _06575_/B vssd1 vssd1 vccd1 vccd1 _06459_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_109_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09058_ _09834_/B vssd1 vssd1 vccd1 vccd1 _10057_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09893__A _09893_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08009_ _08009_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08009_/Y sky130_fd_sc_hd__nand2_1
XFILLER_123_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ _10804_/CLK _10804_/D vssd1 vssd1 vccd1 vccd1 _10804_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10735_ _10751_/CLK _10735_/D vssd1 vssd1 vccd1 vccd1 _10735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05476__A2 _05471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10666_ _10666_/CLK _10666_/D vssd1 vssd1 vccd1 vccd1 _10666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10597_ _10914_/CLK _10597_/D vssd1 vssd1 vccd1 vccd1 _10597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output72_A _10858_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 _10865_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[31] sky130_fd_sc_hd__buf_2
XFILLER_122_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05710_ _08148_/A vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_64_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06690_ _06690_/A _06690_/B vssd1 vssd1 vccd1 vccd1 _06691_/B sky130_fd_sc_hd__or2_1
XANTENNA__09043__A _10966_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05641_ _05641_/A _05641_/B vssd1 vssd1 vccd1 vccd1 _05641_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_91_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08360_ _05528_/A _06011_/A _08037_/A _06115_/B _06024_/A vssd1 vssd1 vccd1 vccd1
+ _08360_/X sky130_fd_sc_hd__a41o_1
X_05572_ _10708_/Q vssd1 vssd1 vccd1 vccd1 _08339_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__08102__A1 _08098_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07311_ _07312_/A _07312_/B vssd1 vssd1 vccd1 vccd1 _07313_/A sky130_fd_sc_hd__nor2_1
X_08291_ _08263_/X _08296_/B _08287_/Y _08290_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08291_/X sky130_fd_sc_hd__o311a_1
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07242_ _07242_/A _07242_/B vssd1 vssd1 vccd1 vccd1 _07246_/B sky130_fd_sc_hd__xnor2_1
X_07173_ _07184_/A _07185_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07175_/B sky130_fd_sc_hd__o21bai_1
XFILLER_157_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06124_ _06124_/A vssd1 vssd1 vccd1 vccd1 _06124_/X sky130_fd_sc_hd__buf_2
XFILLER_133_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06055_ _08173_/A _07981_/A _06050_/X _09104_/A _06054_/X vssd1 vssd1 vccd1 vccd1
+ _06071_/C sky130_fd_sc_hd__a221o_1
XFILLER_160_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09218__A _09218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_141_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09814_ _09825_/B _09814_/B vssd1 vssd1 vccd1 vccd1 _09815_/B sky130_fd_sc_hd__xnor2_2
XFILLER_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09745_ _10493_/A _09810_/A _09745_/C vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__and3_1
X_06957_ _07651_/A _07659_/A _07658_/B vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__nor3_1
XFILLER_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05908_ _05908_/A _05908_/B vssd1 vssd1 vccd1 vccd1 _05909_/B sky130_fd_sc_hd__nor2_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09676_/A _09676_/B _09676_/C _09676_/D vssd1 vssd1 vccd1 vccd1 _09676_/X
+ sky130_fd_sc_hd__and4_1
X_06888_ _06872_/A _07801_/A _06873_/B vssd1 vssd1 vccd1 vccd1 _06891_/B sky130_fd_sc_hd__o21a_2
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08341__A1 _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05839_ _05831_/B _05831_/C _05838_/Y vssd1 vssd1 vccd1 vccd1 _05839_/X sky130_fd_sc_hd__o21a_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08627_ _08627_/A vssd1 vssd1 vccd1 vccd1 _10791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08558_ _08558_/A vssd1 vssd1 vccd1 vccd1 _10772_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07509_ _07509_/A _07509_/B vssd1 vssd1 vccd1 vccd1 _07510_/B sky130_fd_sc_hd__and2_1
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08489_ _08489_/A vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__buf_4
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10520_ _10531_/B _09121_/X _07715_/C vssd1 vssd1 vccd1 vccd1 _10520_/X sky130_fd_sc_hd__o21a_1
XANTENNA__05458__A2 _09078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09400__B _09400_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ _06163_/X _10446_/X _10450_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10953_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08016__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10382_ _10427_/B vssd1 vssd1 vccd1 vccd1 _10405_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08868__C1 _08310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_3_3_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 _10840_/CLK sky130_fd_sc_hd__clkbuf_2
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10718_ _10751_/CLK _10718_/D vssd1 vssd1 vccd1 vccd1 _10718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08207__A _08208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10649_ _10651_/CLK _10649_/D vssd1 vssd1 vccd1 vccd1 _10649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ _06193_/A _07849_/X _07850_/X _07859_/Y _07853_/X vssd1 vssd1 vccd1 vccd1
+ _07860_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_96_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06811_ _06851_/A _06811_/B vssd1 vssd1 vccd1 vccd1 _06813_/A sky130_fd_sc_hd__nand2_1
XFILLER_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07791_ _07791_/A _07791_/B vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__xnor2_1
XFILLER_77_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _10043_/A vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06742_ _06804_/A _06752_/C vssd1 vssd1 vccd1 vccd1 _06743_/B sky130_fd_sc_hd__nand2_1
XFILLER_83_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _09430_/A _09430_/B _09460_/X vssd1 vssd1 vccd1 vccd1 _09462_/C sky130_fd_sc_hd__a21o_1
X_06673_ _06684_/A _06684_/B vssd1 vssd1 vccd1 vccd1 _06941_/B sky130_fd_sc_hd__nand2_1
XFILLER_52_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08412_ _10432_/B vssd1 vssd1 vccd1 vccd1 _10495_/A sky130_fd_sc_hd__clkbuf_4
X_05624_ _10689_/Q vssd1 vssd1 vccd1 vccd1 _08148_/A sky130_fd_sc_hd__clkbuf_2
X_09392_ _09451_/B _09392_/B vssd1 vssd1 vccd1 vccd1 _09393_/B sky130_fd_sc_hd__and2_1
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08343_ _08037_/A _08351_/B _08341_/Y _08342_/Y _08062_/A vssd1 vssd1 vccd1 vccd1
+ _08343_/X sky130_fd_sc_hd__a311o_1
XFILLER_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05555_ _10557_/Q _05612_/A vssd1 vssd1 vccd1 vccd1 _05610_/A sky130_fd_sc_hd__or2_1
XFILLER_20_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08274_ input30/X vssd1 vssd1 vccd1 vccd1 _08274_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05486_ _05910_/B _05470_/B _05495_/A _05455_/X _05485_/Y vssd1 vssd1 vccd1 vccd1
+ _10544_/D sky130_fd_sc_hd__a221o_1
XFILLER_137_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__A _08117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07225_ _07217_/Y _07223_/X _07224_/X _07142_/B _07186_/A vssd1 vssd1 vccd1 vccd1
+ _07225_/X sky130_fd_sc_hd__o2111a_1
XFILLER_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07156_ _07132_/A _07132_/B _07286_/A _07133_/A vssd1 vssd1 vccd1 vccd1 _07355_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_145_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06107_ _10703_/Q _10702_/Q _08278_/B vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__or3_1
XFILLER_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07087_ _07087_/A _07087_/B vssd1 vssd1 vccd1 vccd1 _07089_/B sky130_fd_sc_hd__nor2_1
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06038_ _06038_/A vssd1 vssd1 vccd1 vccd1 _06038_/X sky130_fd_sc_hd__buf_4
XFILLER_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07989_ _06195_/X _07987_/X _07988_/X _07977_/X vssd1 vssd1 vccd1 vccd1 _10661_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09728_ _09665_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09728_/X sky130_fd_sc_hd__and2b_1
XFILLER_74_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09659_ _09716_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _09713_/B sky130_fd_sc_hd__and2_1
XFILLER_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10503_ _06008_/X _10496_/X _10502_/X _10498_/X vssd1 vssd1 vccd1 vccd1 _10972_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10434_ _10947_/Q _10440_/B vssd1 vssd1 vccd1 vccd1 _10434_/X sky130_fd_sc_hd__or2_1
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10365_ _10408_/A vssd1 vssd1 vccd1 vccd1 _10365_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10958_/Q _10942_/Q vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__and2b_1
XFILLER_97_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09292__S _09297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10360__A1 _08491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05340_ _05340_/A _05340_/B vssd1 vssd1 vccd1 vccd1 _05340_/X sky130_fd_sc_hd__and2_1
XANTENNA__07816__B1 _06257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05271_ _10662_/Q vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__clkinv_2
XANTENNA__07292__B2 _07563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07010_ _07567_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07555_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07776__A _10515_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06252__C1 _06247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08961_ _08948_/X _08953_/X _10474_/B _10478_/A vssd1 vssd1 vccd1 vccd1 _08961_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07912_ _10610_/Q _07906_/X _07910_/X _07911_/Y vssd1 vssd1 vccd1 vccd1 _07913_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_08892_ _08890_/X _08891_/X _08889_/X vssd1 vssd1 vccd1 vccd1 _08892_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07843_ _07827_/X _05461_/D _07823_/X _07842_/Y vssd1 vssd1 vccd1 vccd1 _10624_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07774_ _07774_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07775_/S sky130_fd_sc_hd__nor2_1
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09513_ _09613_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09514_/C sky130_fd_sc_hd__nor2_1
XFILLER_25_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06725_ _06725_/A _06725_/B vssd1 vssd1 vccd1 vccd1 _06726_/B sky130_fd_sc_hd__and2_1
XFILLER_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06858__A1 _07780_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09445_/B sky130_fd_sc_hd__and2_1
X_06656_ _06656_/A _06656_/B vssd1 vssd1 vccd1 vccd1 _06660_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05607_ _10697_/Q vssd1 vssd1 vccd1 vccd1 _08224_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06587_ _06587_/A _06587_/B _06587_/C vssd1 vssd1 vccd1 vccd1 _06589_/A sky130_fd_sc_hd__and3_1
X_09375_ _10895_/Q _10911_/Q vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__and2b_1
X_08326_ _08025_/A _08058_/X _08325_/X vssd1 vssd1 vccd1 vccd1 _08326_/X sky130_fd_sc_hd__o21ba_1
XFILLER_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05538_ _10542_/Q vssd1 vssd1 vccd1 vccd1 _05741_/B sky130_fd_sc_hd__inv_2
XFILLER_32_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08257_ _08267_/B _08253_/X _08254_/Y _08256_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08257_/X sky130_fd_sc_hd__a311o_1
XANTENNA__06086__A2 _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05469_ _05472_/B vssd1 vssd1 vccd1 vccd1 _05470_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07208_ _07208_/A _07208_/B vssd1 vssd1 vccd1 vccd1 _07209_/B sky130_fd_sc_hd__and2_1
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08188_ _08188_/A vssd1 vssd1 vccd1 vccd1 _08191_/A sky130_fd_sc_hd__buf_2
XFILLER_118_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07139_ _07138_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _07139_/X sky130_fd_sc_hd__and2b_1
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10150_ _10478_/A _10068_/B _10070_/B _10074_/A vssd1 vssd1 vccd1 vccd1 _10151_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10081_ _10081_/A _10081_/B _10081_/C vssd1 vssd1 vccd1 vccd1 _10082_/B sky130_fd_sc_hd__or3_1
XFILLER_88_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09406__A _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08838__A2 _08785_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10983_ _10984_/CLK _10983_/D vssd1 vssd1 vccd1 vccd1 _10983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09141__A _09153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10287__A _10287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06077__A2 _08352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10417_ _10408_/X _10723_/Q _10414_/X _10416_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10942_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _09634_/A _06352_/A _10192_/X _10917_/Q vssd1 vssd1 vccd1 vccd1 _10917_/D
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06005__A _08483_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _10277_/X _10278_/Y _10279_/S vssd1 vssd1 vccd1 vccd1 _10279_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_40_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10643_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06510_ _06510_/A _06510_/B vssd1 vssd1 vccd1 vccd1 _06511_/B sky130_fd_sc_hd__or2_1
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07490_ _07490_/A _07490_/B vssd1 vssd1 vccd1 vccd1 _07509_/B sky130_fd_sc_hd__xnor2_1
XFILLER_55_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_06441_ _06461_/B _06441_/B _06547_/C _06567_/B vssd1 vssd1 vccd1 vccd1 _06442_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09160_ _07981_/A _09123_/X _09127_/X _09159_/X vssd1 vssd1 vccd1 vccd1 _09160_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06372_ _06804_/A _06387_/A vssd1 vssd1 vccd1 vccd1 _06375_/A sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_55_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10987_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08111_ _08111_/A _08111_/B vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__and2_1
X_05323_ _05830_/A _05831_/B _08342_/A vssd1 vssd1 vccd1 vccd1 _05324_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06068__A2 _07981_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ _07393_/Y _08965_/Y _09209_/B vssd1 vssd1 vccd1 vccd1 _09112_/A sky130_fd_sc_hd__a21oi_2
XFILLER_119_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08042_ _08062_/A _08352_/B vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__nor2_2
XANTENNA__05815__A2 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09993_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__xor2_2
XFILLER_135_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08944_ _08944_/A vssd1 vssd1 vccd1 vccd1 _09124_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08875_ _10823_/Q vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09190__A1 _08198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07826_ _06255_/X _05453_/A _07823_/X _07825_/Y vssd1 vssd1 vccd1 vccd1 _10620_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_45_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07757_ _07757_/A _07757_/B vssd1 vssd1 vccd1 vccd1 _07758_/B sky130_fd_sc_hd__xor2_4
XFILLER_38_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06708_ _06630_/A _06631_/A _06630_/B vssd1 vssd1 vccd1 vccd1 _06717_/B sky130_fd_sc_hd__o21ba_1
X_07688_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09427_ _09427_/A _09427_/B vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__xor2_2
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06639_ _06715_/A _06639_/B vssd1 vssd1 vccd1 vccd1 _06641_/C sky130_fd_sc_hd__and2_1
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09358_ _10886_/Q _10902_/Q vssd1 vssd1 vccd1 vccd1 _09359_/A sky130_fd_sc_hd__or2b_1
XFILLER_138_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08309_ _08305_/A _08315_/C _08308_/Y vssd1 vssd1 vccd1 vccd1 _08309_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06059__A2 _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09289_ _09289_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09290_/A sky130_fd_sc_hd__and2_4
XFILLER_119_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10202_ _10933_/Q _10949_/Q vssd1 vssd1 vccd1 vccd1 _10202_/X sky130_fd_sc_hd__or2b_1
XFILLER_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10133_ _10133_/A _10133_/B vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__xnor2_1
XFILLER_79_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input34_A io_wbs_m2s_data[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _10064_/A _10064_/B vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__xnor2_2
XFILLER_88_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09181__A1 _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10966_ _10967_/CLK _10966_/D vssd1 vssd1 vccd1 vccd1 _10966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10897_ _10909_/CLK _10897_/D vssd1 vssd1 vccd1 vccd1 _10897_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_145_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10480__A _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06990_ _07248_/A vssd1 vssd1 vccd1 vccd1 _07166_/A sky130_fd_sc_hd__buf_2
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05574__A _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05941_ _08318_/A _05941_/B vssd1 vssd1 vccd1 vccd1 _05941_/Y sky130_fd_sc_hd__nand2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09172__B2 _10724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08660_ _10369_/A _08971_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08671_/A sky130_fd_sc_hd__and3_1
X_05872_ _05872_/A _05872_/B vssd1 vssd1 vccd1 vccd1 _05872_/X sky130_fd_sc_hd__and2_1
XFILLER_94_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07611_ _07622_/A _07536_/X _07505_/X vssd1 vssd1 vccd1 vccd1 _07611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08591_ input51/X _10253_/A vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__or2_1
XFILLER_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07542_ _07402_/A _07402_/B _07405_/A vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__a21oi_1
X_07473_ _07473_/A _07473_/B vssd1 vssd1 vccd1 vccd1 _07477_/B sky130_fd_sc_hd__and2_1
XFILLER_22_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09212_ _09275_/A vssd1 vssd1 vccd1 vccd1 _09212_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06424_ _06426_/A _06441_/B _06489_/B _06540_/A vssd1 vssd1 vccd1 vccd1 _06425_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_167_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06355_ _06550_/C vssd1 vssd1 vccd1 vccd1 _06554_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09143_ _10432_/A _09143_/B vssd1 vssd1 vccd1 vccd1 _09143_/Y sky130_fd_sc_hd__nor2_2
XFILLER_148_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05306_ _10668_/Q _10667_/Q _05350_/B vssd1 vssd1 vccd1 vccd1 _05347_/B sky130_fd_sc_hd__or3_1
XFILLER_163_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09074_ _09067_/X _09073_/X _08992_/X vssd1 vssd1 vccd1 vccd1 _10839_/D sky130_fd_sc_hd__o21a_2
XFILLER_136_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06286_ _06270_/A _06276_/A _06284_/X _06272_/Y vssd1 vssd1 vccd1 vccd1 _06287_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_136_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08125__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08025_ _08025_/A _08027_/B vssd1 vssd1 vccd1 vccd1 _08025_/X sky130_fd_sc_hd__or2_1
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08199__C1 _08120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08738__A1 _10537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07964__A _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08738__B2 _10806_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07683__B _09313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09976_ _09977_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _09976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08927_ _08927_/A _08927_/B _08927_/C vssd1 vssd1 vccd1 vccd1 _08927_/X sky130_fd_sc_hd__or3_1
XFILLER_39_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10540__D _10540_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08858_ _10820_/Q _08847_/X _08919_/B vssd1 vssd1 vccd1 vccd1 _08858_/X sky130_fd_sc_hd__o21a_1
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07809_ _10866_/Q _07824_/B vssd1 vssd1 vccd1 vccd1 _07809_/Y sky130_fd_sc_hd__nand2_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08789_ _10813_/Q _08789_/B vssd1 vssd1 vccd1 vccd1 _08803_/C sky130_fd_sc_hd__xor2_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _10822_/CLK _10820_/D vssd1 vssd1 vccd1 vccd1 _10820_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10856__CLK _10856_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09403__B _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10751_ _10751_/CLK _10751_/D vssd1 vssd1 vccd1 vccd1 _10751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10682_ _10682_/CLK _10682_/D vssd1 vssd1 vccd1 vccd1 _10682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07874__A _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10536__A1 _07729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10116_ _10109_/A _10109_/B _09626_/A vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__o21ai_1
XFILLER_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_96_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10047_ _09970_/A _09970_/B _09983_/B _09982_/B _09982_/A vssd1 vssd1 vccd1 vccd1
+ _10051_/A sky130_fd_sc_hd__o32a_1
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09313__B _09313_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10949_ _10971_/CLK _10949_/D vssd1 vssd1 vccd1 vccd1 _10949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10348__A1_N _09634_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06140_ _06140_/A _06145_/B vssd1 vssd1 vccd1 vccd1 _06140_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10194__B _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06071_ _06071_/A _06071_/B _06071_/C _06071_/D vssd1 vssd1 vccd1 vccd1 _06071_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_144_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07784__A _10510_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10527__A1 _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08599__B _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09830_ _09977_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09830_/X sky130_fd_sc_hd__and2_1
XFILLER_141_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09761_ _09647_/A _09834_/A _09761_/C vssd1 vssd1 vccd1 vccd1 _09762_/B sky130_fd_sc_hd__and3b_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _07622_/A vssd1 vssd1 vccd1 vccd1 _07539_/A sky130_fd_sc_hd__buf_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08688_/X _08710_/Y _08711_/X vssd1 vssd1 vccd1 vccd1 _10804_/D sky130_fd_sc_hd__o21a_1
X_05924_ _10690_/Q _05892_/B _05895_/X _08146_/A _05923_/X vssd1 vssd1 vccd1 vccd1
+ _05924_/X sky130_fd_sc_hd__o221a_1
X_09692_ _09692_/A vssd1 vssd1 vccd1 vccd1 _09947_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08643_ _10796_/Q _08686_/A _08643_/C vssd1 vssd1 vccd1 vccd1 _08648_/B sky130_fd_sc_hd__and3_1
X_05855_ _08013_/A _05858_/B _05852_/B vssd1 vssd1 vccd1 vccd1 _05935_/B sky130_fd_sc_hd__o21a_1
XFILLER_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08574_ _08580_/B _08574_/B _08576_/B vssd1 vssd1 vccd1 vccd1 _08575_/A sky130_fd_sc_hd__and3_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05786_ _05768_/X _05770_/X _05786_/C _05786_/D vssd1 vssd1 vccd1 vccd1 _05787_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07024__A _07169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _07525_/A _07525_/B vssd1 vssd1 vccd1 vccd1 _07526_/B sky130_fd_sc_hd__nand2_1
XFILLER_168_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07959__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07456_ _07456_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07499_/A sky130_fd_sc_hd__xnor2_1
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06407_ _06630_/A _06407_/B vssd1 vssd1 vccd1 vccd1 _06408_/C sky130_fd_sc_hd__xor2_1
X_07387_ _07391_/A _07459_/B _07748_/B _07378_/Y _07397_/A vssd1 vssd1 vccd1 vccd1
+ _07456_/B sky130_fd_sc_hd__a41o_1
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09126_ _09126_/A _09211_/A vssd1 vssd1 vccd1 vccd1 _09270_/A sky130_fd_sc_hd__and2_2
X_06338_ _06338_/A vssd1 vssd1 vccd1 vccd1 _06575_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09057_ _10967_/Q vssd1 vssd1 vccd1 vccd1 _09834_/B sky130_fd_sc_hd__clkbuf_2
X_06269_ _10917_/Q _10900_/Q vssd1 vssd1 vccd1 vccd1 _06270_/B sky130_fd_sc_hd__or2_1
XFILLER_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08008_ _08256_/A vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__inv_2
XFILLER_117_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09959_ _09959_/A _09958_/A vssd1 vssd1 vccd1 vccd1 _09960_/B sky130_fd_sc_hd__or2b_1
XANTENNA__05945__A1 _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08895__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _10821_/CLK _10803_/D vssd1 vssd1 vccd1 vccd1 _10803_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10734_ _10751_/CLK _10734_/D vssd1 vssd1 vccd1 vccd1 _10734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10665_ _10665_/CLK _10665_/D vssd1 vssd1 vccd1 vccd1 _10665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10596_ _10652_/CLK _10596_/D vssd1 vssd1 vccd1 vccd1 _10596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10509__A1 _05958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput70 _10856_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[22] sky130_fd_sc_hd__buf_2
Xoutput81 _10837_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[3] sky130_fd_sc_hd__buf_2
XFILLER_95_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05852__A _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05640_ _05910_/B _10543_/Q vssd1 vssd1 vccd1 vccd1 _05641_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05571_ _10570_/Q _05576_/A vssd1 vssd1 vccd1 vccd1 _05571_/X sky130_fd_sc_hd__xor2_1
XFILLER_32_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07310_ _07310_/A _07310_/B vssd1 vssd1 vccd1 vccd1 _07312_/B sky130_fd_sc_hd__or2_1
XFILLER_32_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08290_ _08297_/B _08253_/X _08288_/Y _08289_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08290_/X sky130_fd_sc_hd__a311o_1
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07241_ _07250_/A _07217_/B _07218_/X vssd1 vssd1 vccd1 vccd1 _07242_/A sky130_fd_sc_hd__o21ai_1
XFILLER_164_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07172_ _07192_/B _07192_/A vssd1 vssd1 vccd1 vccd1 _07185_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09994__A _10123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06123_ input16/X vssd1 vssd1 vccd1 vccd1 _06124_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_145_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06054_ _05744_/Y _07998_/A _05883_/A _08181_/A _06053_/X vssd1 vssd1 vccd1 vccd1
+ _06054_/X sky130_fd_sc_hd__a221o_1
XFILLER_160_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09813_ _09743_/A _09743_/B _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09814_/B
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_143_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09744_ _09744_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09745_/C sky130_fd_sc_hd__nand2_1
XFILLER_74_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06956_ _07663_/A _07662_/B vssd1 vssd1 vccd1 vccd1 _07658_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05907_ _05907_/A vssd1 vssd1 vccd1 vccd1 _05908_/A sky130_fd_sc_hd__inv_2
XFILLER_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09675_ _09733_/B _09675_/B vssd1 vssd1 vccd1 vccd1 _09679_/A sky130_fd_sc_hd__nand2_2
X_06887_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _07801_/A sky130_fd_sc_hd__nand2_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _08631_/C _08649_/A _08626_/C vssd1 vssd1 vccd1 vccd1 _08627_/A sky130_fd_sc_hd__and3b_1
X_05838_ _08025_/A _05838_/B vssd1 vssd1 vccd1 vccd1 _05838_/Y sky130_fd_sc_hd__nand2_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08557_ _08557_/A _08557_/B _08557_/C vssd1 vssd1 vccd1 vccd1 _08558_/A sky130_fd_sc_hd__and3_1
X_05769_ _05769_/A vssd1 vssd1 vccd1 vccd1 _05769_/Y sky130_fd_sc_hd__inv_2
XFILLER_168_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07508_ _07508_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07628_/A sky130_fd_sc_hd__xnor2_2
X_08488_ _08488_/A vssd1 vssd1 vccd1 vccd1 _10745_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07439_ _07439_/A vssd1 vssd1 vccd1 vccd1 _07732_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10450_ _10953_/Q _10456_/B vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__or2_1
XFILLER_136_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ _10806_/Q _09168_/A _09112_/A _09103_/Y _09108_/X vssd1 vssd1 vccd1 vccd1
+ _09110_/B sky130_fd_sc_hd__a221o_1
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10381_ _10365_/X _10714_/Q _10379_/X _10380_/X _10373_/X vssd1 vssd1 vccd1 vccd1
+ _10933_/D sky130_fd_sc_hd__o221a_1
XFILLER_163_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08313__A _09154_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08032__B _08034_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09109__A1 _10806_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06040__B1 _07976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10717_ _10751_/CLK _10717_/D vssd1 vssd1 vccd1 vccd1 _10717_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09310__C _09310_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10648_ _10654_/CLK _10648_/D vssd1 vssd1 vccd1 vccd1 _10648_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06008__A _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10579_ _10858_/CLK _10579_/D vssd1 vssd1 vccd1 vccd1 _10579_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08020__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06810_ _10928_/Q _07570_/A vssd1 vssd1 vccd1 vccd1 _06811_/B sky130_fd_sc_hd__nand2_1
XFILLER_56_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07790_ _07790_/A _07790_/B vssd1 vssd1 vccd1 vccd1 _07791_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_45_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06741_ _06741_/A vssd1 vssd1 vccd1 vccd1 _06834_/A sky130_fd_sc_hd__inv_2
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09460_ _09429_/A _09460_/B vssd1 vssd1 vccd1 vccd1 _09460_/X sky130_fd_sc_hd__and2b_1
XFILLER_58_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06672_ _06672_/A _06672_/B vssd1 vssd1 vccd1 vccd1 _06684_/B sky130_fd_sc_hd__xor2_1
XFILLER_92_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08411_ _08419_/A hold8/X _08992_/A _08410_/X vssd1 vssd1 vccd1 vccd1 _10727_/D sky130_fd_sc_hd__o211a_1
X_05623_ _05623_/A _05623_/B vssd1 vssd1 vccd1 vccd1 _05623_/X sky130_fd_sc_hd__and2_1
X_09391_ _09451_/B _09392_/B vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__nor2_1
XFILLER_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08342_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08342_/Y sky130_fd_sc_hd__nor2_1
X_05554_ _10556_/Q _10555_/Q _05663_/A _05663_/B vssd1 vssd1 vccd1 vccd1 _05612_/A
+ sky130_fd_sc_hd__or4_1
X_08273_ _08273_/A vssd1 vssd1 vccd1 vccd1 _10701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05485_ _05485_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05485_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07224_ _10981_/Q _07235_/B vssd1 vssd1 vccd1 vccd1 _07224_/X sky130_fd_sc_hd__and2_1
X_07155_ _07285_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07286_/A sky130_fd_sc_hd__nor2_1
XFILLER_118_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06106_ _10701_/Q _08267_/B vssd1 vssd1 vccd1 vccd1 _08278_/B sky130_fd_sc_hd__or2_2
XFILLER_133_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07086_ _07326_/A _07086_/B _07188_/B _07178_/A vssd1 vssd1 vccd1 vccd1 _07087_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06037_ _06037_/A vssd1 vssd1 vccd1 vccd1 _08105_/A sky130_fd_sc_hd__clkinv_2
XFILLER_160_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07988_ _07988_/A _07988_/B vssd1 vssd1 vccd1 vccd1 _07988_/X sky130_fd_sc_hd__or2_1
XFILLER_86_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09727_ _09727_/A _09727_/B vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__xnor2_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06939_ _06939_/A _06939_/B vssd1 vssd1 vccd1 vccd1 _07630_/A sky130_fd_sc_hd__xor2_4
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09658_ _09760_/B vssd1 vssd1 vccd1 vccd1 _09977_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08609_ _08609_/A vssd1 vssd1 vccd1 vccd1 _10786_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09589_ _09639_/B _09536_/B _09486_/A _09588_/X vssd1 vssd1 vccd1 vccd1 _09590_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07212__A _07415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08027__B _08027_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ _10502_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10502_/X sky130_fd_sc_hd__or2_1
XFILLER_156_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10433_ _10472_/B vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10188__A2 _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08250__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10364_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10408_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10295_ _10942_/Q _10958_/Q vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__or2b_1
XFILLER_78_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08069__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05270_ _10678_/Q vssd1 vssd1 vccd1 vccd1 _08352_/A sky130_fd_sc_hd__buf_2
XANTENNA__09018__A0 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09569__A1 _09527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08960_ _10068_/A vssd1 vssd1 vccd1 vccd1 _10478_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09991__B _10140_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07911_ _07911_/A vssd1 vssd1 vccd1 vccd1 _07911_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_130_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08891_ _08891_/A _08891_/B vssd1 vssd1 vccd1 vccd1 _08891_/X sky130_fd_sc_hd__and2_1
XFILLER_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06004__A0 input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09741__A1 _10480_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09741__B2 _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07842_ _06175_/A _07828_/X _07829_/X _07841_/Y _07832_/X vssd1 vssd1 vccd1 vccd1
+ _07842_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_84_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07773_ _10508_/A _07773_/B vssd1 vssd1 vccd1 vccd1 _07773_/Y sky130_fd_sc_hd__nand2_1
X_09512_ _10069_/A _09692_/A _09761_/C _09736_/B vssd1 vssd1 vccd1 vccd1 _09513_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06724_ _06725_/A _06725_/B vssd1 vssd1 vccd1 vccd1 _07796_/A sky130_fd_sc_hd__nor2_1
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09443_ _10967_/Q _09443_/B vssd1 vssd1 vccd1 vccd1 _09534_/C sky130_fd_sc_hd__nand2_1
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06655_ _06800_/A _06408_/B _06428_/B _06845_/A vssd1 vssd1 vccd1 vccd1 _06656_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_13_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09257__A0 _08298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05606_ _10558_/Q _05610_/A vssd1 vssd1 vccd1 vccd1 _05606_/X sky130_fd_sc_hd__xor2_1
X_09374_ _09923_/A _09674_/B _09372_/X _09373_/Y vssd1 vssd1 vccd1 vccd1 _09922_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06586_ _06591_/A _06591_/B vssd1 vssd1 vccd1 vccd1 _06949_/B sky130_fd_sc_hd__nand2_1
X_08325_ _08332_/B _08058_/A _08324_/Y _08120_/X vssd1 vssd1 vccd1 vccd1 _08325_/X
+ sky130_fd_sc_hd__a31o_1
X_05537_ _10543_/Q vssd1 vssd1 vccd1 vccd1 _05737_/B sky130_fd_sc_hd__inv_2
XFILLER_138_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08256_ _08256_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05468_ _05453_/X _05459_/X _05460_/X _05462_/X _05467_/X vssd1 vssd1 vccd1 vccd1
+ _05472_/B sky130_fd_sc_hd__a2111oi_1
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07207_ _07208_/A _07208_/B vssd1 vssd1 vccd1 vccd1 _07280_/C sky130_fd_sc_hd__nor2_1
X_08187_ _08188_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08196_/B sky130_fd_sc_hd__nand2_1
X_05399_ _10651_/Q _10575_/Q vssd1 vssd1 vccd1 vccd1 _05400_/B sky130_fd_sc_hd__xnor2_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07138_ _07138_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _07147_/B sky130_fd_sc_hd__xnor2_1
XFILLER_145_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07069_ _07149_/C _07186_/B _07312_/A vssd1 vssd1 vccd1 vccd1 _07070_/B sky130_fd_sc_hd__and3_1
XFILLER_0_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10080_ _10081_/A _10081_/B _10081_/C vssd1 vssd1 vccd1 vccd1 _10126_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10982_ _10985_/CLK _10982_/D vssd1 vssd1 vccd1 vccd1 _10982_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08038__A _08038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07877__A _07880_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10416_ input18/X _10399_/X _10415_/X vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__08223__A1 _08157_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10347_ _09312_/X _06281_/B _10346_/X _10916_/Q vssd1 vssd1 vccd1 vccd1 _10916_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_112_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08501__A _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ _10265_/A _10268_/Y _10265_/B vssd1 vssd1 vccd1 vccd1 _10278_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06021__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10478__A _10478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06440_ _06440_/A vssd1 vssd1 vccd1 vccd1 _06567_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06371_ _06371_/A _06371_/B _06371_/C vssd1 vssd1 vccd1 vccd1 _06387_/A sky130_fd_sc_hd__or3_1
XFILLER_159_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08110_ _10533_/A _08086_/X _08109_/X _05728_/X _08166_/A vssd1 vssd1 vccd1 vccd1
+ _08111_/B sky130_fd_sc_hd__o221a_1
X_05322_ _10677_/Q vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_148_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09090_ _09090_/A vssd1 vssd1 vccd1 vccd1 _09228_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08041_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__buf_2
XFILLER_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09992_ _10480_/A _10141_/B vssd1 vssd1 vccd1 vccd1 _10130_/B sky130_fd_sc_hd__nand2_1
XFILLER_103_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ _10518_/B vssd1 vssd1 vccd1 vccd1 _08943_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05984__C1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08874_ _10823_/Q _08888_/B vssd1 vssd1 vccd1 vccd1 _08883_/A sky130_fd_sc_hd__and2_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07825_ _06156_/A _06258_/X _07807_/X _07824_/Y _07811_/X vssd1 vssd1 vccd1 vccd1
+ _07825_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_84_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09190__A2 _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07756_ _07756_/A _07756_/B vssd1 vssd1 vccd1 vccd1 _07757_/B sky130_fd_sc_hd__xnor2_2
XFILLER_37_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06707_ _06719_/B _07791_/A _06706_/X vssd1 vssd1 vccd1 vccd1 _06711_/A sky130_fd_sc_hd__o21a_1
X_07687_ _07687_/A _07687_/B vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09426_ _10963_/Q _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09427_/B sky130_fd_sc_hd__and3_1
XFILLER_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06638_ _06638_/A _06638_/B vssd1 vssd1 vccd1 vccd1 _06639_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09357_ _10903_/Q _10887_/Q vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__or2b_1
X_06569_ _06570_/A _06570_/B vssd1 vssd1 vccd1 vccd1 _06597_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08308_ _08305_/A _08315_/C _08092_/A vssd1 vssd1 vccd1 vccd1 _08308_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09288_ _10828_/Q _09274_/X _09275_/X _09287_/X _09270_/X vssd1 vssd1 vccd1 vccd1
+ _09289_/B sky130_fd_sc_hd__a32o_1
XFILLER_20_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08239_ input25/X _08212_/X _08124_/X _08233_/A _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08240_/B sky130_fd_sc_hd__o221a_1
XFILLER_153_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10201_ _07098_/A _10192_/X _10200_/X vssd1 vssd1 vccd1 vccd1 _10899_/D sky130_fd_sc_hd__a21o_1
XFILLER_107_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10132_ _10480_/A _10068_/B _10131_/X _10068_/A vssd1 vssd1 vccd1 vccd1 _10133_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10063_ _10065_/C _10063_/B vssd1 vssd1 vccd1 vccd1 _10064_/B sky130_fd_sc_hd__nand2_1
XFILLER_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09181__A2 _09226_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input27_A io_wbs_m2s_data[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10965_ _10985_/CLK _10965_/D vssd1 vssd1 vccd1 vccd1 _10965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10896_ _10909_/CLK _10896_/D vssd1 vssd1 vccd1 vccd1 _10896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06016__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05940_ _08315_/B _05940_/B vssd1 vssd1 vccd1 vccd1 _05940_/X sky130_fd_sc_hd__or2_1
XFILLER_140_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05871_ _05848_/B _05823_/A _06052_/A vssd1 vssd1 vccd1 vccd1 _05872_/B sky130_fd_sc_hd__o21ai_1
XFILLER_27_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07610_ _07610_/A _07706_/B vssd1 vssd1 vccd1 vccd1 _09969_/A sky130_fd_sc_hd__xnor2_2
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08590_ _09403_/B vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07541_ _07410_/A _07410_/B _07540_/X vssd1 vssd1 vccd1 vccd1 _07546_/B sky130_fd_sc_hd__o21a_1
XFILLER_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07472_ _07472_/A _07472_/B vssd1 vssd1 vccd1 vccd1 _07473_/B sky130_fd_sc_hd__or2_1
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09211_ _09211_/A _09211_/B vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__nor2_2
XFILLER_22_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10490__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06423_ _06426_/A _06627_/B _06540_/A _06441_/B vssd1 vssd1 vccd1 vccd1 _06425_/A
+ sky130_fd_sc_hd__a22oi_1
X_09142_ _09142_/A _09142_/B _09142_/C _09142_/D vssd1 vssd1 vccd1 vccd1 _09143_/B
+ sky130_fd_sc_hd__or4_1
X_06354_ _06352_/B _06352_/C _06352_/A vssd1 vssd1 vccd1 vccd1 _06550_/C sky130_fd_sc_hd__o21ai_1
XFILLER_136_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05305_ _05353_/A vssd1 vssd1 vccd1 vccd1 _05350_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09073_ _10123_/A _10474_/B _10495_/B _10510_/A _09072_/X vssd1 vssd1 vccd1 vccd1
+ _09073_/X sky130_fd_sc_hd__a221o_1
XFILLER_108_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06285_ _06284_/X _06272_/Y _06270_/A _06276_/A vssd1 vssd1 vccd1 vccd1 _06287_/A
+ sky130_fd_sc_hd__o211a_1
X_08024_ input34/X _08015_/X _08023_/Y _08019_/X vssd1 vssd1 vccd1 vccd1 _10674_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_150_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09975_ _09975_/A _09975_/B vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08926_ _09153_/A _08926_/B vssd1 vssd1 vccd1 vccd1 _10829_/D sky130_fd_sc_hd__nor2_1
XFILLER_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08857_ _08866_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08870_/C sky130_fd_sc_hd__and2_1
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07808_ _07849_/A vssd1 vssd1 vccd1 vccd1 _07824_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08788_ _08783_/Y _08784_/X _08787_/X vssd1 vssd1 vccd1 vccd1 _10812_/D sky130_fd_sc_hd__o21a_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07739_ _07739_/A _07739_/B vssd1 vssd1 vccd1 vccd1 _07740_/B sky130_fd_sc_hd__xnor2_1
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10750_ _10776_/CLK _10750_/D vssd1 vssd1 vccd1 vccd1 _10750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09409_ _09409_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10481__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ _10684_/CLK _10681_/D vssd1 vssd1 vccd1 vccd1 _10681_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07937__A0 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08051__A _08124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10115_ _10115_/A vssd1 vssd1 vccd1 vccd1 _10115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_54_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10693_/CLK sky130_fd_sc_hd__clkbuf_16
X_10046_ _10046_/A _09985_/A vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__or2b_1
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_69_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10545_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10948_ _10971_/CLK _10948_/D vssd1 vssd1 vccd1 vccd1 _10948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10879_ _10879_/CLK _10879_/D vssd1 vssd1 vccd1 vccd1 _10879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06070_ _06070_/A _06070_/B vssd1 vssd1 vccd1 vccd1 _06071_/D sky130_fd_sc_hd__nand2_1
XFILLER_145_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10491__A _10491_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05585__A _08315_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09057__A _10967_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09760_ _09834_/B _09760_/B vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__and2_1
X_06972_ _07715_/D vssd1 vssd1 vccd1 vccd1 _07622_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _10533_/A _08694_/X _08695_/X _10804_/Q _08175_/X vssd1 vssd1 vccd1 vccd1
+ _08711_/X sky130_fd_sc_hd__o221a_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05923_ _06035_/A _05897_/X _05895_/X _08148_/A _05922_/X vssd1 vssd1 vccd1 vccd1
+ _05923_/X sky130_fd_sc_hd__a221o_1
X_09691_ _09761_/C vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08642_ _10795_/Q _10794_/Q _10793_/Q _08642_/D vssd1 vssd1 vccd1 vccd1 _08643_/C
+ sky130_fd_sc_hd__and4_1
X_05854_ _05854_/A _05854_/B vssd1 vssd1 vccd1 vccd1 _05858_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08573_ _08578_/C _08578_/D vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__nand2_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05785_ _05785_/A _05785_/B _05785_/C vssd1 vssd1 vccd1 vccd1 _05786_/D sky130_fd_sc_hd__and3_1
XFILLER_42_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07524_ _07649_/A vssd1 vssd1 vccd1 vccd1 _07527_/B sky130_fd_sc_hd__inv_2
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07455_ _07455_/A _07455_/B vssd1 vssd1 vccd1 vccd1 _07502_/A sky130_fd_sc_hd__nand2_2
XFILLER_50_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06406_ _06690_/A _06426_/A _06428_/B vssd1 vssd1 vccd1 vccd1 _06407_/B sky130_fd_sc_hd__and3b_1
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07386_ _07391_/A _07386_/B vssd1 vssd1 vccd1 vccd1 _07397_/A sky130_fd_sc_hd__nor2_2
XFILLER_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09125_ _05461_/D _09136_/A _09148_/A _06035_/A _08976_/A vssd1 vssd1 vccd1 vccd1
+ _09125_/X sky130_fd_sc_hd__a221o_1
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06337_ _06436_/A _06409_/B vssd1 vssd1 vccd1 vccd1 _06872_/A sky130_fd_sc_hd__and2_1
XFILLER_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ _07713_/A _08965_/Y _09036_/X _09052_/X _09055_/X vssd1 vssd1 vccd1 vccd1
+ _09056_/X sky130_fd_sc_hd__a221o_1
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06268_ _06558_/B _06360_/A _06267_/Y vssd1 vssd1 vccd1 vccd1 _06275_/A sky130_fd_sc_hd__o21ai_1
XFILLER_68_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08007_ input26/X _08002_/X _08005_/X _08006_/X vssd1 vssd1 vccd1 vccd1 _10667_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_135_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06199_ _10441_/A vssd1 vssd1 vccd1 vccd1 _07977_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07395__A1 _07393_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09958_ _09958_/A _09959_/A vssd1 vssd1 vccd1 vccd1 _09960_/A sky130_fd_sc_hd__or2b_1
XFILLER_89_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08909_ _08658_/X _08907_/Y _08908_/X vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__a21oi_1
XFILLER_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _09890_/B _09889_/B vssd1 vssd1 vccd1 vccd1 _09961_/B sky130_fd_sc_hd__and2b_1
XFILLER_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _10804_/CLK _10802_/D vssd1 vssd1 vccd1 vccd1 _10802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ _10751_/CLK _10733_/D vssd1 vssd1 vccd1 vccd1 _10733_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__07869__B _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10664_ _10665_/CLK _10664_/D vssd1 vssd1 vccd1 vccd1 _10664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10595_ _10653_/CLK _10595_/D vssd1 vssd1 vccd1 vccd1 _10595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_127_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput60 _10847_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[13] sky130_fd_sc_hd__buf_2
Xoutput71 _10857_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[23] sky130_fd_sc_hd__buf_2
Xoutput82 _10838_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[4] sky130_fd_sc_hd__buf_2
XFILLER_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08335__B1 _08092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10029_ _10029_/A _10029_/B vssd1 vssd1 vccd1 vccd1 _10105_/B sky130_fd_sc_hd__xor2_2
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05570_ _08339_/A vssd1 vssd1 vccd1 vccd1 _05570_/X sky130_fd_sc_hd__buf_2
XFILLER_91_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07240_ _07235_/C _07235_/B _07515_/A _07239_/Y vssd1 vssd1 vccd1 vccd1 _07246_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_149_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07171_ _07196_/A _07184_/B _07170_/X vssd1 vssd1 vccd1 vccd1 _07192_/A sky130_fd_sc_hd__o21a_1
XFILLER_158_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_41_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06122_ _06122_/A vssd1 vssd1 vccd1 vccd1 _10583_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06053_ _10701_/Q _08268_/A vssd1 vssd1 vccd1 vccd1 _06053_/X sky130_fd_sc_hd__xor2_1
XFILLER_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09812_ _09812_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09825_/B sky130_fd_sc_hd__xnor2_2
XFILLER_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09743_ _09743_/A _09743_/B vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__xor2_1
X_06955_ _07671_/A _07670_/B vssd1 vssd1 vccd1 vccd1 _07662_/B sky130_fd_sc_hd__nor2_1
XFILLER_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07129__A1 _10985_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05906_ _05906_/A _05906_/B vssd1 vssd1 vccd1 vccd1 _05906_/X sky130_fd_sc_hd__and2_1
XFILLER_28_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09674_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09675_/B sky130_fd_sc_hd__nand2_1
X_06886_ _06886_/A _06886_/B vssd1 vssd1 vccd1 vccd1 _06891_/A sky130_fd_sc_hd__xor2_4
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _08600_/X _08628_/C _10791_/Q vssd1 vssd1 vccd1 vccd1 _08626_/C sky130_fd_sc_hd__a21o_1
X_05837_ _08327_/A vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__buf_2
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _10771_/Q _08547_/B _10772_/Q vssd1 vssd1 vccd1 vccd1 _08557_/C sky130_fd_sc_hd__a21o_1
X_05768_ _05766_/Y _10569_/Q _10568_/Q _05767_/Y vssd1 vssd1 vccd1 vccd1 _05768_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09250__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _07534_/C _07507_/B vssd1 vssd1 vccd1 vccd1 _07623_/A sky130_fd_sc_hd__nor2_2
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08487_ _08935_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__and2_1
XFILLER_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05699_ _05896_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__inv_2
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07438_ _07570_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _07726_/B sky130_fd_sc_hd__xnor2_2
XFILLER_168_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07369_ _07369_/A _07369_/B _07462_/A vssd1 vssd1 vccd1 vccd1 _07370_/B sky130_fd_sc_hd__nor3_1
XANTENNA__09054__A1 _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09108_ _08974_/A _09106_/X _09107_/Y _09079_/A _10719_/Q vssd1 vssd1 vccd1 vccd1
+ _09108_/X sky130_fd_sc_hd__a32o_1
X_10380_ _10526_/A _10371_/X _10376_/X vssd1 vssd1 vccd1 vccd1 _10380_/X sky130_fd_sc_hd__a21bo_1
XFILLER_109_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _05455_/X _09020_/B _06129_/B _05733_/X _09263_/A vssd1 vssd1 vccd1 vccd1
+ _09039_/X sky130_fd_sc_hd__o221a_1
XFILLER_123_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06114__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05953__A _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08868__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _10940_/CLK _10716_/D vssd1 vssd1 vccd1 vccd1 _10716_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10647_ _10865_/CLK _10647_/D vssd1 vssd1 vccd1 vccd1 _10647_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10578_ _10914_/CLK _10578_/D vssd1 vssd1 vccd1 vccd1 _10578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06024__A _06024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__B1 _09408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08308__B1 _08092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06740_ _06775_/A _07784_/B vssd1 vssd1 vccd1 vccd1 _06741_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06671_ _06671_/A _06671_/B vssd1 vssd1 vccd1 vccd1 _06684_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08410_ _08547_/A _10761_/Q vssd1 vssd1 vccd1 vccd1 _08410_/X sky130_fd_sc_hd__or2_1
XFILLER_18_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05622_ _10551_/Q _05626_/A vssd1 vssd1 vccd1 vccd1 _05623_/B sky130_fd_sc_hd__nand2_1
X_09390_ _09390_/A _09390_/B vssd1 vssd1 vccd1 vccd1 _09392_/B sky130_fd_sc_hd__xnor2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08341_ _08332_/A _08332_/B _05570_/X vssd1 vssd1 vccd1 vccd1 _08341_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05553_ _10553_/Q _10552_/Q _05623_/A vssd1 vssd1 vccd1 vccd1 _05663_/B sky130_fd_sc_hd__or3_1
XFILLER_149_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ _08270_/X _08272_/B vssd1 vssd1 vccd1 vccd1 _08273_/A sky130_fd_sc_hd__and2b_1
X_05484_ _05482_/X _05470_/B _05495_/A _09020_/A _05483_/Y vssd1 vssd1 vccd1 vccd1
+ _10543_/D sky130_fd_sc_hd__a221o_1
XFILLER_165_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07223_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07223_/X sky130_fd_sc_hd__and2_1
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07154_ _07296_/A _07309_/A _07309_/B _07153_/Y vssd1 vssd1 vccd1 vccd1 _07285_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_118_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06105_ _10700_/Q _06105_/B vssd1 vssd1 vccd1 vccd1 _08267_/B sky130_fd_sc_hd__or2_1
XANTENNA__08795__B1 _08780_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07085_ _07326_/A _07188_/B _07178_/A _07086_/B vssd1 vssd1 vccd1 vccd1 _07087_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06036_ _08115_/A _08119_/A _05405_/A _08059_/A _06035_/X vssd1 vssd1 vccd1 vccd1
+ _06036_/X sky130_fd_sc_hd__a221o_1
XFILLER_105_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10354__B1 _08494_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input1_A io_ba_match vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07987_ _08015_/A vssd1 vssd1 vccd1 vccd1 _07987_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09726_ _09787_/B _09726_/B vssd1 vssd1 vccd1 vccd1 _09727_/B sky130_fd_sc_hd__xnor2_2
X_06938_ _06938_/A _06938_/B vssd1 vssd1 vccd1 vccd1 _07625_/A sky130_fd_sc_hd__xnor2_4
XFILLER_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09657_ _09712_/A _09712_/B vssd1 vssd1 vccd1 vccd1 _09713_/A sky130_fd_sc_hd__xor2_1
X_06869_ _06869_/A _06869_/B vssd1 vssd1 vccd1 vccd1 _07761_/B sky130_fd_sc_hd__xnor2_2
XFILLER_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08611_/B _08649_/A _08608_/C vssd1 vssd1 vccd1 vccd1 _08609_/A sky130_fd_sc_hd__and3b_1
X_09588_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09588_/X sky130_fd_sc_hd__and2_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08539_ _08547_/A _10767_/Q _10768_/Q vssd1 vssd1 vccd1 vccd1 _08540_/C sky130_fd_sc_hd__a21o_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ _10515_/B vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10432_ _10432_/A _10432_/B _10432_/C vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__and3_2
XFILLER_171_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08324__A _08324_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ _08491_/X _07635_/A _09408_/X _10930_/Q vssd1 vssd1 vccd1 vccd1 _10930_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10294_ _07008_/A _10283_/X _10292_/X _10293_/X vssd1 vssd1 vccd1 vccd1 _10908_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_105_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10345__B1 _10184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06013__A1 _06008_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clock_A clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06019__A _06019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06252__A1 input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08529__B1 _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07910_ _07910_/A vssd1 vssd1 vccd1 vccd1 _07910_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_08890_ _10824_/Q _08876_/A _08928_/B vssd1 vssd1 vccd1 vccd1 _08890_/X sky130_fd_sc_hd__o21a_1
XFILLER_97_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07841_ _10874_/Q _07845_/B vssd1 vssd1 vccd1 vccd1 _07841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07772_ _10513_/A _07776_/B _06848_/B _06847_/A vssd1 vssd1 vccd1 vccd1 _07778_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09511_ _09599_/B vssd1 vssd1 vccd1 vccd1 _09761_/C sky130_fd_sc_hd__buf_2
X_06723_ _06638_/A _06638_/B _06721_/Y _06714_/B _06722_/Y vssd1 vssd1 vccd1 vccd1
+ _06725_/B sky130_fd_sc_hd__o32a_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09442_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__nand2_2
XFILLER_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06654_ _06654_/A _06654_/B vssd1 vssd1 vccd1 vccd1 _06700_/B sky130_fd_sc_hd__nor2_1
XFILLER_25_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05605_ _10698_/Q _05605_/B vssd1 vssd1 vccd1 vccd1 _05605_/X sky130_fd_sc_hd__or2_1
X_09373_ _09343_/A _09346_/A _09343_/B vssd1 vssd1 vccd1 vccd1 _09373_/Y sky130_fd_sc_hd__o21bai_1
X_06585_ _06585_/A _06585_/B vssd1 vssd1 vccd1 vccd1 _06591_/B sky130_fd_sc_hd__xnor2_1
XFILLER_40_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08324_ _08324_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05536_ _05818_/B _05536_/B vssd1 vssd1 vccd1 vccd1 _05652_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08255_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08342_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_137_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05467_ _05467_/A _05467_/B _05467_/C _05467_/D vssd1 vssd1 vccd1 vccd1 _05467_/X
+ sky130_fd_sc_hd__or4_4
XFILLER_119_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09009__B2 _10932_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07206_ _07301_/A _07302_/A _07205_/A vssd1 vssd1 vccd1 vccd1 _07208_/B sky130_fd_sc_hd__o21a_1
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08186_ _08186_/A vssd1 vssd1 vccd1 vccd1 _10692_/D sky130_fd_sc_hd__clkbuf_1
X_05398_ _05398_/A _05398_/B vssd1 vssd1 vccd1 vccd1 _05487_/A sky130_fd_sc_hd__xnor2_1
XFILLER_118_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07137_ _07137_/A _07327_/A _07137_/C vssd1 vssd1 vccd1 vccd1 _07139_/B sky130_fd_sc_hd__and3_1
XFILLER_134_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06243__A1 input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07068_ _10983_/Q _07197_/B vssd1 vssd1 vccd1 vccd1 _07312_/A sky130_fd_sc_hd__nand2_1
XFILLER_160_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06019_ _06019_/A _08212_/A vssd1 vssd1 vccd1 vccd1 _08258_/A sky130_fd_sc_hd__and2_1
XFILLER_102_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ _09710_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10981_ _10981_/CLK _10981_/D vssd1 vssd1 vccd1 vccd1 _10981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08054__A _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10415_ _10415_/A vssd1 vssd1 vccd1 vccd1 _10415_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10346_ _10355_/A vssd1 vssd1 vccd1 vccd1 _10346_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07982__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10277_ _10265_/A _10287_/B _10265_/B vssd1 vssd1 vccd1 vccd1 _10277_/X sky130_fd_sc_hd__o21ba_1
XFILLER_155_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06370_ _06409_/B vssd1 vssd1 vccd1 vccd1 _06408_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__06972__A _07715_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05321_ _10676_/Q vssd1 vssd1 vccd1 vccd1 _05830_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10254__C1 _08563_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08040_ _06115_/A _06115_/B _10580_/Q vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__o21a_1
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09991_ _10068_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08942_ _08965_/A _08965_/B vssd1 vssd1 vccd1 vccd1 _10518_/B sky130_fd_sc_hd__or2_2
XFILLER_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08873_ _08873_/A _08873_/B vssd1 vssd1 vccd1 vccd1 _08873_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06212__A _10517_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07725__A1 _07726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07824_ _10870_/Q _07824_/B vssd1 vssd1 vccd1 vccd1 _07824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07755_ _07755_/A _07755_/B vssd1 vssd1 vccd1 vccd1 _07756_/B sky130_fd_sc_hd__xnor2_1
XFILLER_72_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06706_ _06719_/A _06627_/B _06719_/C _06841_/A vssd1 vssd1 vccd1 vccd1 _06706_/X
+ sky130_fd_sc_hd__a22o_1
X_07686_ _09409_/A _09409_/B _07666_/A vssd1 vssd1 vccd1 vccd1 _07689_/A sky130_fd_sc_hd__o21a_1
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09425_ _09424_/A _09418_/A _09677_/B vssd1 vssd1 vccd1 vccd1 _09452_/B sky130_fd_sc_hd__a21o_1
X_06637_ _06638_/A _06638_/B vssd1 vssd1 vccd1 vccd1 _06715_/A sky130_fd_sc_hd__or2_1
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09356_ _09356_/A _10888_/Q vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__xnor2_4
X_06568_ _06568_/A _06568_/B _06581_/A vssd1 vssd1 vccd1 vccd1 _06570_/B sky130_fd_sc_hd__and3_1
XFILLER_166_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05519_ _07911_/A _05471_/X _05474_/Y _05442_/Y vssd1 vssd1 vccd1 vccd1 _10567_/D
+ sky130_fd_sc_hd__a22o_1
X_08307_ _05844_/A _08058_/X _08306_/Y _06011_/X vssd1 vssd1 vccd1 vccd1 _08307_/X
+ sky130_fd_sc_hd__o211a_1
X_09287_ _08342_/A _09286_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06499_ _06561_/B vssd1 vssd1 vccd1 vccd1 _06517_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08238_ _08114_/X _08251_/C _08233_/Y _08237_/X _06020_/X vssd1 vssd1 vccd1 vccd1
+ _08238_/X sky130_fd_sc_hd__o311a_1
XFILLER_166_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08169_ _08169_/A _08169_/B _08169_/C vssd1 vssd1 vccd1 vccd1 _08180_/B sky130_fd_sc_hd__and3_1
XFILLER_134_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10200_ _10197_/Y _10198_/Y _10199_/Y vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__o21a_1
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10131_ _10131_/A _10131_/B _10131_/C vssd1 vssd1 vccd1 vccd1 _10131_/X sky130_fd_sc_hd__and3_1
XANTENNA__08321__B _08355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _10062_/A _09338_/X vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__or2b_1
XFILLER_88_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07716__A1 _07442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10964_ _10985_/CLK _10964_/D vssd1 vssd1 vccd1 vccd1 _10964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08049__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08141__A1 _08058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10895_ _10909_/CLK _10895_/D vssd1 vssd1 vccd1 vccd1 _10895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07888__A _07906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_125_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _10334_/B _10327_/A _10329_/S vssd1 vssd1 vccd1 vccd1 _10330_/B sky130_fd_sc_hd__mux2_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09327__B _10283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06032__A _07910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05870_ _05358_/A _05823_/A _05869_/Y vssd1 vssd1 vccd1 vccd1 _05870_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07540_ _07540_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07540_/X sky130_fd_sc_hd__or2b_1
XFILLER_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07471_ _07471_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09210_ _09274_/A vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06422_ _06506_/B vssd1 vssd1 vccd1 vccd1 _06540_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09141_ _09153_/A _09141_/B vssd1 vssd1 vccd1 vccd1 _10843_/D sky130_fd_sc_hd__nor2_4
X_06353_ _06550_/B vssd1 vssd1 vccd1 vccd1 _06554_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_05304_ _10666_/Q _05358_/A vssd1 vssd1 vccd1 vccd1 _05353_/A sky130_fd_sc_hd__or2_1
X_09072_ _10936_/Q _10394_/C _10430_/B _10952_/Q vssd1 vssd1 vccd1 vccd1 _09072_/X
+ sky130_fd_sc_hd__a22o_1
X_06284_ _10918_/Q _07113_/A vssd1 vssd1 vccd1 vccd1 _06284_/X sky130_fd_sc_hd__and2_1
XANTENNA__06207__A _06238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08023_ _08023_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09974_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09975_/B sky130_fd_sc_hd__and2_1
XFILLER_131_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08925_ _08658_/X _08923_/Y _08924_/X vssd1 vssd1 vccd1 vccd1 _08926_/B sky130_fd_sc_hd__a21oi_1
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08856_ hold4/A _08856_/B vssd1 vssd1 vccd1 vccd1 _08857_/B sky130_fd_sc_hd__or2_1
XFILLER_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07807_ _07850_/A vssd1 vssd1 vccd1 vccd1 _07807_/X sky130_fd_sc_hd__buf_4
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05999_ input41/X vssd1 vssd1 vccd1 vccd1 _10528_/A sky130_fd_sc_hd__buf_6
XFILLER_84_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08787_ _06195_/X _08785_/X _08786_/X _10812_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08787_/X sky130_fd_sc_hd__o221a_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07738_ _07738_/A _07738_/B vssd1 vssd1 vccd1 vccd1 _07739_/B sky130_fd_sc_hd__xnor2_1
XFILLER_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07669_ _07669_/A vssd1 vssd1 vccd1 vccd1 _07673_/A sky130_fd_sc_hd__inv_2
XFILLER_164_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09408_ _10115_/A vssd1 vssd1 vccd1 vccd1 _09408_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_13_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10680_ _10684_/CLK _10680_/D vssd1 vssd1 vccd1 vccd1 _10680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09339_ _10911_/Q _10895_/Q vssd1 vssd1 vccd1 vccd1 _10065_/C sky130_fd_sc_hd__or2b_1
XFILLER_166_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05956__A _05956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08332__A _08332_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07937__A1 _05475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10114_ _10112_/Y _10113_/X _10880_/Q _09406_/X vssd1 vssd1 vccd1 vccd1 _10880_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_103_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10045_ _10045_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10110_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__06787__A _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08362__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08362__B2 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09311__B1 _10192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10947_ _10971_/CLK _10947_/D vssd1 vssd1 vccd1 vccd1 _10947_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10878_ _10970_/CLK _10878_/D vssd1 vssd1 vccd1 vccd1 _10878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06027__A _08201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09338__A _10912_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08242__A _08242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07928__B2 _07874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08050__B1 _10583_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _07655_/A vssd1 vssd1 vccd1 vccd1 _07715_/D sky130_fd_sc_hd__buf_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08710_ _08725_/B _08710_/B vssd1 vssd1 vccd1 vccd1 _08710_/Y sky130_fd_sc_hd__xnor2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05922_ _08130_/A _05900_/X _05897_/X _05896_/A _05921_/X vssd1 vssd1 vccd1 vccd1
+ _05922_/X sky130_fd_sc_hd__o221a_1
X_09690_ _09690_/A _09690_/B vssd1 vssd1 vccd1 vccd1 _09754_/A sky130_fd_sc_hd__xnor2_4
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05853_ _05340_/A _05854_/B _05852_/Y vssd1 vssd1 vccd1 vccd1 _05853_/X sky130_fd_sc_hd__o21a_1
X_08641_ _08641_/A vssd1 vssd1 vccd1 vccd1 _10795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05784_ _05803_/A _05769_/Y _05780_/Y _08304_/A _05783_/X vssd1 vssd1 vccd1 vccd1
+ _05785_/C sky130_fd_sc_hd__o221a_1
X_08572_ _10777_/Q _08572_/B _10775_/Q vssd1 vssd1 vccd1 vccd1 _08578_/D sky130_fd_sc_hd__and3_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07523_ _07525_/B _07523_/B vssd1 vssd1 vccd1 vccd1 _07649_/A sky130_fd_sc_hd__nand2_1
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07454_ _07454_/A _07454_/B _07454_/C vssd1 vssd1 vccd1 vccd1 _07455_/B sky130_fd_sc_hd__or3_1
XFILLER_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06405_ _06513_/D vssd1 vssd1 vccd1 vccd1 _06428_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_07385_ _07378_/Y _07458_/B _09304_/A _07384_/X vssd1 vssd1 vccd1 vccd1 _07386_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06336_ _06522_/B vssd1 vssd1 vccd1 vccd1 _06409_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_09124_ _09124_/A _09124_/B _09124_/C vssd1 vssd1 vccd1 vccd1 _09136_/A sky130_fd_sc_hd__nor3_4
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _05912_/B _08972_/X _08974_/A _09054_/X vssd1 vssd1 vccd1 vccd1 _09055_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_136_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06267_ _10916_/Q _10899_/Q vssd1 vssd1 vccd1 vccd1 _06267_/Y sky130_fd_sc_hd__nand2_1
XFILLER_136_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08006_ _08563_/A vssd1 vssd1 vccd1 vccd1 _08006_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06198_ _09403_/A vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__buf_2
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07395__A2 _07394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _09887_/A _09887_/B _09956_/X vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__a21o_1
XFILLER_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08908_ input36/X _08830_/X _08831_/X hold1/A vssd1 vssd1 vccd1 vccd1 _08908_/X sky130_fd_sc_hd__a22o_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _09626_/A _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09889_/B sky130_fd_sc_hd__a21boi_1
XFILLER_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08835_/Y _08836_/X _08838_/X vssd1 vssd1 vccd1 vccd1 _10818_/D sky130_fd_sc_hd__o21a_1
XFILLER_73_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ _10807_/CLK _10801_/D vssd1 vssd1 vccd1 vccd1 _10801_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10732_ _10807_/CLK _10732_/D vssd1 vssd1 vccd1 vccd1 _10732_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10663_ _10665_/CLK _10663_/D vssd1 vssd1 vccd1 vccd1 _10663_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10594_ _10653_/CLK _10594_/D vssd1 vssd1 vccd1 vccd1 _10594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08062__A _08062_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput61 _10848_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[14] sky130_fd_sc_hd__buf_2
Xoutput72 _10858_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[24] sky130_fd_sc_hd__buf_2
XFILLER_123_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput83 _10839_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[5] sky130_fd_sc_hd__buf_2
XFILLER_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_150_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10028_ _10100_/B _10028_/B vssd1 vssd1 vccd1 vccd1 _10029_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09195__A1_N _10946_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07170_ _07222_/A _07164_/B _07169_/B _07248_/A vssd1 vssd1 vccd1 vccd1 _07170_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_157_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06121_ _08483_/A _06121_/B vssd1 vssd1 vccd1 vccd1 _06122_/A sky130_fd_sc_hd__and2_1
XANTENNA__08271__B1 _08052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09068__A _10968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06052_ _06052_/A vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__buf_2
XFILLER_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09811_ _10493_/A _09811_/B _09811_/C vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__and3_1
XFILLER_98_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09133__A1_N _10940_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07019__C _07416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09742_ _09870_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09743_/B sky130_fd_sc_hd__or2_1
X_06954_ _07675_/B _07676_/B vssd1 vssd1 vccd1 vccd1 _07670_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05905_ _05905_/A _05905_/B vssd1 vssd1 vccd1 vccd1 _05906_/B sky130_fd_sc_hd__nand2_1
X_09673_ _09674_/A _09674_/B vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__or2_1
XFILLER_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06885_ _06885_/A _06885_/B vssd1 vssd1 vccd1 vccd1 _06886_/B sky130_fd_sc_hd__xnor2_4
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08624_ _10791_/Q _08624_/B _08628_/C vssd1 vssd1 vccd1 vccd1 _08631_/C sky130_fd_sc_hd__and3_1
X_05836_ _05836_/A _05836_/B vssd1 vssd1 vccd1 vccd1 _05836_/X sky130_fd_sc_hd__and2_1
XFILLER_82_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05767_ _10707_/Q vssd1 vssd1 vccd1 vccd1 _05767_/Y sky130_fd_sc_hd__clkinv_2
X_08555_ _08531_/X _08559_/B _10772_/Q _08531_/A vssd1 vssd1 vccd1 vccd1 _08557_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07506_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07507_/B sky130_fd_sc_hd__and2_1
XFILLER_23_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08486_ _10782_/Q hold8/A _08486_/S vssd1 vssd1 vccd1 vccd1 _08487_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08147__A _08150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05698_ _08181_/A _10553_/Q _10552_/Q _08173_/A vssd1 vssd1 vccd1 vccd1 _05717_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_168_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07437_ _06993_/A _07570_/C _07678_/A vssd1 vssd1 vccd1 vccd1 _07438_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09039__C1 _09263_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_53_clock _10682_/CLK vssd1 vssd1 vccd1 vccd1 _10851_/CLK sky130_fd_sc_hd__clkbuf_16
X_07368_ _07369_/B _07462_/A _07369_/A vssd1 vssd1 vccd1 vccd1 _07412_/C sky130_fd_sc_hd__o21a_1
XFILLER_109_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09107_ _09107_/A _09107_/B vssd1 vssd1 vccd1 vccd1 _09107_/Y sky130_fd_sc_hd__nand2_1
X_06319_ _10924_/Q _10907_/Q vssd1 vssd1 vccd1 vccd1 _06321_/A sky130_fd_sc_hd__nor2_1
XFILLER_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07299_ _07298_/A _07298_/B _07298_/C vssd1 vssd1 vccd1 vccd1 _07300_/B sky130_fd_sc_hd__a21oi_1
X_09038_ _10715_/Q _08999_/X _09037_/Y _10802_/Q vssd1 vssd1 vccd1 vccd1 _09038_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_68_clock _10840_/CLK vssd1 vssd1 vccd1 vccd1 _10651_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10372__A1 _06124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06040__A2 _08289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06067__A2_N _08235_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08057__A _08352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _10804_/CLK _10715_/D vssd1 vssd1 vccd1 vccd1 _10715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10646_ _10865_/CLK _10646_/D vssd1 vssd1 vccd1 vccd1 _10646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_5_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10577_ _10914_/CLK _10577_/D vssd1 vssd1 vccd1 vccd1 _10577_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_155_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output70_A _10856_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__A1 _08491_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06670_ _06670_/A _06670_/B vssd1 vssd1 vccd1 vccd1 _06671_/B sky130_fd_sc_hd__and2_1
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05621_ _10690_/Q vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_52_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05542__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10497__A _10497_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08340_ _05574_/X _08339_/C _05570_/X vssd1 vssd1 vccd1 vccd1 _08340_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07819__B1 _06257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05552_ _10551_/Q _05626_/A vssd1 vssd1 vccd1 vccd1 _05623_/A sky130_fd_sc_hd__or2_1
XFILLER_149_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08271_ input29/X _08212_/X _08052_/A _08267_/A _08201_/X vssd1 vssd1 vccd1 vccd1
+ _08272_/B sky130_fd_sc_hd__o221a_1
XFILLER_20_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05483_ _05483_/A _05489_/A vssd1 vssd1 vccd1 vccd1 _05483_/Y sky130_fd_sc_hd__nor2_1
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07222_ _07222_/A _07222_/B _07250_/A vssd1 vssd1 vccd1 vccd1 _07233_/B sky130_fd_sc_hd__and3_1
XFILLER_165_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07153_ _07295_/B _07317_/A _07295_/A vssd1 vssd1 vccd1 vccd1 _07153_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06104_ _10699_/Q _08243_/B vssd1 vssd1 vccd1 vccd1 _06105_/B sky130_fd_sc_hd__or2_1
XFILLER_106_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07084_ _07169_/B vssd1 vssd1 vccd1 vccd1 _07178_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06035_ _06035_/A _07974_/A vssd1 vssd1 vccd1 vccd1 _06035_/X sky130_fd_sc_hd__xor2_1
XFILLER_160_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07986_ _06191_/X _07965_/X _07985_/Y _07977_/X vssd1 vssd1 vccd1 vccd1 _10660_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09725_ _09779_/A _09779_/B _09661_/X vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__a21oi_1
XFILLER_41_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06937_ _06937_/A _06937_/B vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__xnor2_4
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09656_ _09656_/A _09656_/B vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__xor2_1
X_06868_ _06868_/A _06868_/B vssd1 vssd1 vccd1 vccd1 _06869_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09261__A _10441_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08607_ _08498_/X _08550_/X _08597_/B _10786_/Q vssd1 vssd1 vccd1 vccd1 _08608_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_82_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05819_ _05907_/A _05909_/A _05908_/B vssd1 vssd1 vccd1 vccd1 _05905_/B sky130_fd_sc_hd__a21o_1
X_09587_ _09587_/A _09587_/B vssd1 vssd1 vccd1 vccd1 _09591_/B sky130_fd_sc_hd__nand2_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ _10508_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07774_/A sky130_fd_sc_hd__nand2_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08567_/D vssd1 vssd1 vccd1 vccd1 _08580_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08469_ _08469_/A vssd1 vssd1 vccd1 vccd1 _10739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ _10517_/A _10500_/B vssd1 vssd1 vccd1 vccd1 _10515_/B sky130_fd_sc_hd__nor2_1
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10431_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10431_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _08491_/X _06855_/A _09408_/X _10929_/Q vssd1 vssd1 vccd1 vccd1 _10929_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06125__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10293_ _10351_/A vssd1 vssd1 vccd1 vccd1 _10293_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09436__A _09436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05964__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10345__A1 _09312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_clock_A clkbuf_3_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10629_ _10657_/CLK _10629_/D vssd1 vssd1 vccd1 vccd1 _10629_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__08226__B1 _06061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06035__A _06035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06252__A2 _06145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08529__A1 _06008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07840_ _07827_/X _05462_/A _07823_/X _07839_/Y vssd1 vssd1 vccd1 vccd1 _10623_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_96_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07771_ _07771_/A _07771_/B vssd1 vssd1 vccd1 vccd1 _07792_/A sky130_fd_sc_hd__xnor2_1
X_09510_ _09555_/B vssd1 vssd1 vccd1 vccd1 _09692_/A sky130_fd_sc_hd__buf_2
XFILLER_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06722_ _06722_/A vssd1 vssd1 vccd1 vccd1 _06722_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09441_ _09441_/A _07689_/A vssd1 vssd1 vccd1 vccd1 _09442_/B sky130_fd_sc_hd__or2b_1
X_06653_ _06650_/A _06650_/C _06650_/B vssd1 vssd1 vccd1 vccd1 _06654_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05604_ _05604_/A _05604_/B vssd1 vssd1 vccd1 vccd1 _05605_/B sky130_fd_sc_hd__and2_1
X_09372_ _09372_/A _09372_/B _09372_/C vssd1 vssd1 vccd1 vccd1 _09372_/X sky130_fd_sc_hd__or3_1
X_06584_ _06584_/A _06584_/B vssd1 vssd1 vccd1 vccd1 _06591_/A sky130_fd_sc_hd__or2_1
XFILLER_80_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08323_ _08881_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _10706_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05535_ _10544_/Q vssd1 vssd1 vccd1 vccd1 _05536_/B sky130_fd_sc_hd__inv_2
XFILLER_21_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10272__B1 _09480_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05466_ _07900_/A _07896_/A _07893_/A _07889_/A vssd1 vssd1 vccd1 vccd1 _05467_/D
+ sky130_fd_sc_hd__or4_1
X_08254_ _08242_/A _08243_/B _05598_/X vssd1 vssd1 vccd1 vccd1 _08254_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_166_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08425__A _08624_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07205_ _07205_/A _07205_/B vssd1 vssd1 vccd1 vccd1 _07302_/A sky130_fd_sc_hd__nand2_2
XANTENNA__06084__A1_N _05291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05397_ _05397_/A _05397_/B vssd1 vssd1 vccd1 vccd1 _05398_/B sky130_fd_sc_hd__nor2_1
X_08185_ _08185_/A _08185_/B vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__and2_1
XANTENNA__08768__A1 _06187_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07136_ _07136_/A _07136_/B vssd1 vssd1 vccd1 vccd1 _07138_/A sky130_fd_sc_hd__xnor2_1
XFILLER_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07067_ _07167_/B vssd1 vssd1 vccd1 vccd1 _07186_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06018_ _06023_/B vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08160__A _08160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10709__CLK _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10840__D _10840_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07969_ _07969_/A vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__05754__B2 _08242_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09708_ _09708_/A _09708_/B vssd1 vssd1 vccd1 vccd1 _09710_/B sky130_fd_sc_hd__nand2_1
X_10980_ _10980_/CLK _10980_/D vssd1 vssd1 vccd1 vccd1 _10980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _09588_/A _09639_/B _09696_/A vssd1 vssd1 vccd1 vccd1 _09640_/B sky130_fd_sc_hd__and3b_1
XFILLER_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07259__A1 _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05959__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06219__C1 _06200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _10942_/Q _10424_/B vssd1 vssd1 vccd1 vccd1 _10414_/X sky130_fd_sc_hd__and2_1
Xclkbuf_opt_4_0_clock clkbuf_3_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _10853_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10345_ _09312_/X _07682_/B _10184_/X _10915_/Q vssd1 vssd1 vccd1 vccd1 _10915_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10276_ _10287_/C _10287_/D vssd1 vssd1 vccd1 vccd1 _10276_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05993__A1 _09107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08931__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05320_ _10645_/Q vssd1 vssd1 vccd1 vccd1 _07922_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08998__A1 _08062_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05869__A _08000_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09990_ _09990_/A _09990_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__xnor2_2
XFILLER_89_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08941_ _09098_/B vssd1 vssd1 vccd1 vccd1 _08965_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_115_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05984__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08872_ _10822_/Q hold4/A _10820_/Q _08847_/X _08840_/B vssd1 vssd1 vccd1 vccd1 _08873_/B
+ sky130_fd_sc_hd__o41a_1
XFILLER_96_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06212__B _06212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07823_ _08557_/A vssd1 vssd1 vccd1 vccd1 _07823_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07754_ _07754_/A _07754_/B vssd1 vssd1 vccd1 vccd1 _07755_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06705_ _06719_/A _06719_/C vssd1 vssd1 vccd1 vccd1 _07791_/A sky130_fd_sc_hd__nand2_1
XFILLER_25_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ _09329_/A _09329_/B _07674_/A vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__o21a_2
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09424_ _09424_/A _09811_/B _09677_/B vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__nand3_1
XFILLER_25_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06636_ _06431_/A _06431_/B _06434_/A vssd1 vssd1 vccd1 vccd1 _06638_/B sky130_fd_sc_hd__o21a_1
XANTENNA__06161__A1 _05982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _10905_/Q _10889_/Q vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__or2b_1
X_06567_ _06567_/A _06567_/B vssd1 vssd1 vccd1 vccd1 _06581_/A sky130_fd_sc_hd__nand2_1
X_08306_ _08317_/B _08306_/B _08306_/C vssd1 vssd1 vccd1 vccd1 _08306_/Y sky130_fd_sc_hd__nand3_1
X_05518_ _05332_/Y _05517_/X _05513_/X _07907_/A vssd1 vssd1 vccd1 vccd1 _10566_/D
+ sky130_fd_sc_hd__a2bb2o_1
X_09286_ _08339_/A _07922_/A _09296_/S vssd1 vssd1 vccd1 vccd1 _09286_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06498_ _10972_/Q vssd1 vssd1 vccd1 vccd1 _06561_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_165_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08237_ _08243_/B _08061_/A _08234_/X _08235_/Y _08236_/X vssd1 vssd1 vccd1 vccd1
+ _08237_/X sky130_fd_sc_hd__a311o_1
XANTENNA__10835__D _10835_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05449_ _10647_/Q _05525_/B _05448_/X vssd1 vssd1 vccd1 vccd1 _05490_/A sky130_fd_sc_hd__o21ai_4
XFILLER_154_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_clock_A _10709_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08168_ _08157_/X _08161_/X _08163_/Y _08167_/X vssd1 vssd1 vccd1 vccd1 _10690_/D
+ sky130_fd_sc_hd__o31a_1
X_07119_ _10983_/Q _07142_/B vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__and2_1
XFILLER_134_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08099_ _08038_/X _08074_/X _08098_/Y _08044_/X _05905_/A vssd1 vssd1 vccd1 vccd1
+ _08099_/X sky130_fd_sc_hd__a32o_1
XANTENNA__08602__B _08649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10130_ _10130_/A _10130_/B vssd1 vssd1 vccd1 vccd1 _10133_/A sky130_fd_sc_hd__nor2_1
XFILLER_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__xor2_1
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_102_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05727__B2 _08117_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05961__B input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10963_ _10967_/CLK _10963_/D vssd1 vssd1 vccd1 vccd1 _10963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ _10909_/CLK _10894_/D vssd1 vssd1 vccd1 vccd1 _10894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ _10312_/A _10310_/X _10320_/A _10327_/Y vssd1 vssd1 vccd1 vccd1 _10334_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_125_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10243_/A _10250_/X _10245_/B vssd1 vssd1 vccd1 vccd1 _10259_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08668__B1 _10799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07470_ _07470_/A _07470_/B _07482_/A vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__nor3_1
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06421_ _06421_/A _06732_/B vssd1 vssd1 vccd1 vccd1 _06506_/B sky130_fd_sc_hd__xnor2_2
XFILLER_50_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09140_ _09112_/X _09135_/Y _09139_/X vssd1 vssd1 vccd1 vccd1 _09141_/B sky130_fd_sc_hd__a21oi_1
X_06352_ _06352_/A _06352_/B _06352_/C vssd1 vssd1 vccd1 vccd1 _06550_/B sky130_fd_sc_hd__or3_1
XFILLER_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05303_ _10665_/Q _10664_/Q _05363_/A vssd1 vssd1 vccd1 vccd1 _05358_/A sky130_fd_sc_hd__or3_2
X_09071_ _09904_/A vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__buf_4
X_06283_ _10901_/Q vssd1 vssd1 vccd1 vccd1 _07113_/A sky130_fd_sc_hd__buf_2
X_08022_ input33/X _08015_/X _08021_/Y _08019_/X vssd1 vssd1 vccd1 vccd1 _10673_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_144_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09973_ _09974_/A _09974_/B vssd1 vssd1 vccd1 vccd1 _09975_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08924_ input39/X _08830_/X _08831_/X hold9/A vssd1 vssd1 vccd1 vccd1 _08924_/X sky130_fd_sc_hd__a22o_1
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09534__A _10968_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08855_ hold4/X _08865_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__nand2_1
XFILLER_130_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07806_ _10160_/A _07804_/Y _07805_/X _10881_/Q vssd1 vssd1 vccd1 vccd1 _07850_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08786_ _08820_/A vssd1 vssd1 vccd1 vccd1 _08786_/X sky130_fd_sc_hd__clkbuf_2
X_05998_ _09090_/A vssd1 vssd1 vccd1 vccd1 _08483_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07737_ _07581_/A _07581_/B _07580_/A vssd1 vssd1 vccd1 vccd1 _07738_/B sky130_fd_sc_hd__o21a_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07668_ _07668_/A _07668_/B vssd1 vssd1 vccd1 vccd1 _07669_/A sky130_fd_sc_hd__xnor2_1
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09407_ _09402_/X _09405_/X _10868_/Q _09406_/X vssd1 vssd1 vccd1 vccd1 _10868_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06619_ _06668_/A _06668_/B _06618_/X vssd1 vssd1 vccd1 vccd1 _06692_/A sky130_fd_sc_hd__a21o_2
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07599_/X sky130_fd_sc_hd__or2_1
X_09338_ _10912_/Q _10896_/Q vssd1 vssd1 vccd1 vccd1 _09338_/X sky130_fd_sc_hd__or2b_1
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09269_ _08318_/A _09268_/X _09287_/S vssd1 vssd1 vccd1 vccd1 _09269_/X sky130_fd_sc_hd__mux2_1
XFILLER_138_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10113_ _10112_/A _10112_/B _09480_/X vssd1 vssd1 vccd1 vccd1 _10113_/X sky130_fd_sc_hd__a21o_1
XFILLER_122_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input32_A io_wbs_m2s_data[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10044_ _10879_/Q _09572_/X _10042_/Y _10043_/X vssd1 vssd1 vccd1 vccd1 _10879_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08898__B1 _08688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09311__A1 _10043_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__A _07899_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10946_ _10958_/CLK _10946_/D vssd1 vssd1 vccd1 vccd1 _10946_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09610__C _09610_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ _10970_/CLK _10877_/D vssd1 vssd1 vccd1 vccd1 _10877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06027__B _09403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_172_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08050__A1 _10369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06970_ _07678_/A vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05921_ _05726_/A _05902_/Y _05900_/X _10687_/Q _05920_/X vssd1 vssd1 vccd1 vccd1
+ _05921_/X sky130_fd_sc_hd__a221o_1
XFILLER_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08640_ _08638_/X _08640_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _08641_/A sky130_fd_sc_hd__and3b_1
X_05852_ _08289_/A _05852_/B vssd1 vssd1 vccd1 vccd1 _05852_/Y sky130_fd_sc_hd__nand2_1
XFILLER_81_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08571_ _08572_/B _08565_/X _10777_/Q vssd1 vssd1 vccd1 vccd1 _08574_/B sky130_fd_sc_hd__a21o_1
X_05783_ _05781_/Y _10566_/Q _10565_/Q _05782_/Y vssd1 vssd1 vccd1 vccd1 _05783_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_19_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07522_ _07522_/A _07522_/B vssd1 vssd1 vccd1 vccd1 _07523_/B sky130_fd_sc_hd__or2_1
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07453_ _07454_/B _07454_/C _07454_/A vssd1 vssd1 vccd1 vccd1 _07455_/A sky130_fd_sc_hd__o21ai_2
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06404_ _06461_/B vssd1 vssd1 vccd1 vccd1 _06426_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07384_ _07384_/A _07384_/B vssd1 vssd1 vccd1 vccd1 _07384_/X sky130_fd_sc_hd__xor2_1
X_09123_ _09263_/A vssd1 vssd1 vccd1 vccd1 _09123_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_06335_ _06515_/B vssd1 vssd1 vccd1 vccd1 _06522_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__08813__B1 _05983_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09054_ _05905_/A _08995_/X _09053_/X _08981_/A vssd1 vssd1 vccd1 vccd1 _09054_/X
+ sky130_fd_sc_hd__a211o_1
X_06266_ _10916_/Q _10899_/Q vssd1 vssd1 vccd1 vccd1 _06360_/A sky130_fd_sc_hd__xnor2_2
XFILLER_135_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08005_ _08244_/A _08005_/B vssd1 vssd1 vccd1 vccd1 _08005_/X sky130_fd_sc_hd__or2_1
X_06197_ _06197_/A _06204_/B vssd1 vssd1 vccd1 vccd1 _06197_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09956_ _09886_/B _09956_/B vssd1 vssd1 vccd1 vccd1 _09956_/X sky130_fd_sc_hd__and2b_1
XFILLER_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08907_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09887_/A _09887_/B vssd1 vssd1 vccd1 vccd1 _09890_/B sky130_fd_sc_hd__xor2_1
XFILLER_57_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ input26/X _08785_/X _08786_/X _10818_/Q _08837_/X vssd1 vssd1 vccd1 vccd1
+ _08838_/X sky130_fd_sc_hd__o221a_1
XFILLER_131_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08769_ _08766_/Y _08767_/X _08768_/X vssd1 vssd1 vccd1 vccd1 _10810_/D sky130_fd_sc_hd__o21a_1
XFILLER_61_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _10833_/CLK _10800_/D vssd1 vssd1 vccd1 vccd1 _10800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10731_ _10807_/CLK _10731_/D vssd1 vssd1 vccd1 vccd1 _10731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10662_ _10665_/CLK _10662_/D vssd1 vssd1 vccd1 vccd1 _10662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_139_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06128__A _09250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10593_ _10652_/CLK _10593_/D vssd1 vssd1 vccd1 vccd1 _10593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_154_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05967__A input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06026__A_N _10581_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput62 _10849_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[15] sky130_fd_sc_hd__buf_2
Xoutput73 _10859_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[25] sky130_fd_sc_hd__buf_2
XFILLER_68_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput84 _10840_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[6] sky130_fd_sc_hd__buf_2
XFILLER_110_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10027_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__or2_1
XFILLER_76_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09296__A0 _06115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08099__B2 _05905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10929_ _10929_/CLK _10929_/D vssd1 vssd1 vccd1 vccd1 _10929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06120_ input16/X _06019_/A _06120_/S vssd1 vssd1 vccd1 vccd1 _06121_/B sky130_fd_sc_hd__mux2_1
XFILLER_173_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08271__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08271__B2 _08267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_79_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06051_ _08130_/A vssd1 vssd1 vccd1 vccd1 _09104_/A sky130_fd_sc_hd__inv_2
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09220__A0 _08233_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09810_ _09810_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09811_/C sky130_fd_sc_hd__nand2_1
XFILLER_99_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09741_ _10480_/A _10129_/B _10122_/B _10478_/A vssd1 vssd1 vccd1 vccd1 _09742_/B
+ sky130_fd_sc_hd__a22oi_1
X_06953_ _06769_/A _06460_/B _06558_/X vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08326__A2 _08058_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05904_ _05904_/A _05904_/B vssd1 vssd1 vccd1 vccd1 _05904_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09672_ _09670_/Y _09672_/B vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__and2b_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06884_ _06884_/A _06884_/B vssd1 vssd1 vccd1 vccd1 _06886_/A sky130_fd_sc_hd__or2_2
XFILLER_95_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08623_ _10790_/Q _10789_/Q _08623_/C _08623_/D vssd1 vssd1 vccd1 vccd1 _08628_/C
+ sky130_fd_sc_hd__and4_1
X_05835_ _08025_/A _05838_/B _08027_/A vssd1 vssd1 vccd1 vccd1 _05836_/B sky130_fd_sc_hd__o21ai_1
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09287__A0 _08342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08554_ _08583_/A _08554_/B vssd1 vssd1 vccd1 vccd1 _10771_/D sky130_fd_sc_hd__nor2_1
XFILLER_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05766_ _10708_/Q vssd1 vssd1 vccd1 vccd1 _05766_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07505_ _07505_/A _07505_/B vssd1 vssd1 vccd1 vccd1 _07505_/X sky130_fd_sc_hd__and2_1
XFILLER_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ _09090_/A vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05697_ _05885_/A vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__clkinv_2
XFILLER_50_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07436_ _07727_/A _07433_/A _07729_/B _07713_/A vssd1 vssd1 vccd1 vccd1 _07445_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07367_ _07412_/B _07367_/B vssd1 vssd1 vccd1 vccd1 _07369_/A sky130_fd_sc_hd__nor2_1
XFILLER_164_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09106_ _06050_/X _08995_/A _09105_/X _09107_/B vssd1 vssd1 vccd1 vccd1 _09106_/X
+ sky130_fd_sc_hd__a211o_1
X_06318_ _06755_/A _06729_/A vssd1 vssd1 vccd1 vccd1 _06318_/X sky130_fd_sc_hd__or2_1
X_07298_ _07298_/A _07298_/B _07298_/C vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__and3_1
XFILLER_164_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10843__D _10843_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09037_ _09037_/A _09079_/A vssd1 vssd1 vccd1 vccd1 _09037_/Y sky130_fd_sc_hd__nor2_1
X_06249_ _10613_/Q _06249_/B vssd1 vssd1 vccd1 vccd1 _06249_/X sky130_fd_sc_hd__or2_1
XFILLER_136_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08014__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09939_ _09940_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _10009_/B sky130_fd_sc_hd__or2_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07941__S _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10804_/CLK _10714_/D vssd1 vssd1 vccd1 vccd1 _10714_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10645_ _10865_/CLK _10645_/D vssd1 vssd1 vccd1 vccd1 _10645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09345__A_N _09344_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09169__A _09270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10576_ _10652_/CLK _10576_/D vssd1 vssd1 vccd1 vccd1 _10576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_155_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_80_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10363__A2 _07635_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09632__A _09757_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09269__A0 _08318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05620_ _10692_/Q vssd1 vssd1 vccd1 vccd1 _05885_/A sky130_fd_sc_hd__buf_2
XANTENNA__08248__A _08248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05551_ _10550_/Q _10549_/Q _05630_/A vssd1 vssd1 vccd1 vccd1 _05626_/A sky130_fd_sc_hd__or3_1
XFILLER_33_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08270_ _08263_/X _08276_/B _08266_/Y _08269_/X _08258_/X vssd1 vssd1 vccd1 vccd1
+ _08270_/X sky130_fd_sc_hd__o311a_1
XANTENNA__06991__A _07166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05482_ _10574_/Q vssd1 vssd1 vccd1 vccd1 _05482_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_149_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07221_ _07250_/A _07217_/B _07218_/X _07242_/B vssd1 vssd1 vccd1 vccd1 _07233_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_146_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07152_ _07309_/A _07152_/B _07322_/A vssd1 vssd1 vccd1 vccd1 _07317_/A sky130_fd_sc_hd__and3_1
XFILLER_121_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06103_ _10698_/Q _10697_/Q _10696_/Q _08218_/B vssd1 vssd1 vccd1 vccd1 _08243_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_161_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07083_ _07083_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07169_/B sky130_fd_sc_hd__xnor2_4
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06034_ _10686_/Q vssd1 vssd1 vccd1 vccd1 _08115_/A sky130_fd_sc_hd__inv_2
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07985_ _07985_/A _07985_/B vssd1 vssd1 vccd1 vccd1 _07985_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09724_ _09724_/A _09723_/Y vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__or2b_1
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06936_ _06936_/A _06936_/B vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__xnor2_4
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09655_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09656_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06867_ _06866_/B _06867_/B vssd1 vssd1 vccd1 vccd1 _06868_/B sky130_fd_sc_hd__and2b_1
XFILLER_28_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08606_ _10786_/Q _10785_/Q _08617_/B vssd1 vssd1 vccd1 vccd1 _08611_/B sky130_fd_sc_hd__and3_1
X_05818_ _05818_/A _05818_/B vssd1 vssd1 vccd1 vccd1 _05908_/B sky130_fd_sc_hd__nor2_1
X_09586_ _09639_/B _09834_/B _09642_/A _09696_/A vssd1 vssd1 vccd1 vccd1 _09587_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ _06845_/A vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__buf_2
XANTENNA__08158__A _08160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07062__A _07164_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10838__D _10838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _10291_/S _08686_/A _08462_/A vssd1 vssd1 vccd1 vccd1 _08567_/D sky130_fd_sc_hd__a21oi_2
X_05749_ _05749_/A _10564_/Q vssd1 vssd1 vccd1 vccd1 _05749_/X sky130_fd_sc_hd__and2_1
XFILLER_168_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08468_ _08477_/A _08468_/B vssd1 vssd1 vccd1 vccd1 _08469_/A sky130_fd_sc_hd__or2_1
XFILLER_168_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07419_ _07416_/A _07727_/B _07713_/B _07567_/A vssd1 vssd1 vccd1 vccd1 _07419_/X
+ sky130_fd_sc_hd__a22o_1
X_08399_ _08408_/A _10756_/Q vssd1 vssd1 vccd1 vccd1 _08399_/X sky130_fd_sc_hd__or2_1
XFILLER_7_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10430_ _10495_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__nand2_1
XFILLER_109_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ _08491_/X _06853_/B _10355_/X _10928_/Q vssd1 vssd1 vccd1 vccd1 _10928_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09717__A _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10292_/X sky130_fd_sc_hd__xor2_2
XFILLER_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__05964__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10345__A2 _07682_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_1_1_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05980__A input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_clock_A _10977_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08171__B1 _05692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10628_ _10657_/CLK _10628_/D vssd1 vssd1 vccd1 vccd1 _10628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_128_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10559_ _10562_/CLK _10559_/D vssd1 vssd1 vccd1 vccd1 _10559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__06788__A1 _10506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06035__B _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05874__B _05883_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07770_ _06864_/A _06864_/B _06863_/A vssd1 vssd1 vccd1 vccd1 _07771_/B sky130_fd_sc_hd__a21oi_1
XFILLER_110_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_clock _10709_/CLK vssd1 vssd1 vccd1 vccd1 _10562_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06721_ _06721_/A vssd1 vssd1 vccd1 vccd1 _06721_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08162__B1 _08067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _10869_/Q _09408_/X _09438_/Y _09439_/X vssd1 vssd1 vccd1 vccd1 _10869_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06652_ _06702_/B _06652_/B vssd1 vssd1 vccd1 vccd1 _06893_/A sky130_fd_sc_hd__xnor2_4
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05603_ _10558_/Q _05610_/A _10559_/Q vssd1 vssd1 vccd1 vccd1 _05604_/B sky130_fd_sc_hd__o21ai_1
X_09371_ _09371_/A _09371_/B vssd1 vssd1 vccd1 vccd1 _09372_/C sky130_fd_sc_hd__nor2_1
X_06583_ _06568_/A _06459_/B _06576_/B _10973_/Q vssd1 vssd1 vccd1 vccd1 _06584_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_67_clock clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _10970_/CLK sky130_fd_sc_hd__clkbuf_16
X_08322_ _08314_/Y _08086_/X _08157_/A _08320_/X _08321_/X vssd1 vssd1 vccd1 vccd1
+ _08323_/B sky130_fd_sc_hd__o221a_1
X_05534_ _09107_/A _10544_/Q vssd1 vssd1 vccd1 vccd1 _05652_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10272__A1 _10287_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08253_ _08255_/A vssd1 vssd1 vccd1 vccd1 _08253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05465_ _07885_/A _07882_/A _07878_/A _07875_/A vssd1 vssd1 vccd1 vccd1 _05467_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_21_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07204_ _07204_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07205_/B sky130_fd_sc_hd__nand2_1
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08184_ input19/X _08123_/X _08109_/X _08180_/A _08125_/X vssd1 vssd1 vccd1 vccd1
+ _08185_/B sky130_fd_sc_hd__o221a_1
XANTENNA__06226__A _06253_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05396_ _10652_/Q _05452_/A vssd1 vssd1 vccd1 vccd1 _05397_/A sky130_fd_sc_hd__nor2_1
XFILLER_146_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07135_ _07135_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07136_/B sky130_fd_sc_hd__nor2_1
XFILLER_134_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07066_ _07066_/A _07066_/B vssd1 vssd1 vccd1 vccd1 _07167_/B sky130_fd_sc_hd__xnor2_4
XFILLER_160_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06017_ _10341_/A _09124_/B _09098_/A vssd1 vssd1 vccd1 vccd1 _06023_/B sky130_fd_sc_hd__or3_4
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07968_ _08971_/B _08989_/A vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__nand2_1
XFILLER_102_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09707_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__or2_1
X_06919_ _06748_/X _06940_/B _06918_/X vssd1 vssd1 vccd1 vccd1 _06939_/B sky130_fd_sc_hd__a21oi_4
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07899_ _07899_/A vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09638_ _09769_/A _09744_/B _09638_/C vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__and3_1
XFILLER_71_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09569_ _09527_/A _09527_/B _09568_/X vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__a21bo_1
XFILLER_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05959__B input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06136__A _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05690__A1 _05528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _10408_/X _10722_/Q _10410_/X _10411_/X _10412_/X vssd1 vssd1 vccd1 vccd1
+ _10941_/D sky130_fd_sc_hd__o221a_1
XFILLER_125_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10344_ _10344_/A vssd1 vssd1 vccd1 vccd1 _10914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08351__A _08351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10275_ _10940_/Q _10956_/Q vssd1 vssd1 vccd1 vccd1 _10287_/D sky130_fd_sc_hd__or2b_1
XFILLER_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10254__A1 _07061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07958__A0 _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08940_ _09142_/D vssd1 vssd1 vccd1 vccd1 _09098_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08871_ _08871_/A _08871_/B vssd1 vssd1 vccd1 vccd1 _08871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07822_ _06255_/X _05455_/X _06257_/X _07821_/Y vssd1 vssd1 vccd1 vccd1 _10619_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_29_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__07605__A _07708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _07753_/A _07753_/B vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__xor2_1
XFILLER_65_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ _06885_/A _06885_/B _06642_/A vssd1 vssd1 vccd1 vccd1 _06876_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__08280__A1_N _05851_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ _07681_/A _07681_/B _09314_/A vssd1 vssd1 vccd1 vccd1 _09329_/B sky130_fd_sc_hd__o21ba_2
XFILLER_80_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09423_ _09423_/A vssd1 vssd1 vccd1 vccd1 _09677_/B sky130_fd_sc_hd__inv_2
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06635_ _06719_/B _06635_/B vssd1 vssd1 vccd1 vccd1 _06638_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09354_ _09372_/A _09734_/A _09674_/A vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__or3_1
XFILLER_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06566_ _06571_/B _06571_/C _06571_/A vssd1 vssd1 vccd1 vccd1 _06570_/A sky130_fd_sc_hd__a21bo_1
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08436__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ _08305_/A _08305_/B vssd1 vssd1 vccd1 vccd1 _08306_/C sky130_fd_sc_hd__nand2_1
X_05517_ _05517_/A vssd1 vssd1 vccd1 vccd1 _05517_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_09285_ _09285_/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__clkbuf_1
XFILLER_138_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06497_ _06502_/B _06515_/B vssd1 vssd1 vccd1 vccd1 _06517_/C sky130_fd_sc_hd__and2_1
XFILLER_166_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08236_ _08236_/A vssd1 vssd1 vccd1 vccd1 _08236_/X sky130_fd_sc_hd__clkbuf_2
X_05448_ _10647_/Q _05525_/B _05318_/X _07925_/A _05447_/X vssd1 vssd1 vccd1 vccd1
+ _05448_/X sky130_fd_sc_hd__a221o_1
XFILLER_166_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ input17/X _08164_/X _08165_/X _08158_/X _08394_/A vssd1 vssd1 vccd1 vccd1
+ _08167_/X sky130_fd_sc_hd__o221a_1
X_05379_ _10657_/Q _05383_/A vssd1 vssd1 vccd1 vccd1 _05380_/B sky130_fd_sc_hd__and2_1
XFILLER_107_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09267__A _09267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ _07150_/A _07135_/B _07117_/X vssd1 vssd1 vccd1 vccd1 _07145_/A sky130_fd_sc_hd__o21ai_1
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08098_ _08098_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08098_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07049_ _07473_/A _07463_/B vssd1 vssd1 vccd1 vccd1 _07464_/A sky130_fd_sc_hd__nor2_1
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10060_ _10491_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__nand2_1
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08126__B1 _08124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10962_ _10962_/CLK _10962_/D vssd1 vssd1 vccd1 vccd1 _10962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10893_ _10909_/CLK _10893_/D vssd1 vssd1 vccd1 vccd1 _10893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10327_ _10327_/A vssd1 vssd1 vccd1 vccd1 _10327_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _10243_/A _10249_/A _10245_/B vssd1 vssd1 vccd1 vccd1 _10258_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_59_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10189_ _10931_/Q _10947_/Q vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__and2b_1
XFILLER_66_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__06083__A1_N _05766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06420_ _06420_/A _06420_/B vssd1 vssd1 vccd1 vccd1 _06732_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08256__A _08256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06351_ _06895_/A vssd1 vssd1 vccd1 vccd1 _06365_/B sky130_fd_sc_hd__clkinv_2
XFILLER_148_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05302_ _10663_/Q _05362_/B vssd1 vssd1 vccd1 vccd1 _05363_/A sky130_fd_sc_hd__or2_1
X_09070_ _09834_/A vssd1 vssd1 vccd1 vccd1 _09904_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06282_ _06352_/A _06352_/B vssd1 vssd1 vccd1 vccd1 _06371_/B sky130_fd_sc_hd__nand2_1
XFILLER_129_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08021_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09972_ _09971_/Y _09906_/A _09905_/B vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__a21o_1
XFILLER_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08923_ _08927_/C _08923_/B vssd1 vssd1 vccd1 vccd1 _08923_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_103_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08356__B1 _08157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08854_ _08814_/X _08852_/X _08853_/X vssd1 vssd1 vccd1 vccd1 _10820_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07805_ _10160_/A _10117_/A _10117_/B vssd1 vssd1 vccd1 vccd1 _07805_/X sky130_fd_sc_hd__and3b_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_08785_ _08819_/A vssd1 vssd1 vccd1 vccd1 _08785_/X sky130_fd_sc_hd__buf_2
XFILLER_38_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05997_ _09403_/A vssd1 vssd1 vccd1 vccd1 _09090_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07736_ _07729_/A _07728_/B _07565_/B _07563_/X vssd1 vssd1 vccd1 vccd1 _07738_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09550__A _09610_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10466__A1 _06191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _07678_/A _07667_/B vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09406_ _10192_/A vssd1 vssd1 vccd1 vccd1 _09406_/X sky130_fd_sc_hd__buf_2
X_06618_ _06618_/A _06618_/B vssd1 vssd1 vccd1 vccd1 _06618_/X sky130_fd_sc_hd__and2_1
XFILLER_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07598_ _07598_/A vssd1 vssd1 vccd1 vccd1 _07598_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08166__A _08166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10846__D _10846_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ _09387_/A _09337_/B vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__or2_2
X_06549_ _06549_/A _06549_/B vssd1 vssd1 vccd1 vccd1 _06571_/B sky130_fd_sc_hd__nor2_1
XFILLER_166_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09268_ _08317_/A _07911_/A _09276_/S vssd1 vssd1 vccd1 vccd1 _09268_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08292__C1 _08175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06117__C _06117_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ _07998_/A _08306_/B _08217_/X _08228_/B _06011_/X vssd1 vssd1 vccd1 vccd1
+ _08219_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ _08209_/A _09226_/S _09203_/A _09198_/X vssd1 vssd1 vccd1 vccd1 _09199_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10112_ _10112_/A _10112_/B vssd1 vssd1 vccd1 vccd1 _10112_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07944__S _07964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10043_ _10043_/A vssd1 vssd1 vccd1 vccd1 _10043_/X sky130_fd_sc_hd__buf_2
XFILLER_76_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input25_A io_wbs_m2s_data[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10945_ _10945_/CLK _10945_/D vssd1 vssd1 vccd1 vccd1 _10945_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__D _09717_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ _10970_/CLK _10876_/D vssd1 vssd1 vccd1 vccd1 _10876_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__05884__A1 _07988_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08035__C1 _08030_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ _06037_/A _05904_/Y _05902_/Y _10686_/Q _05919_/X vssd1 vssd1 vccd1 vccd1
+ _05920_/X sky130_fd_sc_hd__o221a_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_05851_ _05851_/A _10669_/Q _05857_/B vssd1 vssd1 vccd1 vccd1 _05852_/B sky130_fd_sc_hd__or3_1
XFILLER_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08570_ _08572_/B _08565_/X _08569_/Y vssd1 vssd1 vccd1 vccd1 _10776_/D sky130_fd_sc_hd__o21a_1
XFILLER_54_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05782_ _10704_/Q vssd1 vssd1 vccd1 vccd1 _05782_/Y sky130_fd_sc_hd__inv_2
XFILLER_148_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_75_clock_A clkbuf_3_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07521_ _07657_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07648_/B sky130_fd_sc_hd__or2_1
XFILLER_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07452_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07454_/A sky130_fd_sc_hd__xor2_1
XFILLER_35_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06403_ _10976_/Q vssd1 vssd1 vccd1 vccd1 _06461_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__05875__A1 _08198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07383_ _07459_/B _07748_/B _07381_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07384_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09066__A1 _05482_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09122_ _09113_/X _09120_/X _09121_/X vssd1 vssd1 vccd1 vccd1 _09122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06334_ _06371_/A _06334_/B vssd1 vssd1 vccd1 vccd1 _06515_/B sky130_fd_sc_hd__xor2_4
XFILLER_109_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _05453_/A _08978_/A _06129_/B _08098_/A _09179_/A vssd1 vssd1 vccd1 vccd1
+ _09053_/X sky130_fd_sc_hd__o221a_1
XFILLER_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06265_ _10915_/Q _10898_/Q vssd1 vssd1 vccd1 vccd1 _06558_/B sky130_fd_sc_hd__nand2_2
XFILLER_117_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08004_ input25/X _08002_/X _08003_/X _07993_/X vssd1 vssd1 vccd1 vccd1 _10666_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06196_ _10597_/Q vssd1 vssd1 vccd1 vccd1 _06197_/A sky130_fd_sc_hd__inv_2
XFILLER_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09955_ _09955_/A _09955_/B vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__xnor2_1
X_08906_ _08889_/X _08891_/X _08896_/X _08905_/X vssd1 vssd1 vccd1 vccd1 _08907_/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_98_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09956_/B _09886_/B vssd1 vssd1 vccd1 vccd1 _09887_/B sky130_fd_sc_hd__xnor2_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08837_/A vssd1 vssd1 vccd1 vccd1 _08837_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _06187_/X _08694_/X _08695_/X _10810_/Q _08737_/X vssd1 vssd1 vccd1 vccd1
+ _08768_/X sky130_fd_sc_hd__o221a_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09280__A _09280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_07719_ _07391_/A _07391_/B _07588_/B _07596_/A _07718_/Y vssd1 vssd1 vccd1 vccd1
+ _07720_/B sky130_fd_sc_hd__a32o_1
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _10803_/Q _08732_/B vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__and2_1
XFILLER_26_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__08608__B _08649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10730_ _10807_/CLK _10730_/D vssd1 vssd1 vccd1 vccd1 _10730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10661_ _10665_/CLK _10661_/D vssd1 vssd1 vccd1 vccd1 _10661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10592_ _10652_/CLK _10592_/D vssd1 vssd1 vccd1 vccd1 _10592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05967__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput52 _10581_/Q vssd1 vssd1 vccd1 vccd1 io_motor_irq sky130_fd_sc_hd__buf_2
XANTENNA__05983__A _08445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput63 _10850_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[16] sky130_fd_sc_hd__buf_2
Xoutput74 _10860_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[26] sky130_fd_sc_hd__buf_2
XFILLER_96_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput85 _10841_/Q vssd1 vssd1 vccd1 vccd1 io_wbs_data_o[7] sky130_fd_sc_hd__buf_2
XFILLER_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10026_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10928_ _10929_/CLK _10928_/D vssd1 vssd1 vccd1 vccd1 _10928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10859_ _10859_/CLK _10859_/D vssd1 vssd1 vccd1 vccd1 _10859_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08534__A _10251_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_06050_ _10655_/Q vssd1 vssd1 vccd1 vccd1 _06050_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06952_ _06952_/A _06952_/B vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__nor2_1
X_09740_ _09930_/C vssd1 vssd1 vccd1 vccd1 _10122_/B sky130_fd_sc_hd__dlymetal6s2s_1
.ends

