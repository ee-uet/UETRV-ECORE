magic
tech sky130A
magscale 1 2
timestamp 1649144880
<< obsli1 >>
rect 1104 2159 108836 107729
<< obsm1 >>
rect 1104 1980 108836 107760
<< metal2 >>
rect 6090 109200 6146 110000
rect 18234 109200 18290 110000
rect 30470 109200 30526 110000
rect 42706 109200 42762 110000
rect 54942 109200 54998 110000
rect 67178 109200 67234 110000
rect 79414 109200 79470 110000
rect 91650 109200 91706 110000
rect 103886 109200 103942 110000
rect 4250 0 4306 800
rect 12714 0 12770 800
rect 21178 0 21234 800
rect 29642 0 29698 800
rect 38106 0 38162 800
rect 46570 0 46626 800
rect 55034 0 55090 800
rect 63498 0 63554 800
rect 71962 0 72018 800
rect 80426 0 80482 800
rect 88890 0 88946 800
rect 97354 0 97410 800
rect 105818 0 105874 800
<< obsm2 >>
rect 1398 109144 6034 109290
rect 6202 109144 18178 109290
rect 18346 109144 30414 109290
rect 30582 109144 42650 109290
rect 42818 109144 54886 109290
rect 55054 109144 67122 109290
rect 67290 109144 79358 109290
rect 79526 109144 91594 109290
rect 91762 109144 103830 109290
rect 103998 109144 108266 109290
rect 1398 856 108266 109144
rect 1398 800 4194 856
rect 4362 800 12658 856
rect 12826 800 21122 856
rect 21290 800 29586 856
rect 29754 800 38050 856
rect 38218 800 46514 856
rect 46682 800 54978 856
rect 55146 800 63442 856
rect 63610 800 71906 856
rect 72074 800 80370 856
rect 80538 800 88834 856
rect 89002 800 97298 856
rect 97466 800 105762 856
rect 105930 800 108266 856
<< metal3 >>
rect 0 109080 800 109200
rect 0 107448 800 107568
rect 0 105816 800 105936
rect 0 104184 800 104304
rect 109200 102960 110000 103080
rect 0 102552 800 102672
rect 0 100920 800 101040
rect 0 99288 800 99408
rect 0 97656 800 97776
rect 0 96024 800 96144
rect 0 94392 800 94512
rect 0 92760 800 92880
rect 0 91128 800 91248
rect 0 89496 800 89616
rect 109200 89224 110000 89344
rect 0 87728 800 87848
rect 0 86096 800 86216
rect 0 84464 800 84584
rect 0 82832 800 82952
rect 0 81200 800 81320
rect 0 79568 800 79688
rect 0 77936 800 78056
rect 0 76304 800 76424
rect 109200 75488 110000 75608
rect 0 74672 800 74792
rect 0 73040 800 73160
rect 0 71408 800 71528
rect 0 69776 800 69896
rect 0 68144 800 68264
rect 0 66376 800 66496
rect 0 64744 800 64864
rect 0 63112 800 63232
rect 109200 61752 110000 61872
rect 0 61480 800 61600
rect 0 59848 800 59968
rect 0 58216 800 58336
rect 0 56584 800 56704
rect 0 54952 800 55072
rect 0 53320 800 53440
rect 0 51688 800 51808
rect 0 50056 800 50176
rect 0 48424 800 48544
rect 109200 48016 110000 48136
rect 0 46792 800 46912
rect 0 45160 800 45280
rect 0 43392 800 43512
rect 0 41760 800 41880
rect 0 40128 800 40248
rect 0 38496 800 38616
rect 0 36864 800 36984
rect 0 35232 800 35352
rect 109200 34280 110000 34400
rect 0 33600 800 33720
rect 0 31968 800 32088
rect 0 30336 800 30456
rect 0 28704 800 28824
rect 0 27072 800 27192
rect 0 25440 800 25560
rect 0 23808 800 23928
rect 0 22040 800 22160
rect 0 20408 800 20528
rect 109200 20544 110000 20664
rect 0 18776 800 18896
rect 0 17144 800 17264
rect 0 15512 800 15632
rect 0 13880 800 14000
rect 0 12248 800 12368
rect 0 10616 800 10736
rect 0 8984 800 9104
rect 0 7352 800 7472
rect 109200 6808 110000 6928
rect 0 5720 800 5840
rect 0 4088 800 4208
rect 0 2456 800 2576
rect 0 824 800 944
<< obsm3 >>
rect 880 109000 109200 109173
rect 800 107648 109200 109000
rect 880 107368 109200 107648
rect 800 106016 109200 107368
rect 880 105736 109200 106016
rect 800 104384 109200 105736
rect 880 104104 109200 104384
rect 800 103160 109200 104104
rect 800 102880 109120 103160
rect 800 102752 109200 102880
rect 880 102472 109200 102752
rect 800 101120 109200 102472
rect 880 100840 109200 101120
rect 800 99488 109200 100840
rect 880 99208 109200 99488
rect 800 97856 109200 99208
rect 880 97576 109200 97856
rect 800 96224 109200 97576
rect 880 95944 109200 96224
rect 800 94592 109200 95944
rect 880 94312 109200 94592
rect 800 92960 109200 94312
rect 880 92680 109200 92960
rect 800 91328 109200 92680
rect 880 91048 109200 91328
rect 800 89696 109200 91048
rect 880 89424 109200 89696
rect 880 89416 109120 89424
rect 800 89144 109120 89416
rect 800 87928 109200 89144
rect 880 87648 109200 87928
rect 800 86296 109200 87648
rect 880 86016 109200 86296
rect 800 84664 109200 86016
rect 880 84384 109200 84664
rect 800 83032 109200 84384
rect 880 82752 109200 83032
rect 800 81400 109200 82752
rect 880 81120 109200 81400
rect 800 79768 109200 81120
rect 880 79488 109200 79768
rect 800 78136 109200 79488
rect 880 77856 109200 78136
rect 800 76504 109200 77856
rect 880 76224 109200 76504
rect 800 75688 109200 76224
rect 800 75408 109120 75688
rect 800 74872 109200 75408
rect 880 74592 109200 74872
rect 800 73240 109200 74592
rect 880 72960 109200 73240
rect 800 71608 109200 72960
rect 880 71328 109200 71608
rect 800 69976 109200 71328
rect 880 69696 109200 69976
rect 800 68344 109200 69696
rect 880 68064 109200 68344
rect 800 66576 109200 68064
rect 880 66296 109200 66576
rect 800 64944 109200 66296
rect 880 64664 109200 64944
rect 800 63312 109200 64664
rect 880 63032 109200 63312
rect 800 61952 109200 63032
rect 800 61680 109120 61952
rect 880 61672 109120 61680
rect 880 61400 109200 61672
rect 800 60048 109200 61400
rect 880 59768 109200 60048
rect 800 58416 109200 59768
rect 880 58136 109200 58416
rect 800 56784 109200 58136
rect 880 56504 109200 56784
rect 800 55152 109200 56504
rect 880 54872 109200 55152
rect 800 53520 109200 54872
rect 880 53240 109200 53520
rect 800 51888 109200 53240
rect 880 51608 109200 51888
rect 800 50256 109200 51608
rect 880 49976 109200 50256
rect 800 48624 109200 49976
rect 880 48344 109200 48624
rect 800 48216 109200 48344
rect 800 47936 109120 48216
rect 800 46992 109200 47936
rect 880 46712 109200 46992
rect 800 45360 109200 46712
rect 880 45080 109200 45360
rect 800 43592 109200 45080
rect 880 43312 109200 43592
rect 800 41960 109200 43312
rect 880 41680 109200 41960
rect 800 40328 109200 41680
rect 880 40048 109200 40328
rect 800 38696 109200 40048
rect 880 38416 109200 38696
rect 800 37064 109200 38416
rect 880 36784 109200 37064
rect 800 35432 109200 36784
rect 880 35152 109200 35432
rect 800 34480 109200 35152
rect 800 34200 109120 34480
rect 800 33800 109200 34200
rect 880 33520 109200 33800
rect 800 32168 109200 33520
rect 880 31888 109200 32168
rect 800 30536 109200 31888
rect 880 30256 109200 30536
rect 800 28904 109200 30256
rect 880 28624 109200 28904
rect 800 27272 109200 28624
rect 880 26992 109200 27272
rect 800 25640 109200 26992
rect 880 25360 109200 25640
rect 800 24008 109200 25360
rect 880 23728 109200 24008
rect 800 22240 109200 23728
rect 880 21960 109200 22240
rect 800 20744 109200 21960
rect 800 20608 109120 20744
rect 880 20464 109120 20608
rect 880 20328 109200 20464
rect 800 18976 109200 20328
rect 880 18696 109200 18976
rect 800 17344 109200 18696
rect 880 17064 109200 17344
rect 800 15712 109200 17064
rect 880 15432 109200 15712
rect 800 14080 109200 15432
rect 880 13800 109200 14080
rect 800 12448 109200 13800
rect 880 12168 109200 12448
rect 800 10816 109200 12168
rect 880 10536 109200 10816
rect 800 9184 109200 10536
rect 880 8904 109200 9184
rect 800 7552 109200 8904
rect 880 7272 109200 7552
rect 800 7008 109200 7272
rect 800 6728 109120 7008
rect 800 5920 109200 6728
rect 880 5640 109200 5920
rect 800 4288 109200 5640
rect 880 4008 109200 4288
rect 800 2656 109200 4008
rect 880 2376 109200 2656
rect 800 1024 109200 2376
rect 880 851 109200 1024
<< metal4 >>
rect 4208 2128 4528 107760
rect 19568 2128 19888 107760
rect 34928 2128 35248 107760
rect 50288 2128 50608 107760
rect 65648 2128 65968 107760
rect 81008 2128 81328 107760
rect 96368 2128 96688 107760
<< obsm4 >>
rect 10179 2347 19488 91765
rect 19968 2347 34848 91765
rect 35328 2347 50208 91765
rect 50688 2347 60661 91765
<< labels >>
rlabel metal2 s 6090 109200 6146 110000 6 clock
port 1 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 io_ba_match
port 2 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 io_motor_gpio_pwm_high
port 3 nsew signal output
rlabel metal2 s 12714 0 12770 800 6 io_motor_gpio_pwm_high_en
port 4 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 io_motor_gpio_pwm_low
port 5 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 io_motor_gpio_pwm_low_en
port 6 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 io_motor_gpio_qei_ch_a
port 7 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 io_motor_gpio_qei_ch_b
port 8 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 io_motor_irq
port 9 nsew signal output
rlabel metal3 s 109200 6808 110000 6928 6 io_wbs_ack_o
port 10 nsew signal output
rlabel metal3 s 109200 20544 110000 20664 6 io_wbs_data_o[0]
port 11 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 io_wbs_data_o[10]
port 12 nsew signal output
rlabel metal2 s 63498 0 63554 800 6 io_wbs_data_o[11]
port 13 nsew signal output
rlabel metal2 s 42706 109200 42762 110000 6 io_wbs_data_o[12]
port 14 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 io_wbs_data_o[13]
port 15 nsew signal output
rlabel metal3 s 109200 102960 110000 103080 6 io_wbs_data_o[14]
port 16 nsew signal output
rlabel metal2 s 54942 109200 54998 110000 6 io_wbs_data_o[15]
port 17 nsew signal output
rlabel metal2 s 80426 0 80482 800 6 io_wbs_data_o[16]
port 18 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 io_wbs_data_o[17]
port 19 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 io_wbs_data_o[18]
port 20 nsew signal output
rlabel metal2 s 67178 109200 67234 110000 6 io_wbs_data_o[19]
port 21 nsew signal output
rlabel metal3 s 109200 34280 110000 34400 6 io_wbs_data_o[1]
port 22 nsew signal output
rlabel metal2 s 88890 0 88946 800 6 io_wbs_data_o[20]
port 23 nsew signal output
rlabel metal2 s 79414 109200 79470 110000 6 io_wbs_data_o[21]
port 24 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 io_wbs_data_o[22]
port 25 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 io_wbs_data_o[23]
port 26 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 io_wbs_data_o[24]
port 27 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 io_wbs_data_o[25]
port 28 nsew signal output
rlabel metal3 s 0 105816 800 105936 6 io_wbs_data_o[26]
port 29 nsew signal output
rlabel metal2 s 91650 109200 91706 110000 6 io_wbs_data_o[27]
port 30 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 io_wbs_data_o[28]
port 31 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 io_wbs_data_o[29]
port 32 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 io_wbs_data_o[2]
port 33 nsew signal output
rlabel metal2 s 103886 109200 103942 110000 6 io_wbs_data_o[30]
port 34 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 io_wbs_data_o[31]
port 35 nsew signal output
rlabel metal2 s 30470 109200 30526 110000 6 io_wbs_data_o[3]
port 36 nsew signal output
rlabel metal3 s 109200 48016 110000 48136 6 io_wbs_data_o[4]
port 37 nsew signal output
rlabel metal3 s 109200 61752 110000 61872 6 io_wbs_data_o[5]
port 38 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 io_wbs_data_o[6]
port 39 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 io_wbs_data_o[7]
port 40 nsew signal output
rlabel metal3 s 109200 75488 110000 75608 6 io_wbs_data_o[8]
port 41 nsew signal output
rlabel metal3 s 109200 89224 110000 89344 6 io_wbs_data_o[9]
port 42 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_wbs_m2s_addr[0]
port 43 nsew signal input
rlabel metal3 s 0 43392 800 43512 6 io_wbs_m2s_addr[10]
port 44 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 io_wbs_m2s_addr[11]
port 45 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 io_wbs_m2s_addr[12]
port 46 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 io_wbs_m2s_addr[13]
port 47 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 io_wbs_m2s_addr[14]
port 48 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 io_wbs_m2s_addr[15]
port 49 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 io_wbs_m2s_addr[1]
port 50 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 io_wbs_m2s_addr[2]
port 51 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 io_wbs_m2s_addr[3]
port 52 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 io_wbs_m2s_addr[4]
port 53 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 io_wbs_m2s_addr[5]
port 54 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 io_wbs_m2s_addr[6]
port 55 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 io_wbs_m2s_addr[7]
port 56 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 io_wbs_m2s_addr[8]
port 57 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 io_wbs_m2s_addr[9]
port 58 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 io_wbs_m2s_data[0]
port 59 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 io_wbs_m2s_data[10]
port 60 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 io_wbs_m2s_data[11]
port 61 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 io_wbs_m2s_data[12]
port 62 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 io_wbs_m2s_data[13]
port 63 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 io_wbs_m2s_data[14]
port 64 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 io_wbs_m2s_data[15]
port 65 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 io_wbs_m2s_data[16]
port 66 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 io_wbs_m2s_data[17]
port 67 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 io_wbs_m2s_data[18]
port 68 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 io_wbs_m2s_data[19]
port 69 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 io_wbs_m2s_data[1]
port 70 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 io_wbs_m2s_data[20]
port 71 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 io_wbs_m2s_data[21]
port 72 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 io_wbs_m2s_data[22]
port 73 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 io_wbs_m2s_data[23]
port 74 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 io_wbs_m2s_data[24]
port 75 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 io_wbs_m2s_data[25]
port 76 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 io_wbs_m2s_data[26]
port 77 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 io_wbs_m2s_data[27]
port 78 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 io_wbs_m2s_data[28]
port 79 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 io_wbs_m2s_data[29]
port 80 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 io_wbs_m2s_data[2]
port 81 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 io_wbs_m2s_data[30]
port 82 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 io_wbs_m2s_data[31]
port 83 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_wbs_m2s_data[3]
port 84 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 io_wbs_m2s_data[4]
port 85 nsew signal input
rlabel metal3 s 0 28704 800 28824 6 io_wbs_m2s_data[5]
port 86 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 io_wbs_m2s_data[6]
port 87 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 io_wbs_m2s_data[7]
port 88 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 io_wbs_m2s_data[8]
port 89 nsew signal input
rlabel metal3 s 0 41760 800 41880 6 io_wbs_m2s_data[9]
port 90 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 io_wbs_m2s_sel[0]
port 91 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 io_wbs_m2s_sel[1]
port 92 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 io_wbs_m2s_sel[2]
port 93 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 io_wbs_m2s_sel[3]
port 94 nsew signal input
rlabel metal3 s 0 824 800 944 6 io_wbs_m2s_stb
port 95 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 io_wbs_m2s_we
port 96 nsew signal input
rlabel metal2 s 18234 109200 18290 110000 6 reset
port 97 nsew signal input
rlabel metal4 s 4208 2128 4528 107760 6 vccd1
port 98 nsew power input
rlabel metal4 s 34928 2128 35248 107760 6 vccd1
port 98 nsew power input
rlabel metal4 s 65648 2128 65968 107760 6 vccd1
port 98 nsew power input
rlabel metal4 s 96368 2128 96688 107760 6 vccd1
port 98 nsew power input
rlabel metal4 s 19568 2128 19888 107760 6 vssd1
port 99 nsew ground input
rlabel metal4 s 50288 2128 50608 107760 6 vssd1
port 99 nsew ground input
rlabel metal4 s 81008 2128 81328 107760 6 vssd1
port 99 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 110000 110000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18336108
string GDS_FILE /home/ali112000/Desktop/mpw/UETRV-ECORE/openlane/Motor_Top/runs/Motor_Top/results/finishing/Motor_Top.magic.gds
string GDS_START 1104644
<< end >>

