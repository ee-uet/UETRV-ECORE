magic
tech sky130A
magscale 1 2
timestamp 1647720188
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 14 1844 199718 197668
<< metal2 >>
rect 1306 199200 1362 200000
rect 3238 199200 3294 200000
rect 4526 199200 4582 200000
rect 6458 199200 6514 200000
rect 8390 199200 8446 200000
rect 10322 199200 10378 200000
rect 11610 199200 11666 200000
rect 13542 199200 13598 200000
rect 15474 199200 15530 200000
rect 17406 199200 17462 200000
rect 18694 199200 18750 200000
rect 20626 199200 20682 200000
rect 22558 199200 22614 200000
rect 23846 199200 23902 200000
rect 25778 199200 25834 200000
rect 27710 199200 27766 200000
rect 29642 199200 29698 200000
rect 30930 199200 30986 200000
rect 32862 199200 32918 200000
rect 34794 199200 34850 200000
rect 36726 199200 36782 200000
rect 38014 199200 38070 200000
rect 39946 199200 40002 200000
rect 41878 199200 41934 200000
rect 43810 199200 43866 200000
rect 45098 199200 45154 200000
rect 47030 199200 47086 200000
rect 48962 199200 49018 200000
rect 50894 199200 50950 200000
rect 52182 199200 52238 200000
rect 54114 199200 54170 200000
rect 56046 199200 56102 200000
rect 57978 199200 58034 200000
rect 59266 199200 59322 200000
rect 61198 199200 61254 200000
rect 63130 199200 63186 200000
rect 65062 199200 65118 200000
rect 66350 199200 66406 200000
rect 68282 199200 68338 200000
rect 70214 199200 70270 200000
rect 72146 199200 72202 200000
rect 73434 199200 73490 200000
rect 75366 199200 75422 200000
rect 77298 199200 77354 200000
rect 79230 199200 79286 200000
rect 80518 199200 80574 200000
rect 82450 199200 82506 200000
rect 84382 199200 84438 200000
rect 86314 199200 86370 200000
rect 87602 199200 87658 200000
rect 89534 199200 89590 200000
rect 91466 199200 91522 200000
rect 93398 199200 93454 200000
rect 94686 199200 94742 200000
rect 96618 199200 96674 200000
rect 98550 199200 98606 200000
rect 99838 199200 99894 200000
rect 101770 199200 101826 200000
rect 103702 199200 103758 200000
rect 105634 199200 105690 200000
rect 106922 199200 106978 200000
rect 108854 199200 108910 200000
rect 110786 199200 110842 200000
rect 112718 199200 112774 200000
rect 114006 199200 114062 200000
rect 115938 199200 115994 200000
rect 117870 199200 117926 200000
rect 119802 199200 119858 200000
rect 121090 199200 121146 200000
rect 123022 199200 123078 200000
rect 124954 199200 125010 200000
rect 126886 199200 126942 200000
rect 128174 199200 128230 200000
rect 130106 199200 130162 200000
rect 132038 199200 132094 200000
rect 133970 199200 134026 200000
rect 135258 199200 135314 200000
rect 137190 199200 137246 200000
rect 139122 199200 139178 200000
rect 141054 199200 141110 200000
rect 142342 199200 142398 200000
rect 144274 199200 144330 200000
rect 146206 199200 146262 200000
rect 148138 199200 148194 200000
rect 149426 199200 149482 200000
rect 151358 199200 151414 200000
rect 153290 199200 153346 200000
rect 155222 199200 155278 200000
rect 156510 199200 156566 200000
rect 158442 199200 158498 200000
rect 160374 199200 160430 200000
rect 162306 199200 162362 200000
rect 163594 199200 163650 200000
rect 165526 199200 165582 200000
rect 167458 199200 167514 200000
rect 168746 199200 168802 200000
rect 170678 199200 170734 200000
rect 172610 199200 172666 200000
rect 174542 199200 174598 200000
rect 175830 199200 175886 200000
rect 177762 199200 177818 200000
rect 179694 199200 179750 200000
rect 181626 199200 181682 200000
rect 182914 199200 182970 200000
rect 184846 199200 184902 200000
rect 186778 199200 186834 200000
rect 188710 199200 188766 200000
rect 189998 199200 190054 200000
rect 191930 199200 191986 200000
rect 193862 199200 193918 200000
rect 195794 199200 195850 200000
rect 197082 199200 197138 200000
rect 199014 199200 199070 200000
rect 18 0 74 800
rect 1306 0 1362 800
rect 3238 0 3294 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 29642 0 29698 800
rect 31574 0 31630 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36726 0 36782 800
rect 38658 0 38714 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 48962 0 49018 800
rect 50894 0 50950 800
rect 52826 0 52882 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 57978 0 58034 800
rect 59910 0 59966 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 65062 0 65118 800
rect 66994 0 67050 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 72146 0 72202 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 77298 0 77354 800
rect 79230 0 79286 800
rect 81162 0 81218 800
rect 82450 0 82506 800
rect 84382 0 84438 800
rect 86314 0 86370 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 91466 0 91522 800
rect 93398 0 93454 800
rect 95330 0 95386 800
rect 96618 0 96674 800
rect 98550 0 98606 800
rect 100482 0 100538 800
rect 102414 0 102470 800
rect 103702 0 103758 800
rect 105634 0 105690 800
rect 107566 0 107622 800
rect 109498 0 109554 800
rect 110786 0 110842 800
rect 112718 0 112774 800
rect 114650 0 114706 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 119802 0 119858 800
rect 121734 0 121790 800
rect 123666 0 123722 800
rect 124954 0 125010 800
rect 126886 0 126942 800
rect 128818 0 128874 800
rect 130750 0 130806 800
rect 132038 0 132094 800
rect 133970 0 134026 800
rect 135902 0 135958 800
rect 137834 0 137890 800
rect 139122 0 139178 800
rect 141054 0 141110 800
rect 142986 0 143042 800
rect 144274 0 144330 800
rect 146206 0 146262 800
rect 148138 0 148194 800
rect 150070 0 150126 800
rect 151358 0 151414 800
rect 153290 0 153346 800
rect 155222 0 155278 800
rect 157154 0 157210 800
rect 158442 0 158498 800
rect 160374 0 160430 800
rect 162306 0 162362 800
rect 164238 0 164294 800
rect 165526 0 165582 800
rect 167458 0 167514 800
rect 169390 0 169446 800
rect 171322 0 171378 800
rect 172610 0 172666 800
rect 174542 0 174598 800
rect 176474 0 176530 800
rect 178406 0 178462 800
rect 179694 0 179750 800
rect 181626 0 181682 800
rect 183558 0 183614 800
rect 185490 0 185546 800
rect 186778 0 186834 800
rect 188710 0 188766 800
rect 190642 0 190698 800
rect 192574 0 192630 800
rect 193862 0 193918 800
rect 195794 0 195850 800
rect 197726 0 197782 800
rect 199658 0 199714 800
<< obsm2 >>
rect 20 199144 1250 199345
rect 1418 199144 3182 199345
rect 3350 199144 4470 199345
rect 4638 199144 6402 199345
rect 6570 199144 8334 199345
rect 8502 199144 10266 199345
rect 10434 199144 11554 199345
rect 11722 199144 13486 199345
rect 13654 199144 15418 199345
rect 15586 199144 17350 199345
rect 17518 199144 18638 199345
rect 18806 199144 20570 199345
rect 20738 199144 22502 199345
rect 22670 199144 23790 199345
rect 23958 199144 25722 199345
rect 25890 199144 27654 199345
rect 27822 199144 29586 199345
rect 29754 199144 30874 199345
rect 31042 199144 32806 199345
rect 32974 199144 34738 199345
rect 34906 199144 36670 199345
rect 36838 199144 37958 199345
rect 38126 199144 39890 199345
rect 40058 199144 41822 199345
rect 41990 199144 43754 199345
rect 43922 199144 45042 199345
rect 45210 199144 46974 199345
rect 47142 199144 48906 199345
rect 49074 199144 50838 199345
rect 51006 199144 52126 199345
rect 52294 199144 54058 199345
rect 54226 199144 55990 199345
rect 56158 199144 57922 199345
rect 58090 199144 59210 199345
rect 59378 199144 61142 199345
rect 61310 199144 63074 199345
rect 63242 199144 65006 199345
rect 65174 199144 66294 199345
rect 66462 199144 68226 199345
rect 68394 199144 70158 199345
rect 70326 199144 72090 199345
rect 72258 199144 73378 199345
rect 73546 199144 75310 199345
rect 75478 199144 77242 199345
rect 77410 199144 79174 199345
rect 79342 199144 80462 199345
rect 80630 199144 82394 199345
rect 82562 199144 84326 199345
rect 84494 199144 86258 199345
rect 86426 199144 87546 199345
rect 87714 199144 89478 199345
rect 89646 199144 91410 199345
rect 91578 199144 93342 199345
rect 93510 199144 94630 199345
rect 94798 199144 96562 199345
rect 96730 199144 98494 199345
rect 98662 199144 99782 199345
rect 99950 199144 101714 199345
rect 101882 199144 103646 199345
rect 103814 199144 105578 199345
rect 105746 199144 106866 199345
rect 107034 199144 108798 199345
rect 108966 199144 110730 199345
rect 110898 199144 112662 199345
rect 112830 199144 113950 199345
rect 114118 199144 115882 199345
rect 116050 199144 117814 199345
rect 117982 199144 119746 199345
rect 119914 199144 121034 199345
rect 121202 199144 122966 199345
rect 123134 199144 124898 199345
rect 125066 199144 126830 199345
rect 126998 199144 128118 199345
rect 128286 199144 130050 199345
rect 130218 199144 131982 199345
rect 132150 199144 133914 199345
rect 134082 199144 135202 199345
rect 135370 199144 137134 199345
rect 137302 199144 139066 199345
rect 139234 199144 140998 199345
rect 141166 199144 142286 199345
rect 142454 199144 144218 199345
rect 144386 199144 146150 199345
rect 146318 199144 148082 199345
rect 148250 199144 149370 199345
rect 149538 199144 151302 199345
rect 151470 199144 153234 199345
rect 153402 199144 155166 199345
rect 155334 199144 156454 199345
rect 156622 199144 158386 199345
rect 158554 199144 160318 199345
rect 160486 199144 162250 199345
rect 162418 199144 163538 199345
rect 163706 199144 165470 199345
rect 165638 199144 167402 199345
rect 167570 199144 168690 199345
rect 168858 199144 170622 199345
rect 170790 199144 172554 199345
rect 172722 199144 174486 199345
rect 174654 199144 175774 199345
rect 175942 199144 177706 199345
rect 177874 199144 179638 199345
rect 179806 199144 181570 199345
rect 181738 199144 182858 199345
rect 183026 199144 184790 199345
rect 184958 199144 186722 199345
rect 186890 199144 188654 199345
rect 188822 199144 189942 199345
rect 190110 199144 191874 199345
rect 192042 199144 193806 199345
rect 193974 199144 195738 199345
rect 195906 199144 197026 199345
rect 197194 199144 198958 199345
rect 199126 199144 199712 199345
rect 20 856 199712 199144
rect 130 711 1250 856
rect 1418 711 3182 856
rect 3350 711 5114 856
rect 5282 711 6402 856
rect 6570 711 8334 856
rect 8502 711 10266 856
rect 10434 711 12198 856
rect 12366 711 13486 856
rect 13654 711 15418 856
rect 15586 711 17350 856
rect 17518 711 19282 856
rect 19450 711 20570 856
rect 20738 711 22502 856
rect 22670 711 24434 856
rect 24602 711 26366 856
rect 26534 711 27654 856
rect 27822 711 29586 856
rect 29754 711 31518 856
rect 31686 711 33450 856
rect 33618 711 34738 856
rect 34906 711 36670 856
rect 36838 711 38602 856
rect 38770 711 40534 856
rect 40702 711 41822 856
rect 41990 711 43754 856
rect 43922 711 45686 856
rect 45854 711 47618 856
rect 47786 711 48906 856
rect 49074 711 50838 856
rect 51006 711 52770 856
rect 52938 711 54702 856
rect 54870 711 55990 856
rect 56158 711 57922 856
rect 58090 711 59854 856
rect 60022 711 61786 856
rect 61954 711 63074 856
rect 63242 711 65006 856
rect 65174 711 66938 856
rect 67106 711 68870 856
rect 69038 711 70158 856
rect 70326 711 72090 856
rect 72258 711 74022 856
rect 74190 711 75310 856
rect 75478 711 77242 856
rect 77410 711 79174 856
rect 79342 711 81106 856
rect 81274 711 82394 856
rect 82562 711 84326 856
rect 84494 711 86258 856
rect 86426 711 88190 856
rect 88358 711 89478 856
rect 89646 711 91410 856
rect 91578 711 93342 856
rect 93510 711 95274 856
rect 95442 711 96562 856
rect 96730 711 98494 856
rect 98662 711 100426 856
rect 100594 711 102358 856
rect 102526 711 103646 856
rect 103814 711 105578 856
rect 105746 711 107510 856
rect 107678 711 109442 856
rect 109610 711 110730 856
rect 110898 711 112662 856
rect 112830 711 114594 856
rect 114762 711 116526 856
rect 116694 711 117814 856
rect 117982 711 119746 856
rect 119914 711 121678 856
rect 121846 711 123610 856
rect 123778 711 124898 856
rect 125066 711 126830 856
rect 126998 711 128762 856
rect 128930 711 130694 856
rect 130862 711 131982 856
rect 132150 711 133914 856
rect 134082 711 135846 856
rect 136014 711 137778 856
rect 137946 711 139066 856
rect 139234 711 140998 856
rect 141166 711 142930 856
rect 143098 711 144218 856
rect 144386 711 146150 856
rect 146318 711 148082 856
rect 148250 711 150014 856
rect 150182 711 151302 856
rect 151470 711 153234 856
rect 153402 711 155166 856
rect 155334 711 157098 856
rect 157266 711 158386 856
rect 158554 711 160318 856
rect 160486 711 162250 856
rect 162418 711 164182 856
rect 164350 711 165470 856
rect 165638 711 167402 856
rect 167570 711 169334 856
rect 169502 711 171266 856
rect 171434 711 172554 856
rect 172722 711 174486 856
rect 174654 711 176418 856
rect 176586 711 178350 856
rect 178518 711 179638 856
rect 179806 711 181570 856
rect 181738 711 183502 856
rect 183670 711 185434 856
rect 185602 711 186722 856
rect 186890 711 188654 856
rect 188822 711 190586 856
rect 190754 711 192518 856
rect 192686 711 193806 856
rect 193974 711 195738 856
rect 195906 711 197670 856
rect 197838 711 199602 856
<< metal3 >>
rect 0 199248 800 199368
rect 199200 198568 200000 198688
rect 0 197208 800 197328
rect 199200 196528 200000 196648
rect 0 195848 800 195968
rect 199200 195168 200000 195288
rect 0 193808 800 193928
rect 199200 193128 200000 193248
rect 0 191768 800 191888
rect 199200 191088 200000 191208
rect 0 189728 800 189848
rect 199200 189048 200000 189168
rect 0 188368 800 188488
rect 199200 187688 200000 187808
rect 0 186328 800 186448
rect 199200 185648 200000 185768
rect 0 184288 800 184408
rect 199200 183608 200000 183728
rect 0 182248 800 182368
rect 199200 181568 200000 181688
rect 0 180888 800 181008
rect 199200 180208 200000 180328
rect 0 178848 800 178968
rect 199200 178168 200000 178288
rect 0 176808 800 176928
rect 199200 176128 200000 176248
rect 0 174768 800 174888
rect 199200 174088 200000 174208
rect 0 173408 800 173528
rect 199200 172728 200000 172848
rect 0 171368 800 171488
rect 199200 170688 200000 170808
rect 0 169328 800 169448
rect 199200 168648 200000 168768
rect 0 167288 800 167408
rect 199200 166608 200000 166728
rect 0 165928 800 166048
rect 199200 165248 200000 165368
rect 0 163888 800 164008
rect 199200 163208 200000 163328
rect 0 161848 800 161968
rect 199200 161168 200000 161288
rect 0 159808 800 159928
rect 199200 159808 200000 159928
rect 0 158448 800 158568
rect 199200 157768 200000 157888
rect 0 156408 800 156528
rect 199200 155728 200000 155848
rect 0 154368 800 154488
rect 199200 153688 200000 153808
rect 0 152328 800 152448
rect 199200 152328 200000 152448
rect 0 150968 800 151088
rect 199200 150288 200000 150408
rect 0 148928 800 149048
rect 199200 148248 200000 148368
rect 0 146888 800 147008
rect 199200 146208 200000 146328
rect 0 145528 800 145648
rect 199200 144848 200000 144968
rect 0 143488 800 143608
rect 199200 142808 200000 142928
rect 0 141448 800 141568
rect 199200 140768 200000 140888
rect 0 139408 800 139528
rect 199200 138728 200000 138848
rect 0 138048 800 138168
rect 199200 137368 200000 137488
rect 0 136008 800 136128
rect 199200 135328 200000 135448
rect 0 133968 800 134088
rect 199200 133288 200000 133408
rect 0 131928 800 132048
rect 199200 131248 200000 131368
rect 0 130568 800 130688
rect 199200 129888 200000 130008
rect 0 128528 800 128648
rect 199200 127848 200000 127968
rect 0 126488 800 126608
rect 199200 125808 200000 125928
rect 0 124448 800 124568
rect 199200 123768 200000 123888
rect 0 123088 800 123208
rect 199200 122408 200000 122528
rect 0 121048 800 121168
rect 199200 120368 200000 120488
rect 0 119008 800 119128
rect 199200 118328 200000 118448
rect 0 116968 800 117088
rect 199200 116288 200000 116408
rect 0 115608 800 115728
rect 199200 114928 200000 115048
rect 0 113568 800 113688
rect 199200 112888 200000 113008
rect 0 111528 800 111648
rect 199200 110848 200000 110968
rect 0 109488 800 109608
rect 199200 108808 200000 108928
rect 0 108128 800 108248
rect 199200 107448 200000 107568
rect 0 106088 800 106208
rect 199200 105408 200000 105528
rect 0 104048 800 104168
rect 199200 103368 200000 103488
rect 0 102008 800 102128
rect 199200 101328 200000 101448
rect 0 100648 800 100768
rect 199200 99968 200000 100088
rect 0 98608 800 98728
rect 199200 97928 200000 98048
rect 0 96568 800 96688
rect 199200 95888 200000 96008
rect 0 94528 800 94648
rect 199200 93848 200000 93968
rect 0 93168 800 93288
rect 199200 92488 200000 92608
rect 0 91128 800 91248
rect 199200 90448 200000 90568
rect 0 89088 800 89208
rect 199200 88408 200000 88528
rect 0 87048 800 87168
rect 199200 87048 200000 87168
rect 0 85688 800 85808
rect 199200 85008 200000 85128
rect 0 83648 800 83768
rect 199200 82968 200000 83088
rect 0 81608 800 81728
rect 199200 80928 200000 81048
rect 0 79568 800 79688
rect 199200 79568 200000 79688
rect 0 78208 800 78328
rect 199200 77528 200000 77648
rect 0 76168 800 76288
rect 199200 75488 200000 75608
rect 0 74128 800 74248
rect 199200 73448 200000 73568
rect 0 72768 800 72888
rect 199200 72088 200000 72208
rect 0 70728 800 70848
rect 199200 70048 200000 70168
rect 0 68688 800 68808
rect 199200 68008 200000 68128
rect 0 66648 800 66768
rect 199200 65968 200000 66088
rect 0 65288 800 65408
rect 199200 64608 200000 64728
rect 0 63248 800 63368
rect 199200 62568 200000 62688
rect 0 61208 800 61328
rect 199200 60528 200000 60648
rect 0 59168 800 59288
rect 199200 58488 200000 58608
rect 0 57808 800 57928
rect 199200 57128 200000 57248
rect 0 55768 800 55888
rect 199200 55088 200000 55208
rect 0 53728 800 53848
rect 199200 53048 200000 53168
rect 0 51688 800 51808
rect 199200 51008 200000 51128
rect 0 50328 800 50448
rect 199200 49648 200000 49768
rect 0 48288 800 48408
rect 199200 47608 200000 47728
rect 0 46248 800 46368
rect 199200 45568 200000 45688
rect 0 44208 800 44328
rect 199200 43528 200000 43648
rect 0 42848 800 42968
rect 199200 42168 200000 42288
rect 0 40808 800 40928
rect 199200 40128 200000 40248
rect 0 38768 800 38888
rect 199200 38088 200000 38208
rect 0 36728 800 36848
rect 199200 36048 200000 36168
rect 0 35368 800 35488
rect 199200 34688 200000 34808
rect 0 33328 800 33448
rect 199200 32648 200000 32768
rect 0 31288 800 31408
rect 199200 30608 200000 30728
rect 0 29248 800 29368
rect 199200 28568 200000 28688
rect 0 27888 800 28008
rect 199200 27208 200000 27328
rect 0 25848 800 25968
rect 199200 25168 200000 25288
rect 0 23808 800 23928
rect 199200 23128 200000 23248
rect 0 21768 800 21888
rect 199200 21088 200000 21208
rect 0 20408 800 20528
rect 199200 19728 200000 19848
rect 0 18368 800 18488
rect 199200 17688 200000 17808
rect 0 16328 800 16448
rect 199200 15648 200000 15768
rect 0 14288 800 14408
rect 199200 13608 200000 13728
rect 0 12928 800 13048
rect 199200 12248 200000 12368
rect 0 10888 800 11008
rect 199200 10208 200000 10328
rect 0 8848 800 8968
rect 199200 8168 200000 8288
rect 0 6808 800 6928
rect 199200 6808 200000 6928
rect 0 5448 800 5568
rect 199200 4768 200000 4888
rect 0 3408 800 3528
rect 199200 2728 200000 2848
rect 0 1368 800 1488
rect 199200 688 200000 808
<< obsm3 >>
rect 880 199168 199200 199341
rect 800 198768 199200 199168
rect 800 198488 199120 198768
rect 800 197408 199200 198488
rect 880 197128 199200 197408
rect 800 196728 199200 197128
rect 800 196448 199120 196728
rect 800 196048 199200 196448
rect 880 195768 199200 196048
rect 800 195368 199200 195768
rect 800 195088 199120 195368
rect 800 194008 199200 195088
rect 880 193728 199200 194008
rect 800 193328 199200 193728
rect 800 193048 199120 193328
rect 800 191968 199200 193048
rect 880 191688 199200 191968
rect 800 191288 199200 191688
rect 800 191008 199120 191288
rect 800 189928 199200 191008
rect 880 189648 199200 189928
rect 800 189248 199200 189648
rect 800 188968 199120 189248
rect 800 188568 199200 188968
rect 880 188288 199200 188568
rect 800 187888 199200 188288
rect 800 187608 199120 187888
rect 800 186528 199200 187608
rect 880 186248 199200 186528
rect 800 185848 199200 186248
rect 800 185568 199120 185848
rect 800 184488 199200 185568
rect 880 184208 199200 184488
rect 800 183808 199200 184208
rect 800 183528 199120 183808
rect 800 182448 199200 183528
rect 880 182168 199200 182448
rect 800 181768 199200 182168
rect 800 181488 199120 181768
rect 800 181088 199200 181488
rect 880 180808 199200 181088
rect 800 180408 199200 180808
rect 800 180128 199120 180408
rect 800 179048 199200 180128
rect 880 178768 199200 179048
rect 800 178368 199200 178768
rect 800 178088 199120 178368
rect 800 177008 199200 178088
rect 880 176728 199200 177008
rect 800 176328 199200 176728
rect 800 176048 199120 176328
rect 800 174968 199200 176048
rect 880 174688 199200 174968
rect 800 174288 199200 174688
rect 800 174008 199120 174288
rect 800 173608 199200 174008
rect 880 173328 199200 173608
rect 800 172928 199200 173328
rect 800 172648 199120 172928
rect 800 171568 199200 172648
rect 880 171288 199200 171568
rect 800 170888 199200 171288
rect 800 170608 199120 170888
rect 800 169528 199200 170608
rect 880 169248 199200 169528
rect 800 168848 199200 169248
rect 800 168568 199120 168848
rect 800 167488 199200 168568
rect 880 167208 199200 167488
rect 800 166808 199200 167208
rect 800 166528 199120 166808
rect 800 166128 199200 166528
rect 880 165848 199200 166128
rect 800 165448 199200 165848
rect 800 165168 199120 165448
rect 800 164088 199200 165168
rect 880 163808 199200 164088
rect 800 163408 199200 163808
rect 800 163128 199120 163408
rect 800 162048 199200 163128
rect 880 161768 199200 162048
rect 800 161368 199200 161768
rect 800 161088 199120 161368
rect 800 160008 199200 161088
rect 880 159728 199120 160008
rect 800 158648 199200 159728
rect 880 158368 199200 158648
rect 800 157968 199200 158368
rect 800 157688 199120 157968
rect 800 156608 199200 157688
rect 880 156328 199200 156608
rect 800 155928 199200 156328
rect 800 155648 199120 155928
rect 800 154568 199200 155648
rect 880 154288 199200 154568
rect 800 153888 199200 154288
rect 800 153608 199120 153888
rect 800 152528 199200 153608
rect 880 152248 199120 152528
rect 800 151168 199200 152248
rect 880 150888 199200 151168
rect 800 150488 199200 150888
rect 800 150208 199120 150488
rect 800 149128 199200 150208
rect 880 148848 199200 149128
rect 800 148448 199200 148848
rect 800 148168 199120 148448
rect 800 147088 199200 148168
rect 880 146808 199200 147088
rect 800 146408 199200 146808
rect 800 146128 199120 146408
rect 800 145728 199200 146128
rect 880 145448 199200 145728
rect 800 145048 199200 145448
rect 800 144768 199120 145048
rect 800 143688 199200 144768
rect 880 143408 199200 143688
rect 800 143008 199200 143408
rect 800 142728 199120 143008
rect 800 141648 199200 142728
rect 880 141368 199200 141648
rect 800 140968 199200 141368
rect 800 140688 199120 140968
rect 800 139608 199200 140688
rect 880 139328 199200 139608
rect 800 138928 199200 139328
rect 800 138648 199120 138928
rect 800 138248 199200 138648
rect 880 137968 199200 138248
rect 800 137568 199200 137968
rect 800 137288 199120 137568
rect 800 136208 199200 137288
rect 880 135928 199200 136208
rect 800 135528 199200 135928
rect 800 135248 199120 135528
rect 800 134168 199200 135248
rect 880 133888 199200 134168
rect 800 133488 199200 133888
rect 800 133208 199120 133488
rect 800 132128 199200 133208
rect 880 131848 199200 132128
rect 800 131448 199200 131848
rect 800 131168 199120 131448
rect 800 130768 199200 131168
rect 880 130488 199200 130768
rect 800 130088 199200 130488
rect 800 129808 199120 130088
rect 800 128728 199200 129808
rect 880 128448 199200 128728
rect 800 128048 199200 128448
rect 800 127768 199120 128048
rect 800 126688 199200 127768
rect 880 126408 199200 126688
rect 800 126008 199200 126408
rect 800 125728 199120 126008
rect 800 124648 199200 125728
rect 880 124368 199200 124648
rect 800 123968 199200 124368
rect 800 123688 199120 123968
rect 800 123288 199200 123688
rect 880 123008 199200 123288
rect 800 122608 199200 123008
rect 800 122328 199120 122608
rect 800 121248 199200 122328
rect 880 120968 199200 121248
rect 800 120568 199200 120968
rect 800 120288 199120 120568
rect 800 119208 199200 120288
rect 880 118928 199200 119208
rect 800 118528 199200 118928
rect 800 118248 199120 118528
rect 800 117168 199200 118248
rect 880 116888 199200 117168
rect 800 116488 199200 116888
rect 800 116208 199120 116488
rect 800 115808 199200 116208
rect 880 115528 199200 115808
rect 800 115128 199200 115528
rect 800 114848 199120 115128
rect 800 113768 199200 114848
rect 880 113488 199200 113768
rect 800 113088 199200 113488
rect 800 112808 199120 113088
rect 800 111728 199200 112808
rect 880 111448 199200 111728
rect 800 111048 199200 111448
rect 800 110768 199120 111048
rect 800 109688 199200 110768
rect 880 109408 199200 109688
rect 800 109008 199200 109408
rect 800 108728 199120 109008
rect 800 108328 199200 108728
rect 880 108048 199200 108328
rect 800 107648 199200 108048
rect 800 107368 199120 107648
rect 800 106288 199200 107368
rect 880 106008 199200 106288
rect 800 105608 199200 106008
rect 800 105328 199120 105608
rect 800 104248 199200 105328
rect 880 103968 199200 104248
rect 800 103568 199200 103968
rect 800 103288 199120 103568
rect 800 102208 199200 103288
rect 880 101928 199200 102208
rect 800 101528 199200 101928
rect 800 101248 199120 101528
rect 800 100848 199200 101248
rect 880 100568 199200 100848
rect 800 100168 199200 100568
rect 800 99888 199120 100168
rect 800 98808 199200 99888
rect 880 98528 199200 98808
rect 800 98128 199200 98528
rect 800 97848 199120 98128
rect 800 96768 199200 97848
rect 880 96488 199200 96768
rect 800 96088 199200 96488
rect 800 95808 199120 96088
rect 800 94728 199200 95808
rect 880 94448 199200 94728
rect 800 94048 199200 94448
rect 800 93768 199120 94048
rect 800 93368 199200 93768
rect 880 93088 199200 93368
rect 800 92688 199200 93088
rect 800 92408 199120 92688
rect 800 91328 199200 92408
rect 880 91048 199200 91328
rect 800 90648 199200 91048
rect 800 90368 199120 90648
rect 800 89288 199200 90368
rect 880 89008 199200 89288
rect 800 88608 199200 89008
rect 800 88328 199120 88608
rect 800 87248 199200 88328
rect 880 86968 199120 87248
rect 800 85888 199200 86968
rect 880 85608 199200 85888
rect 800 85208 199200 85608
rect 800 84928 199120 85208
rect 800 83848 199200 84928
rect 880 83568 199200 83848
rect 800 83168 199200 83568
rect 800 82888 199120 83168
rect 800 81808 199200 82888
rect 880 81528 199200 81808
rect 800 81128 199200 81528
rect 800 80848 199120 81128
rect 800 79768 199200 80848
rect 880 79488 199120 79768
rect 800 78408 199200 79488
rect 880 78128 199200 78408
rect 800 77728 199200 78128
rect 800 77448 199120 77728
rect 800 76368 199200 77448
rect 880 76088 199200 76368
rect 800 75688 199200 76088
rect 800 75408 199120 75688
rect 800 74328 199200 75408
rect 880 74048 199200 74328
rect 800 73648 199200 74048
rect 800 73368 199120 73648
rect 800 72968 199200 73368
rect 880 72688 199200 72968
rect 800 72288 199200 72688
rect 800 72008 199120 72288
rect 800 70928 199200 72008
rect 880 70648 199200 70928
rect 800 70248 199200 70648
rect 800 69968 199120 70248
rect 800 68888 199200 69968
rect 880 68608 199200 68888
rect 800 68208 199200 68608
rect 800 67928 199120 68208
rect 800 66848 199200 67928
rect 880 66568 199200 66848
rect 800 66168 199200 66568
rect 800 65888 199120 66168
rect 800 65488 199200 65888
rect 880 65208 199200 65488
rect 800 64808 199200 65208
rect 800 64528 199120 64808
rect 800 63448 199200 64528
rect 880 63168 199200 63448
rect 800 62768 199200 63168
rect 800 62488 199120 62768
rect 800 61408 199200 62488
rect 880 61128 199200 61408
rect 800 60728 199200 61128
rect 800 60448 199120 60728
rect 800 59368 199200 60448
rect 880 59088 199200 59368
rect 800 58688 199200 59088
rect 800 58408 199120 58688
rect 800 58008 199200 58408
rect 880 57728 199200 58008
rect 800 57328 199200 57728
rect 800 57048 199120 57328
rect 800 55968 199200 57048
rect 880 55688 199200 55968
rect 800 55288 199200 55688
rect 800 55008 199120 55288
rect 800 53928 199200 55008
rect 880 53648 199200 53928
rect 800 53248 199200 53648
rect 800 52968 199120 53248
rect 800 51888 199200 52968
rect 880 51608 199200 51888
rect 800 51208 199200 51608
rect 800 50928 199120 51208
rect 800 50528 199200 50928
rect 880 50248 199200 50528
rect 800 49848 199200 50248
rect 800 49568 199120 49848
rect 800 48488 199200 49568
rect 880 48208 199200 48488
rect 800 47808 199200 48208
rect 800 47528 199120 47808
rect 800 46448 199200 47528
rect 880 46168 199200 46448
rect 800 45768 199200 46168
rect 800 45488 199120 45768
rect 800 44408 199200 45488
rect 880 44128 199200 44408
rect 800 43728 199200 44128
rect 800 43448 199120 43728
rect 800 43048 199200 43448
rect 880 42768 199200 43048
rect 800 42368 199200 42768
rect 800 42088 199120 42368
rect 800 41008 199200 42088
rect 880 40728 199200 41008
rect 800 40328 199200 40728
rect 800 40048 199120 40328
rect 800 38968 199200 40048
rect 880 38688 199200 38968
rect 800 38288 199200 38688
rect 800 38008 199120 38288
rect 800 36928 199200 38008
rect 880 36648 199200 36928
rect 800 36248 199200 36648
rect 800 35968 199120 36248
rect 800 35568 199200 35968
rect 880 35288 199200 35568
rect 800 34888 199200 35288
rect 800 34608 199120 34888
rect 800 33528 199200 34608
rect 880 33248 199200 33528
rect 800 32848 199200 33248
rect 800 32568 199120 32848
rect 800 31488 199200 32568
rect 880 31208 199200 31488
rect 800 30808 199200 31208
rect 800 30528 199120 30808
rect 800 29448 199200 30528
rect 880 29168 199200 29448
rect 800 28768 199200 29168
rect 800 28488 199120 28768
rect 800 28088 199200 28488
rect 880 27808 199200 28088
rect 800 27408 199200 27808
rect 800 27128 199120 27408
rect 800 26048 199200 27128
rect 880 25768 199200 26048
rect 800 25368 199200 25768
rect 800 25088 199120 25368
rect 800 24008 199200 25088
rect 880 23728 199200 24008
rect 800 23328 199200 23728
rect 800 23048 199120 23328
rect 800 21968 199200 23048
rect 880 21688 199200 21968
rect 800 21288 199200 21688
rect 800 21008 199120 21288
rect 800 20608 199200 21008
rect 880 20328 199200 20608
rect 800 19928 199200 20328
rect 800 19648 199120 19928
rect 800 18568 199200 19648
rect 880 18288 199200 18568
rect 800 17888 199200 18288
rect 800 17608 199120 17888
rect 800 16528 199200 17608
rect 880 16248 199200 16528
rect 800 15848 199200 16248
rect 800 15568 199120 15848
rect 800 14488 199200 15568
rect 880 14208 199200 14488
rect 800 13808 199200 14208
rect 800 13528 199120 13808
rect 800 13128 199200 13528
rect 880 12848 199200 13128
rect 800 12448 199200 12848
rect 800 12168 199120 12448
rect 800 11088 199200 12168
rect 880 10808 199200 11088
rect 800 10408 199200 10808
rect 800 10128 199120 10408
rect 800 9048 199200 10128
rect 880 8768 199200 9048
rect 800 8368 199200 8768
rect 800 8088 199120 8368
rect 800 7008 199200 8088
rect 880 6728 199120 7008
rect 800 5648 199200 6728
rect 880 5368 199200 5648
rect 800 4968 199200 5368
rect 800 4688 199120 4968
rect 800 3608 199200 4688
rect 880 3328 199200 3608
rect 800 2928 199200 3328
rect 800 2648 199120 2928
rect 800 1568 199200 2648
rect 880 1288 199200 1568
rect 800 888 199200 1288
rect 800 715 199120 888
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< obsm4 >>
rect 80467 2483 80928 197165
rect 81408 2483 96288 197165
rect 96768 2483 111648 197165
rect 112128 2483 127008 197165
rect 127488 2483 137021 197165
<< labels >>
rlabel metal3 s 0 42848 800 42968 6 clock
port 1 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 io_dbus_addr[0]
port 2 nsew signal input
rlabel metal3 s 199200 13608 200000 13728 6 io_dbus_addr[10]
port 3 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 io_dbus_addr[11]
port 4 nsew signal input
rlabel metal2 s 128174 199200 128230 200000 6 io_dbus_addr[12]
port 5 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 io_dbus_addr[13]
port 6 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 io_dbus_addr[14]
port 7 nsew signal input
rlabel metal2 s 172610 0 172666 800 6 io_dbus_addr[15]
port 8 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 io_dbus_addr[16]
port 9 nsew signal input
rlabel metal2 s 183558 0 183614 800 6 io_dbus_addr[17]
port 10 nsew signal input
rlabel metal3 s 199200 170688 200000 170808 6 io_dbus_addr[18]
port 11 nsew signal input
rlabel metal2 s 3238 199200 3294 200000 6 io_dbus_addr[19]
port 12 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 io_dbus_addr[1]
port 13 nsew signal input
rlabel metal2 s 56046 199200 56102 200000 6 io_dbus_addr[20]
port 14 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 io_dbus_addr[21]
port 15 nsew signal input
rlabel metal2 s 115938 199200 115994 200000 6 io_dbus_addr[22]
port 16 nsew signal input
rlabel metal3 s 199200 93848 200000 93968 6 io_dbus_addr[23]
port 17 nsew signal input
rlabel metal3 s 199200 79568 200000 79688 6 io_dbus_addr[24]
port 18 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 io_dbus_addr[25]
port 19 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 io_dbus_addr[26]
port 20 nsew signal input
rlabel metal3 s 199200 193128 200000 193248 6 io_dbus_addr[27]
port 21 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 io_dbus_addr[28]
port 22 nsew signal input
rlabel metal3 s 199200 172728 200000 172848 6 io_dbus_addr[29]
port 23 nsew signal input
rlabel metal2 s 158442 199200 158498 200000 6 io_dbus_addr[2]
port 24 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_dbus_addr[30]
port 25 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_dbus_addr[31]
port 26 nsew signal input
rlabel metal2 s 135258 199200 135314 200000 6 io_dbus_addr[3]
port 27 nsew signal input
rlabel metal3 s 199200 114928 200000 115048 6 io_dbus_addr[4]
port 28 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 io_dbus_addr[5]
port 29 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 io_dbus_addr[6]
port 30 nsew signal input
rlabel metal2 s 18694 199200 18750 200000 6 io_dbus_addr[7]
port 31 nsew signal input
rlabel metal2 s 199014 199200 199070 200000 6 io_dbus_addr[8]
port 32 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 io_dbus_addr[9]
port 33 nsew signal input
rlabel metal2 s 174542 0 174598 800 6 io_dbus_ld_type[0]
port 34 nsew signal input
rlabel metal2 s 151358 199200 151414 200000 6 io_dbus_ld_type[1]
port 35 nsew signal input
rlabel metal2 s 189998 199200 190054 200000 6 io_dbus_ld_type[2]
port 36 nsew signal input
rlabel metal3 s 199200 80928 200000 81048 6 io_dbus_rd_en
port 37 nsew signal input
rlabel metal2 s 4526 199200 4582 200000 6 io_dbus_rdata[0]
port 38 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 io_dbus_rdata[10]
port 39 nsew signal output
rlabel metal2 s 160374 199200 160430 200000 6 io_dbus_rdata[11]
port 40 nsew signal output
rlabel metal2 s 94686 199200 94742 200000 6 io_dbus_rdata[12]
port 41 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_dbus_rdata[13]
port 42 nsew signal output
rlabel metal3 s 199200 49648 200000 49768 6 io_dbus_rdata[14]
port 43 nsew signal output
rlabel metal3 s 0 188368 800 188488 6 io_dbus_rdata[15]
port 44 nsew signal output
rlabel metal2 s 75366 199200 75422 200000 6 io_dbus_rdata[16]
port 45 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_dbus_rdata[17]
port 46 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 io_dbus_rdata[18]
port 47 nsew signal output
rlabel metal3 s 199200 65968 200000 66088 6 io_dbus_rdata[19]
port 48 nsew signal output
rlabel metal3 s 199200 142808 200000 142928 6 io_dbus_rdata[1]
port 49 nsew signal output
rlabel metal3 s 199200 195168 200000 195288 6 io_dbus_rdata[20]
port 50 nsew signal output
rlabel metal2 s 181626 0 181682 800 6 io_dbus_rdata[21]
port 51 nsew signal output
rlabel metal2 s 17406 199200 17462 200000 6 io_dbus_rdata[22]
port 52 nsew signal output
rlabel metal2 s 80518 199200 80574 200000 6 io_dbus_rdata[23]
port 53 nsew signal output
rlabel metal2 s 34794 199200 34850 200000 6 io_dbus_rdata[24]
port 54 nsew signal output
rlabel metal3 s 199200 198568 200000 198688 6 io_dbus_rdata[25]
port 55 nsew signal output
rlabel metal3 s 199200 23128 200000 23248 6 io_dbus_rdata[26]
port 56 nsew signal output
rlabel metal2 s 48962 199200 49018 200000 6 io_dbus_rdata[27]
port 57 nsew signal output
rlabel metal2 s 170678 199200 170734 200000 6 io_dbus_rdata[28]
port 58 nsew signal output
rlabel metal3 s 199200 148248 200000 148368 6 io_dbus_rdata[29]
port 59 nsew signal output
rlabel metal2 s 182914 199200 182970 200000 6 io_dbus_rdata[2]
port 60 nsew signal output
rlabel metal3 s 199200 68008 200000 68128 6 io_dbus_rdata[30]
port 61 nsew signal output
rlabel metal2 s 79230 199200 79286 200000 6 io_dbus_rdata[31]
port 62 nsew signal output
rlabel metal2 s 124954 199200 125010 200000 6 io_dbus_rdata[3]
port 63 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 io_dbus_rdata[4]
port 64 nsew signal output
rlabel metal3 s 199200 97928 200000 98048 6 io_dbus_rdata[5]
port 65 nsew signal output
rlabel metal2 s 41878 199200 41934 200000 6 io_dbus_rdata[6]
port 66 nsew signal output
rlabel metal2 s 15474 199200 15530 200000 6 io_dbus_rdata[7]
port 67 nsew signal output
rlabel metal2 s 77298 199200 77354 200000 6 io_dbus_rdata[8]
port 68 nsew signal output
rlabel metal2 s 175830 199200 175886 200000 6 io_dbus_rdata[9]
port 69 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 io_dbus_st_type[0]
port 70 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 io_dbus_st_type[1]
port 71 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 io_dbus_valid
port 72 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 io_dbus_wdata[0]
port 73 nsew signal input
rlabel metal2 s 193862 199200 193918 200000 6 io_dbus_wdata[10]
port 74 nsew signal input
rlabel metal3 s 199200 191088 200000 191208 6 io_dbus_wdata[11]
port 75 nsew signal input
rlabel metal3 s 199200 88408 200000 88528 6 io_dbus_wdata[12]
port 76 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 io_dbus_wdata[13]
port 77 nsew signal input
rlabel metal3 s 199200 165248 200000 165368 6 io_dbus_wdata[14]
port 78 nsew signal input
rlabel metal2 s 101770 199200 101826 200000 6 io_dbus_wdata[15]
port 79 nsew signal input
rlabel metal2 s 72146 199200 72202 200000 6 io_dbus_wdata[16]
port 80 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 io_dbus_wdata[17]
port 81 nsew signal input
rlabel metal2 s 119802 199200 119858 200000 6 io_dbus_wdata[18]
port 82 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_dbus_wdata[19]
port 83 nsew signal input
rlabel metal3 s 199200 155728 200000 155848 6 io_dbus_wdata[1]
port 84 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 io_dbus_wdata[20]
port 85 nsew signal input
rlabel metal3 s 199200 12248 200000 12368 6 io_dbus_wdata[21]
port 86 nsew signal input
rlabel metal2 s 106922 199200 106978 200000 6 io_dbus_wdata[22]
port 87 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 io_dbus_wdata[23]
port 88 nsew signal input
rlabel metal3 s 199200 688 200000 808 6 io_dbus_wdata[24]
port 89 nsew signal input
rlabel metal2 s 108854 199200 108910 200000 6 io_dbus_wdata[25]
port 90 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 io_dbus_wdata[26]
port 91 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 io_dbus_wdata[27]
port 92 nsew signal input
rlabel metal2 s 87602 199200 87658 200000 6 io_dbus_wdata[28]
port 93 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 io_dbus_wdata[29]
port 94 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 io_dbus_wdata[2]
port 95 nsew signal input
rlabel metal3 s 199200 28568 200000 28688 6 io_dbus_wdata[30]
port 96 nsew signal input
rlabel metal3 s 199200 51008 200000 51128 6 io_dbus_wdata[31]
port 97 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 io_dbus_wdata[3]
port 98 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 io_dbus_wdata[4]
port 99 nsew signal input
rlabel metal3 s 199200 73448 200000 73568 6 io_dbus_wdata[5]
port 100 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 io_dbus_wdata[6]
port 101 nsew signal input
rlabel metal3 s 0 163888 800 164008 6 io_dbus_wdata[7]
port 102 nsew signal input
rlabel metal3 s 199200 36048 200000 36168 6 io_dbus_wdata[8]
port 103 nsew signal input
rlabel metal3 s 199200 77528 200000 77648 6 io_dbus_wdata[9]
port 104 nsew signal input
rlabel metal2 s 141054 199200 141110 200000 6 io_dbus_wr_en
port 105 nsew signal input
rlabel metal3 s 199200 60528 200000 60648 6 io_dmem_io_addr[0]
port 106 nsew signal output
rlabel metal3 s 199200 42168 200000 42288 6 io_dmem_io_addr[1]
port 107 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 io_dmem_io_addr[2]
port 108 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 io_dmem_io_addr[3]
port 109 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 io_dmem_io_addr[4]
port 110 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 io_dmem_io_addr[5]
port 111 nsew signal output
rlabel metal3 s 199200 15648 200000 15768 6 io_dmem_io_addr[6]
port 112 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 io_dmem_io_addr[7]
port 113 nsew signal output
rlabel metal3 s 199200 43528 200000 43648 6 io_dmem_io_rdata[0]
port 114 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 io_dmem_io_rdata[10]
port 115 nsew signal input
rlabel metal3 s 199200 21088 200000 21208 6 io_dmem_io_rdata[11]
port 116 nsew signal input
rlabel metal2 s 172610 199200 172666 200000 6 io_dmem_io_rdata[12]
port 117 nsew signal input
rlabel metal3 s 199200 4768 200000 4888 6 io_dmem_io_rdata[13]
port 118 nsew signal input
rlabel metal3 s 199200 166608 200000 166728 6 io_dmem_io_rdata[14]
port 119 nsew signal input
rlabel metal2 s 32862 199200 32918 200000 6 io_dmem_io_rdata[15]
port 120 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 io_dmem_io_rdata[16]
port 121 nsew signal input
rlabel metal2 s 22558 199200 22614 200000 6 io_dmem_io_rdata[17]
port 122 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 io_dmem_io_rdata[18]
port 123 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 io_dmem_io_rdata[19]
port 124 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 io_dmem_io_rdata[1]
port 125 nsew signal input
rlabel metal3 s 199200 135328 200000 135448 6 io_dmem_io_rdata[20]
port 126 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 io_dmem_io_rdata[21]
port 127 nsew signal input
rlabel metal3 s 199200 108808 200000 108928 6 io_dmem_io_rdata[22]
port 128 nsew signal input
rlabel metal2 s 27710 199200 27766 200000 6 io_dmem_io_rdata[23]
port 129 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 io_dmem_io_rdata[24]
port 130 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 io_dmem_io_rdata[25]
port 131 nsew signal input
rlabel metal3 s 199200 40128 200000 40248 6 io_dmem_io_rdata[26]
port 132 nsew signal input
rlabel metal3 s 199200 32648 200000 32768 6 io_dmem_io_rdata[27]
port 133 nsew signal input
rlabel metal3 s 199200 58488 200000 58608 6 io_dmem_io_rdata[28]
port 134 nsew signal input
rlabel metal2 s 11610 199200 11666 200000 6 io_dmem_io_rdata[29]
port 135 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 io_dmem_io_rdata[2]
port 136 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 io_dmem_io_rdata[30]
port 137 nsew signal input
rlabel metal3 s 199200 176128 200000 176248 6 io_dmem_io_rdata[31]
port 138 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 io_dmem_io_rdata[3]
port 139 nsew signal input
rlabel metal2 s 112718 199200 112774 200000 6 io_dmem_io_rdata[4]
port 140 nsew signal input
rlabel metal3 s 199200 27208 200000 27328 6 io_dmem_io_rdata[5]
port 141 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 io_dmem_io_rdata[6]
port 142 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 io_dmem_io_rdata[7]
port 143 nsew signal input
rlabel metal2 s 68282 199200 68338 200000 6 io_dmem_io_rdata[8]
port 144 nsew signal input
rlabel metal2 s 70214 199200 70270 200000 6 io_dmem_io_rdata[9]
port 145 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 io_dmem_io_st_type[0]
port 146 nsew signal output
rlabel metal2 s 121090 199200 121146 200000 6 io_dmem_io_st_type[1]
port 147 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 io_dmem_io_st_type[2]
port 148 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 io_dmem_io_st_type[3]
port 149 nsew signal output
rlabel metal3 s 199200 161168 200000 161288 6 io_dmem_io_wdata[0]
port 150 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 io_dmem_io_wdata[10]
port 151 nsew signal output
rlabel metal3 s 199200 70048 200000 70168 6 io_dmem_io_wdata[11]
port 152 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_dmem_io_wdata[12]
port 153 nsew signal output
rlabel metal2 s 195794 199200 195850 200000 6 io_dmem_io_wdata[13]
port 154 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 io_dmem_io_wdata[14]
port 155 nsew signal output
rlabel metal2 s 195794 0 195850 800 6 io_dmem_io_wdata[15]
port 156 nsew signal output
rlabel metal2 s 137834 0 137890 800 6 io_dmem_io_wdata[16]
port 157 nsew signal output
rlabel metal2 s 193862 0 193918 800 6 io_dmem_io_wdata[17]
port 158 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 io_dmem_io_wdata[18]
port 159 nsew signal output
rlabel metal3 s 199200 157768 200000 157888 6 io_dmem_io_wdata[19]
port 160 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 io_dmem_io_wdata[1]
port 161 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 io_dmem_io_wdata[20]
port 162 nsew signal output
rlabel metal2 s 117870 199200 117926 200000 6 io_dmem_io_wdata[21]
port 163 nsew signal output
rlabel metal3 s 0 143488 800 143608 6 io_dmem_io_wdata[22]
port 164 nsew signal output
rlabel metal2 s 82450 199200 82506 200000 6 io_dmem_io_wdata[23]
port 165 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 io_dmem_io_wdata[24]
port 166 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 io_dmem_io_wdata[25]
port 167 nsew signal output
rlabel metal3 s 199200 168648 200000 168768 6 io_dmem_io_wdata[26]
port 168 nsew signal output
rlabel metal2 s 114006 199200 114062 200000 6 io_dmem_io_wdata[27]
port 169 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 io_dmem_io_wdata[28]
port 170 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 io_dmem_io_wdata[29]
port 171 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 io_dmem_io_wdata[2]
port 172 nsew signal output
rlabel metal3 s 199200 92488 200000 92608 6 io_dmem_io_wdata[30]
port 173 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_dmem_io_wdata[31]
port 174 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 io_dmem_io_wdata[3]
port 175 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 io_dmem_io_wdata[4]
port 176 nsew signal output
rlabel metal3 s 199200 150288 200000 150408 6 io_dmem_io_wdata[5]
port 177 nsew signal output
rlabel metal2 s 188710 199200 188766 200000 6 io_dmem_io_wdata[6]
port 178 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 io_dmem_io_wdata[7]
port 179 nsew signal output
rlabel metal2 s 65062 199200 65118 200000 6 io_dmem_io_wdata[8]
port 180 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 io_dmem_io_wdata[9]
port 181 nsew signal output
rlabel metal2 s 171322 0 171378 800 6 io_dmem_io_wr_en
port 182 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 io_ibus_addr[0]
port 183 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 io_ibus_addr[10]
port 184 nsew signal input
rlabel metal2 s 66350 199200 66406 200000 6 io_ibus_addr[11]
port 185 nsew signal input
rlabel metal2 s 98550 0 98606 800 6 io_ibus_addr[12]
port 186 nsew signal input
rlabel metal3 s 199200 87048 200000 87168 6 io_ibus_addr[13]
port 187 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 io_ibus_addr[14]
port 188 nsew signal input
rlabel metal3 s 199200 75488 200000 75608 6 io_ibus_addr[15]
port 189 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 io_ibus_addr[16]
port 190 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 io_ibus_addr[17]
port 191 nsew signal input
rlabel metal3 s 0 195848 800 195968 6 io_ibus_addr[18]
port 192 nsew signal input
rlabel metal2 s 45098 199200 45154 200000 6 io_ibus_addr[19]
port 193 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 io_ibus_addr[1]
port 194 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 io_ibus_addr[20]
port 195 nsew signal input
rlabel metal3 s 0 154368 800 154488 6 io_ibus_addr[21]
port 196 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 io_ibus_addr[22]
port 197 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 io_ibus_addr[23]
port 198 nsew signal input
rlabel metal3 s 199200 120368 200000 120488 6 io_ibus_addr[24]
port 199 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 io_ibus_addr[25]
port 200 nsew signal input
rlabel metal2 s 177762 199200 177818 200000 6 io_ibus_addr[26]
port 201 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 io_ibus_addr[27]
port 202 nsew signal input
rlabel metal2 s 192574 0 192630 800 6 io_ibus_addr[28]
port 203 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 io_ibus_addr[29]
port 204 nsew signal input
rlabel metal3 s 199200 127848 200000 127968 6 io_ibus_addr[2]
port 205 nsew signal input
rlabel metal2 s 1306 199200 1362 200000 6 io_ibus_addr[30]
port 206 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 io_ibus_addr[31]
port 207 nsew signal input
rlabel metal2 s 191930 199200 191986 200000 6 io_ibus_addr[3]
port 208 nsew signal input
rlabel metal3 s 199200 99968 200000 100088 6 io_ibus_addr[4]
port 209 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 io_ibus_addr[5]
port 210 nsew signal input
rlabel metal3 s 199200 129888 200000 130008 6 io_ibus_addr[6]
port 211 nsew signal input
rlabel metal2 s 52182 199200 52238 200000 6 io_ibus_addr[7]
port 212 nsew signal input
rlabel metal3 s 199200 189048 200000 189168 6 io_ibus_addr[8]
port 213 nsew signal input
rlabel metal3 s 0 184288 800 184408 6 io_ibus_addr[9]
port 214 nsew signal input
rlabel metal2 s 98550 199200 98606 200000 6 io_ibus_inst[0]
port 215 nsew signal output
rlabel metal3 s 199200 38088 200000 38208 6 io_ibus_inst[10]
port 216 nsew signal output
rlabel metal3 s 199200 163208 200000 163328 6 io_ibus_inst[11]
port 217 nsew signal output
rlabel metal3 s 199200 144848 200000 144968 6 io_ibus_inst[12]
port 218 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 io_ibus_inst[13]
port 219 nsew signal output
rlabel metal2 s 96618 199200 96674 200000 6 io_ibus_inst[14]
port 220 nsew signal output
rlabel metal2 s 146206 199200 146262 200000 6 io_ibus_inst[15]
port 221 nsew signal output
rlabel metal2 s 86314 199200 86370 200000 6 io_ibus_inst[16]
port 222 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_ibus_inst[17]
port 223 nsew signal output
rlabel metal2 s 59266 199200 59322 200000 6 io_ibus_inst[18]
port 224 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 io_ibus_inst[19]
port 225 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 io_ibus_inst[1]
port 226 nsew signal output
rlabel metal2 s 29642 199200 29698 200000 6 io_ibus_inst[20]
port 227 nsew signal output
rlabel metal2 s 148138 199200 148194 200000 6 io_ibus_inst[21]
port 228 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 io_ibus_inst[22]
port 229 nsew signal output
rlabel metal3 s 199200 47608 200000 47728 6 io_ibus_inst[23]
port 230 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 io_ibus_inst[24]
port 231 nsew signal output
rlabel metal2 s 91466 199200 91522 200000 6 io_ibus_inst[25]
port 232 nsew signal output
rlabel metal3 s 199200 181568 200000 181688 6 io_ibus_inst[26]
port 233 nsew signal output
rlabel metal3 s 199200 90448 200000 90568 6 io_ibus_inst[27]
port 234 nsew signal output
rlabel metal3 s 199200 10208 200000 10328 6 io_ibus_inst[28]
port 235 nsew signal output
rlabel metal3 s 0 197208 800 197328 6 io_ibus_inst[29]
port 236 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 io_ibus_inst[2]
port 237 nsew signal output
rlabel metal2 s 199658 0 199714 800 6 io_ibus_inst[30]
port 238 nsew signal output
rlabel metal3 s 0 193808 800 193928 6 io_ibus_inst[31]
port 239 nsew signal output
rlabel metal3 s 199200 187688 200000 187808 6 io_ibus_inst[3]
port 240 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 io_ibus_inst[4]
port 241 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 io_ibus_inst[5]
port 242 nsew signal output
rlabel metal2 s 103702 199200 103758 200000 6 io_ibus_inst[6]
port 243 nsew signal output
rlabel metal2 s 8390 199200 8446 200000 6 io_ibus_inst[7]
port 244 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 io_ibus_inst[8]
port 245 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 io_ibus_inst[9]
port 246 nsew signal output
rlabel metal3 s 0 161848 800 161968 6 io_ibus_valid
port 247 nsew signal output
rlabel metal3 s 199200 116288 200000 116408 6 io_imem_io_addr[0]
port 248 nsew signal output
rlabel metal3 s 199200 30608 200000 30728 6 io_imem_io_addr[10]
port 249 nsew signal output
rlabel metal3 s 0 186328 800 186448 6 io_imem_io_addr[11]
port 250 nsew signal output
rlabel metal3 s 199200 17688 200000 17808 6 io_imem_io_addr[12]
port 251 nsew signal output
rlabel metal2 s 13542 199200 13598 200000 6 io_imem_io_addr[13]
port 252 nsew signal output
rlabel metal2 s 137190 199200 137246 200000 6 io_imem_io_addr[14]
port 253 nsew signal output
rlabel metal3 s 0 156408 800 156528 6 io_imem_io_addr[15]
port 254 nsew signal output
rlabel metal3 s 199200 55088 200000 55208 6 io_imem_io_addr[16]
port 255 nsew signal output
rlabel metal2 s 93398 199200 93454 200000 6 io_imem_io_addr[17]
port 256 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 io_imem_io_addr[18]
port 257 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 io_imem_io_addr[19]
port 258 nsew signal output
rlabel metal2 s 89534 199200 89590 200000 6 io_imem_io_addr[1]
port 259 nsew signal output
rlabel metal2 s 144274 199200 144330 200000 6 io_imem_io_addr[20]
port 260 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 io_imem_io_addr[21]
port 261 nsew signal output
rlabel metal2 s 176474 0 176530 800 6 io_imem_io_addr[22]
port 262 nsew signal output
rlabel metal2 s 99838 199200 99894 200000 6 io_imem_io_addr[23]
port 263 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 io_imem_io_addr[24]
port 264 nsew signal output
rlabel metal2 s 174542 199200 174598 200000 6 io_imem_io_addr[25]
port 265 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 io_imem_io_addr[26]
port 266 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 io_imem_io_addr[27]
port 267 nsew signal output
rlabel metal3 s 199200 82968 200000 83088 6 io_imem_io_addr[28]
port 268 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 io_imem_io_addr[29]
port 269 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 io_imem_io_addr[2]
port 270 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 io_imem_io_addr[30]
port 271 nsew signal output
rlabel metal3 s 199200 125808 200000 125928 6 io_imem_io_addr[31]
port 272 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 io_imem_io_addr[3]
port 273 nsew signal output
rlabel metal2 s 178406 0 178462 800 6 io_imem_io_addr[4]
port 274 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 io_imem_io_addr[5]
port 275 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 io_imem_io_addr[6]
port 276 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 io_imem_io_addr[7]
port 277 nsew signal output
rlabel metal2 s 23846 199200 23902 200000 6 io_imem_io_addr[8]
port 278 nsew signal output
rlabel metal3 s 199200 110848 200000 110968 6 io_imem_io_addr[9]
port 279 nsew signal output
rlabel metal2 s 168746 199200 168802 200000 6 io_imem_io_rdata[0]
port 280 nsew signal input
rlabel metal2 s 162306 199200 162362 200000 6 io_imem_io_rdata[10]
port 281 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 io_imem_io_rdata[11]
port 282 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 io_imem_io_rdata[12]
port 283 nsew signal input
rlabel metal3 s 199200 131248 200000 131368 6 io_imem_io_rdata[13]
port 284 nsew signal input
rlabel metal2 s 179694 0 179750 800 6 io_imem_io_rdata[14]
port 285 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 io_imem_io_rdata[15]
port 286 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 io_imem_io_rdata[16]
port 287 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 io_imem_io_rdata[17]
port 288 nsew signal input
rlabel metal2 s 197082 199200 197138 200000 6 io_imem_io_rdata[18]
port 289 nsew signal input
rlabel metal2 s 184846 199200 184902 200000 6 io_imem_io_rdata[19]
port 290 nsew signal input
rlabel metal3 s 199200 183608 200000 183728 6 io_imem_io_rdata[1]
port 291 nsew signal input
rlabel metal2 s 73434 199200 73490 200000 6 io_imem_io_rdata[20]
port 292 nsew signal input
rlabel metal3 s 199200 174088 200000 174208 6 io_imem_io_rdata[21]
port 293 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 io_imem_io_rdata[22]
port 294 nsew signal input
rlabel metal2 s 165526 199200 165582 200000 6 io_imem_io_rdata[23]
port 295 nsew signal input
rlabel metal2 s 36726 199200 36782 200000 6 io_imem_io_rdata[24]
port 296 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 io_imem_io_rdata[25]
port 297 nsew signal input
rlabel metal2 s 38014 199200 38070 200000 6 io_imem_io_rdata[26]
port 298 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 io_imem_io_rdata[27]
port 299 nsew signal input
rlabel metal3 s 199200 8168 200000 8288 6 io_imem_io_rdata[28]
port 300 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_imem_io_rdata[29]
port 301 nsew signal input
rlabel metal3 s 199200 25168 200000 25288 6 io_imem_io_rdata[2]
port 302 nsew signal input
rlabel metal3 s 0 199248 800 199368 6 io_imem_io_rdata[30]
port 303 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 io_imem_io_rdata[31]
port 304 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 io_imem_io_rdata[3]
port 305 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 io_imem_io_rdata[4]
port 306 nsew signal input
rlabel metal2 s 155222 199200 155278 200000 6 io_imem_io_rdata[5]
port 307 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 io_imem_io_rdata[6]
port 308 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 io_imem_io_rdata[7]
port 309 nsew signal input
rlabel metal2 s 150070 0 150126 800 6 io_imem_io_rdata[8]
port 310 nsew signal input
rlabel metal3 s 199200 101328 200000 101448 6 io_imem_io_rdata[9]
port 311 nsew signal input
rlabel metal3 s 199200 140768 200000 140888 6 io_imem_io_wdata[0]
port 312 nsew signal output
rlabel metal3 s 0 145528 800 145648 6 io_imem_io_wdata[10]
port 313 nsew signal output
rlabel metal2 s 54114 199200 54170 200000 6 io_imem_io_wdata[11]
port 314 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 io_imem_io_wdata[12]
port 315 nsew signal output
rlabel metal3 s 199200 133288 200000 133408 6 io_imem_io_wdata[13]
port 316 nsew signal output
rlabel metal3 s 0 191768 800 191888 6 io_imem_io_wdata[14]
port 317 nsew signal output
rlabel metal3 s 199200 107448 200000 107568 6 io_imem_io_wdata[15]
port 318 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 io_imem_io_wdata[16]
port 319 nsew signal output
rlabel metal2 s 167458 199200 167514 200000 6 io_imem_io_wdata[17]
port 320 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 io_imem_io_wdata[18]
port 321 nsew signal output
rlabel metal2 s 110786 199200 110842 200000 6 io_imem_io_wdata[19]
port 322 nsew signal output
rlabel metal2 s 185490 0 185546 800 6 io_imem_io_wdata[1]
port 323 nsew signal output
rlabel metal2 s 39946 199200 40002 200000 6 io_imem_io_wdata[20]
port 324 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 io_imem_io_wdata[21]
port 325 nsew signal output
rlabel metal3 s 199200 103368 200000 103488 6 io_imem_io_wdata[22]
port 326 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 io_imem_io_wdata[23]
port 327 nsew signal output
rlabel metal3 s 199200 137368 200000 137488 6 io_imem_io_wdata[24]
port 328 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 io_imem_io_wdata[25]
port 329 nsew signal output
rlabel metal2 s 188710 0 188766 800 6 io_imem_io_wdata[26]
port 330 nsew signal output
rlabel metal2 s 50894 199200 50950 200000 6 io_imem_io_wdata[27]
port 331 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 io_imem_io_wdata[28]
port 332 nsew signal output
rlabel metal3 s 0 102008 800 102128 6 io_imem_io_wdata[29]
port 333 nsew signal output
rlabel metal2 s 43810 199200 43866 200000 6 io_imem_io_wdata[2]
port 334 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 io_imem_io_wdata[30]
port 335 nsew signal output
rlabel metal3 s 199200 34688 200000 34808 6 io_imem_io_wdata[31]
port 336 nsew signal output
rlabel metal2 s 30930 199200 30986 200000 6 io_imem_io_wdata[3]
port 337 nsew signal output
rlabel metal3 s 199200 72088 200000 72208 6 io_imem_io_wdata[4]
port 338 nsew signal output
rlabel metal2 s 126886 199200 126942 200000 6 io_imem_io_wdata[5]
port 339 nsew signal output
rlabel metal2 s 84382 199200 84438 200000 6 io_imem_io_wdata[6]
port 340 nsew signal output
rlabel metal2 s 6458 199200 6514 200000 6 io_imem_io_wdata[7]
port 341 nsew signal output
rlabel metal2 s 17406 0 17462 800 6 io_imem_io_wdata[8]
port 342 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 io_imem_io_wdata[9]
port 343 nsew signal output
rlabel metal3 s 199200 152328 200000 152448 6 io_imem_io_wr_en
port 344 nsew signal output
rlabel metal3 s 199200 138728 200000 138848 6 io_motor_ack_i
port 345 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 io_motor_addr_sel
port 346 nsew signal output
rlabel metal3 s 199200 123768 200000 123888 6 io_motor_data_i[0]
port 347 nsew signal input
rlabel metal3 s 199200 62568 200000 62688 6 io_motor_data_i[10]
port 348 nsew signal input
rlabel metal2 s 190642 0 190698 800 6 io_motor_data_i[11]
port 349 nsew signal input
rlabel metal2 s 123022 199200 123078 200000 6 io_motor_data_i[12]
port 350 nsew signal input
rlabel metal2 s 179694 199200 179750 200000 6 io_motor_data_i[13]
port 351 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 io_motor_data_i[14]
port 352 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 io_motor_data_i[15]
port 353 nsew signal input
rlabel metal3 s 199200 45568 200000 45688 6 io_motor_data_i[16]
port 354 nsew signal input
rlabel metal2 s 20626 199200 20682 200000 6 io_motor_data_i[17]
port 355 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 io_motor_data_i[18]
port 356 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 io_motor_data_i[19]
port 357 nsew signal input
rlabel metal2 s 63130 199200 63186 200000 6 io_motor_data_i[1]
port 358 nsew signal input
rlabel metal3 s 199200 118328 200000 118448 6 io_motor_data_i[20]
port 359 nsew signal input
rlabel metal3 s 199200 196528 200000 196648 6 io_motor_data_i[21]
port 360 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 io_motor_data_i[22]
port 361 nsew signal input
rlabel metal2 s 153290 199200 153346 200000 6 io_motor_data_i[23]
port 362 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 io_motor_data_i[24]
port 363 nsew signal input
rlabel metal2 s 153290 0 153346 800 6 io_motor_data_i[25]
port 364 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 io_motor_data_i[26]
port 365 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 io_motor_data_i[27]
port 366 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 io_motor_data_i[28]
port 367 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_motor_data_i[29]
port 368 nsew signal input
rlabel metal2 s 197726 0 197782 800 6 io_motor_data_i[2]
port 369 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 io_motor_data_i[30]
port 370 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_motor_data_i[31]
port 371 nsew signal input
rlabel metal3 s 199200 178168 200000 178288 6 io_motor_data_i[3]
port 372 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 io_motor_data_i[4]
port 373 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 io_motor_data_i[5]
port 374 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 io_motor_data_i[6]
port 375 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_motor_data_i[7]
port 376 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 io_motor_data_i[8]
port 377 nsew signal input
rlabel metal3 s 199200 105408 200000 105528 6 io_motor_data_i[9]
port 378 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 io_spi_clk
port 379 nsew signal output
rlabel metal2 s 133970 199200 134026 200000 6 io_spi_cs
port 380 nsew signal output
rlabel metal2 s 181626 199200 181682 200000 6 io_spi_irq
port 381 nsew signal output
rlabel metal2 s 10322 199200 10378 200000 6 io_spi_miso
port 382 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 io_spi_mosi
port 383 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 io_uart_irq
port 384 nsew signal output
rlabel metal2 s 186778 199200 186834 200000 6 io_uart_rx
port 385 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 io_uart_tx
port 386 nsew signal output
rlabel metal3 s 199200 159808 200000 159928 6 io_wbm_m2s_addr[0]
port 387 nsew signal output
rlabel metal3 s 199200 64608 200000 64728 6 io_wbm_m2s_addr[10]
port 388 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 io_wbm_m2s_addr[11]
port 389 nsew signal output
rlabel metal2 s 163594 199200 163650 200000 6 io_wbm_m2s_addr[12]
port 390 nsew signal output
rlabel metal2 s 47030 199200 47086 200000 6 io_wbm_m2s_addr[13]
port 391 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 io_wbm_m2s_addr[14]
port 392 nsew signal output
rlabel metal3 s 199200 122408 200000 122528 6 io_wbm_m2s_addr[15]
port 393 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 io_wbm_m2s_addr[1]
port 394 nsew signal output
rlabel metal3 s 199200 57128 200000 57248 6 io_wbm_m2s_addr[2]
port 395 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 io_wbm_m2s_addr[3]
port 396 nsew signal output
rlabel metal3 s 199200 2728 200000 2848 6 io_wbm_m2s_addr[4]
port 397 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 io_wbm_m2s_addr[5]
port 398 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 io_wbm_m2s_addr[6]
port 399 nsew signal output
rlabel metal3 s 199200 85008 200000 85128 6 io_wbm_m2s_addr[7]
port 400 nsew signal output
rlabel metal2 s 156510 199200 156566 200000 6 io_wbm_m2s_addr[8]
port 401 nsew signal output
rlabel metal3 s 199200 180208 200000 180328 6 io_wbm_m2s_addr[9]
port 402 nsew signal output
rlabel metal3 s 199200 6808 200000 6928 6 io_wbm_m2s_data[0]
port 403 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 io_wbm_m2s_data[10]
port 404 nsew signal output
rlabel metal3 s 199200 112888 200000 113008 6 io_wbm_m2s_data[11]
port 405 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 io_wbm_m2s_data[12]
port 406 nsew signal output
rlabel metal3 s 199200 185648 200000 185768 6 io_wbm_m2s_data[13]
port 407 nsew signal output
rlabel metal2 s 149426 199200 149482 200000 6 io_wbm_m2s_data[14]
port 408 nsew signal output
rlabel metal3 s 199200 19728 200000 19848 6 io_wbm_m2s_data[15]
port 409 nsew signal output
rlabel metal2 s 142342 199200 142398 200000 6 io_wbm_m2s_data[16]
port 410 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 io_wbm_m2s_data[17]
port 411 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 io_wbm_m2s_data[18]
port 412 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 io_wbm_m2s_data[19]
port 413 nsew signal output
rlabel metal2 s 18 0 74 800 6 io_wbm_m2s_data[1]
port 414 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 io_wbm_m2s_data[20]
port 415 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 io_wbm_m2s_data[21]
port 416 nsew signal output
rlabel metal3 s 0 174768 800 174888 6 io_wbm_m2s_data[22]
port 417 nsew signal output
rlabel metal2 s 57978 199200 58034 200000 6 io_wbm_m2s_data[23]
port 418 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 io_wbm_m2s_data[24]
port 419 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 io_wbm_m2s_data[25]
port 420 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 io_wbm_m2s_data[26]
port 421 nsew signal output
rlabel metal2 s 105634 199200 105690 200000 6 io_wbm_m2s_data[27]
port 422 nsew signal output
rlabel metal2 s 61198 199200 61254 200000 6 io_wbm_m2s_data[28]
port 423 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 io_wbm_m2s_data[29]
port 424 nsew signal output
rlabel metal2 s 139122 199200 139178 200000 6 io_wbm_m2s_data[2]
port 425 nsew signal output
rlabel metal3 s 199200 53048 200000 53168 6 io_wbm_m2s_data[30]
port 426 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 io_wbm_m2s_data[31]
port 427 nsew signal output
rlabel metal3 s 199200 153688 200000 153808 6 io_wbm_m2s_data[3]
port 428 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 io_wbm_m2s_data[4]
port 429 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 io_wbm_m2s_data[5]
port 430 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 io_wbm_m2s_data[6]
port 431 nsew signal output
rlabel metal3 s 199200 146208 200000 146328 6 io_wbm_m2s_data[7]
port 432 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 io_wbm_m2s_data[8]
port 433 nsew signal output
rlabel metal2 s 132038 199200 132094 200000 6 io_wbm_m2s_data[9]
port 434 nsew signal output
rlabel metal2 s 130106 199200 130162 200000 6 io_wbm_m2s_sel[0]
port 435 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 io_wbm_m2s_sel[1]
port 436 nsew signal output
rlabel metal2 s 25778 199200 25834 200000 6 io_wbm_m2s_sel[2]
port 437 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 io_wbm_m2s_sel[3]
port 438 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 io_wbm_m2s_stb
port 439 nsew signal output
rlabel metal3 s 0 169328 800 169448 6 io_wbm_m2s_we
port 440 nsew signal output
rlabel metal3 s 199200 95888 200000 96008 6 reset
port 441 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 442 nsew power input
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 442 nsew power input
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 442 nsew power input
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 442 nsew power input
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 442 nsew power input
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 442 nsew power input
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 442 nsew power input
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 443 nsew ground input
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 443 nsew ground input
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 443 nsew ground input
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 443 nsew ground input
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 443 nsew ground input
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 443 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 20137934
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Wishbone_InterConnect/runs/Wishbone_InterConnect/results/finishing/WB_InterConnect.magic.gds
string GDS_START 849388
<< end >>

