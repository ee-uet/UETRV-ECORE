magic
tech sky130A
magscale 1 2
timestamp 1647753841
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 14 1844 139826 138032
<< metal2 >>
rect 662 139200 718 140000
rect 1950 139200 2006 140000
rect 3238 139200 3294 140000
rect 5170 139200 5226 140000
rect 6458 139200 6514 140000
rect 7746 139200 7802 140000
rect 9034 139200 9090 140000
rect 10322 139200 10378 140000
rect 11610 139200 11666 140000
rect 12898 139200 12954 140000
rect 14186 139200 14242 140000
rect 15474 139200 15530 140000
rect 16762 139200 16818 140000
rect 18050 139200 18106 140000
rect 19338 139200 19394 140000
rect 20626 139200 20682 140000
rect 21914 139200 21970 140000
rect 23202 139200 23258 140000
rect 24490 139200 24546 140000
rect 25778 139200 25834 140000
rect 27066 139200 27122 140000
rect 28354 139200 28410 140000
rect 29642 139200 29698 140000
rect 30930 139200 30986 140000
rect 32218 139200 32274 140000
rect 33506 139200 33562 140000
rect 34794 139200 34850 140000
rect 36082 139200 36138 140000
rect 37370 139200 37426 140000
rect 38658 139200 38714 140000
rect 39946 139200 40002 140000
rect 41234 139200 41290 140000
rect 42522 139200 42578 140000
rect 43810 139200 43866 140000
rect 45098 139200 45154 140000
rect 46386 139200 46442 140000
rect 47674 139200 47730 140000
rect 48962 139200 49018 140000
rect 50250 139200 50306 140000
rect 51538 139200 51594 140000
rect 52826 139200 52882 140000
rect 54114 139200 54170 140000
rect 55402 139200 55458 140000
rect 56690 139200 56746 140000
rect 57978 139200 58034 140000
rect 59266 139200 59322 140000
rect 60554 139200 60610 140000
rect 61842 139200 61898 140000
rect 63130 139200 63186 140000
rect 64418 139200 64474 140000
rect 65706 139200 65762 140000
rect 66994 139200 67050 140000
rect 68282 139200 68338 140000
rect 69570 139200 69626 140000
rect 70858 139200 70914 140000
rect 72790 139200 72846 140000
rect 74078 139200 74134 140000
rect 75366 139200 75422 140000
rect 76654 139200 76710 140000
rect 77942 139200 77998 140000
rect 79230 139200 79286 140000
rect 80518 139200 80574 140000
rect 81806 139200 81862 140000
rect 83094 139200 83150 140000
rect 84382 139200 84438 140000
rect 85670 139200 85726 140000
rect 86958 139200 87014 140000
rect 88246 139200 88302 140000
rect 89534 139200 89590 140000
rect 90822 139200 90878 140000
rect 92110 139200 92166 140000
rect 93398 139200 93454 140000
rect 94686 139200 94742 140000
rect 95974 139200 96030 140000
rect 97262 139200 97318 140000
rect 98550 139200 98606 140000
rect 99838 139200 99894 140000
rect 101126 139200 101182 140000
rect 102414 139200 102470 140000
rect 103702 139200 103758 140000
rect 104990 139200 105046 140000
rect 106278 139200 106334 140000
rect 107566 139200 107622 140000
rect 108854 139200 108910 140000
rect 110142 139200 110198 140000
rect 111430 139200 111486 140000
rect 112718 139200 112774 140000
rect 114006 139200 114062 140000
rect 115294 139200 115350 140000
rect 116582 139200 116638 140000
rect 117870 139200 117926 140000
rect 119158 139200 119214 140000
rect 120446 139200 120502 140000
rect 121734 139200 121790 140000
rect 123022 139200 123078 140000
rect 124310 139200 124366 140000
rect 125598 139200 125654 140000
rect 126886 139200 126942 140000
rect 128174 139200 128230 140000
rect 129462 139200 129518 140000
rect 130750 139200 130806 140000
rect 132038 139200 132094 140000
rect 133326 139200 133382 140000
rect 134614 139200 134670 140000
rect 135902 139200 135958 140000
rect 137190 139200 137246 140000
rect 138478 139200 138534 140000
rect 139766 139200 139822 140000
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 32218 0 32274 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 42522 0 42578 800
rect 43810 0 43866 800
rect 45098 0 45154 800
rect 46386 0 46442 800
rect 47674 0 47730 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 54114 0 54170 800
rect 55402 0 55458 800
rect 56690 0 56746 800
rect 57978 0 58034 800
rect 59266 0 59322 800
rect 60554 0 60610 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66994 0 67050 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 77942 0 77998 800
rect 79230 0 79286 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 83094 0 83150 800
rect 84382 0 84438 800
rect 85670 0 85726 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 90822 0 90878 800
rect 92110 0 92166 800
rect 93398 0 93454 800
rect 94686 0 94742 800
rect 95974 0 96030 800
rect 97262 0 97318 800
rect 98550 0 98606 800
rect 99838 0 99894 800
rect 101126 0 101182 800
rect 102414 0 102470 800
rect 103702 0 103758 800
rect 104990 0 105046 800
rect 106278 0 106334 800
rect 107566 0 107622 800
rect 108854 0 108910 800
rect 110142 0 110198 800
rect 111430 0 111486 800
rect 112718 0 112774 800
rect 114006 0 114062 800
rect 115294 0 115350 800
rect 116582 0 116638 800
rect 117870 0 117926 800
rect 119158 0 119214 800
rect 120446 0 120502 800
rect 121734 0 121790 800
rect 123022 0 123078 800
rect 124310 0 124366 800
rect 125598 0 125654 800
rect 126886 0 126942 800
rect 128174 0 128230 800
rect 129462 0 129518 800
rect 130750 0 130806 800
rect 132038 0 132094 800
rect 133326 0 133382 800
rect 134614 0 134670 800
rect 136546 0 136602 800
rect 137834 0 137890 800
rect 139122 0 139178 800
<< obsm2 >>
rect 20 139144 606 139505
rect 774 139144 1894 139505
rect 2062 139144 3182 139505
rect 3350 139144 5114 139505
rect 5282 139144 6402 139505
rect 6570 139144 7690 139505
rect 7858 139144 8978 139505
rect 9146 139144 10266 139505
rect 10434 139144 11554 139505
rect 11722 139144 12842 139505
rect 13010 139144 14130 139505
rect 14298 139144 15418 139505
rect 15586 139144 16706 139505
rect 16874 139144 17994 139505
rect 18162 139144 19282 139505
rect 19450 139144 20570 139505
rect 20738 139144 21858 139505
rect 22026 139144 23146 139505
rect 23314 139144 24434 139505
rect 24602 139144 25722 139505
rect 25890 139144 27010 139505
rect 27178 139144 28298 139505
rect 28466 139144 29586 139505
rect 29754 139144 30874 139505
rect 31042 139144 32162 139505
rect 32330 139144 33450 139505
rect 33618 139144 34738 139505
rect 34906 139144 36026 139505
rect 36194 139144 37314 139505
rect 37482 139144 38602 139505
rect 38770 139144 39890 139505
rect 40058 139144 41178 139505
rect 41346 139144 42466 139505
rect 42634 139144 43754 139505
rect 43922 139144 45042 139505
rect 45210 139144 46330 139505
rect 46498 139144 47618 139505
rect 47786 139144 48906 139505
rect 49074 139144 50194 139505
rect 50362 139144 51482 139505
rect 51650 139144 52770 139505
rect 52938 139144 54058 139505
rect 54226 139144 55346 139505
rect 55514 139144 56634 139505
rect 56802 139144 57922 139505
rect 58090 139144 59210 139505
rect 59378 139144 60498 139505
rect 60666 139144 61786 139505
rect 61954 139144 63074 139505
rect 63242 139144 64362 139505
rect 64530 139144 65650 139505
rect 65818 139144 66938 139505
rect 67106 139144 68226 139505
rect 68394 139144 69514 139505
rect 69682 139144 70802 139505
rect 70970 139144 72734 139505
rect 72902 139144 74022 139505
rect 74190 139144 75310 139505
rect 75478 139144 76598 139505
rect 76766 139144 77886 139505
rect 78054 139144 79174 139505
rect 79342 139144 80462 139505
rect 80630 139144 81750 139505
rect 81918 139144 83038 139505
rect 83206 139144 84326 139505
rect 84494 139144 85614 139505
rect 85782 139144 86902 139505
rect 87070 139144 88190 139505
rect 88358 139144 89478 139505
rect 89646 139144 90766 139505
rect 90934 139144 92054 139505
rect 92222 139144 93342 139505
rect 93510 139144 94630 139505
rect 94798 139144 95918 139505
rect 96086 139144 97206 139505
rect 97374 139144 98494 139505
rect 98662 139144 99782 139505
rect 99950 139144 101070 139505
rect 101238 139144 102358 139505
rect 102526 139144 103646 139505
rect 103814 139144 104934 139505
rect 105102 139144 106222 139505
rect 106390 139144 107510 139505
rect 107678 139144 108798 139505
rect 108966 139144 110086 139505
rect 110254 139144 111374 139505
rect 111542 139144 112662 139505
rect 112830 139144 113950 139505
rect 114118 139144 115238 139505
rect 115406 139144 116526 139505
rect 116694 139144 117814 139505
rect 117982 139144 119102 139505
rect 119270 139144 120390 139505
rect 120558 139144 121678 139505
rect 121846 139144 122966 139505
rect 123134 139144 124254 139505
rect 124422 139144 125542 139505
rect 125710 139144 126830 139505
rect 126998 139144 128118 139505
rect 128286 139144 129406 139505
rect 129574 139144 130694 139505
rect 130862 139144 131982 139505
rect 132150 139144 133270 139505
rect 133438 139144 134558 139505
rect 134726 139144 135846 139505
rect 136014 139144 137134 139505
rect 137302 139144 138422 139505
rect 138590 139144 139710 139505
rect 20 856 139820 139144
rect 130 31 1250 856
rect 1418 31 2538 856
rect 2706 31 3826 856
rect 3994 31 5114 856
rect 5282 31 6402 856
rect 6570 31 7690 856
rect 7858 31 8978 856
rect 9146 31 10266 856
rect 10434 31 11554 856
rect 11722 31 12842 856
rect 13010 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16706 856
rect 16874 31 17994 856
rect 18162 31 19282 856
rect 19450 31 20570 856
rect 20738 31 21858 856
rect 22026 31 23146 856
rect 23314 31 24434 856
rect 24602 31 25722 856
rect 25890 31 27010 856
rect 27178 31 28298 856
rect 28466 31 29586 856
rect 29754 31 30874 856
rect 31042 31 32162 856
rect 32330 31 33450 856
rect 33618 31 34738 856
rect 34906 31 36026 856
rect 36194 31 37314 856
rect 37482 31 38602 856
rect 38770 31 39890 856
rect 40058 31 41178 856
rect 41346 31 42466 856
rect 42634 31 43754 856
rect 43922 31 45042 856
rect 45210 31 46330 856
rect 46498 31 47618 856
rect 47786 31 48906 856
rect 49074 31 50194 856
rect 50362 31 51482 856
rect 51650 31 52770 856
rect 52938 31 54058 856
rect 54226 31 55346 856
rect 55514 31 56634 856
rect 56802 31 57922 856
rect 58090 31 59210 856
rect 59378 31 60498 856
rect 60666 31 61786 856
rect 61954 31 63074 856
rect 63242 31 64362 856
rect 64530 31 65650 856
rect 65818 31 66938 856
rect 67106 31 68870 856
rect 69038 31 70158 856
rect 70326 31 71446 856
rect 71614 31 72734 856
rect 72902 31 74022 856
rect 74190 31 75310 856
rect 75478 31 76598 856
rect 76766 31 77886 856
rect 78054 31 79174 856
rect 79342 31 80462 856
rect 80630 31 81750 856
rect 81918 31 83038 856
rect 83206 31 84326 856
rect 84494 31 85614 856
rect 85782 31 86902 856
rect 87070 31 88190 856
rect 88358 31 89478 856
rect 89646 31 90766 856
rect 90934 31 92054 856
rect 92222 31 93342 856
rect 93510 31 94630 856
rect 94798 31 95918 856
rect 96086 31 97206 856
rect 97374 31 98494 856
rect 98662 31 99782 856
rect 99950 31 101070 856
rect 101238 31 102358 856
rect 102526 31 103646 856
rect 103814 31 104934 856
rect 105102 31 106222 856
rect 106390 31 107510 856
rect 107678 31 108798 856
rect 108966 31 110086 856
rect 110254 31 111374 856
rect 111542 31 112662 856
rect 112830 31 113950 856
rect 114118 31 115238 856
rect 115406 31 116526 856
rect 116694 31 117814 856
rect 117982 31 119102 856
rect 119270 31 120390 856
rect 120558 31 121678 856
rect 121846 31 122966 856
rect 123134 31 124254 856
rect 124422 31 125542 856
rect 125710 31 126830 856
rect 126998 31 128118 856
rect 128286 31 129406 856
rect 129574 31 130694 856
rect 130862 31 131982 856
rect 132150 31 133270 856
rect 133438 31 134558 856
rect 134726 31 136490 856
rect 136658 31 137778 856
rect 137946 31 139066 856
rect 139234 31 139820 856
<< metal3 >>
rect 0 139408 800 139528
rect 0 138048 800 138168
rect 139200 138048 140000 138168
rect 0 136688 800 136808
rect 139200 136688 140000 136808
rect 0 135328 800 135448
rect 139200 135328 140000 135448
rect 0 133968 800 134088
rect 139200 133968 140000 134088
rect 0 132608 800 132728
rect 139200 132608 140000 132728
rect 0 131248 800 131368
rect 139200 131248 140000 131368
rect 0 129888 800 130008
rect 139200 129888 140000 130008
rect 0 128528 800 128648
rect 139200 128528 140000 128648
rect 0 127168 800 127288
rect 139200 127168 140000 127288
rect 0 125808 800 125928
rect 139200 125808 140000 125928
rect 0 124448 800 124568
rect 139200 124448 140000 124568
rect 0 123088 800 123208
rect 139200 123088 140000 123208
rect 0 121728 800 121848
rect 139200 121728 140000 121848
rect 0 120368 800 120488
rect 139200 120368 140000 120488
rect 0 119008 800 119128
rect 139200 119008 140000 119128
rect 0 117648 800 117768
rect 139200 117648 140000 117768
rect 0 116288 800 116408
rect 139200 116288 140000 116408
rect 0 114928 800 115048
rect 139200 114928 140000 115048
rect 0 113568 800 113688
rect 139200 113568 140000 113688
rect 0 112208 800 112328
rect 139200 112208 140000 112328
rect 0 110848 800 110968
rect 139200 110848 140000 110968
rect 0 109488 800 109608
rect 139200 109488 140000 109608
rect 0 108128 800 108248
rect 139200 108128 140000 108248
rect 0 106768 800 106888
rect 139200 106768 140000 106888
rect 0 105408 800 105528
rect 139200 105408 140000 105528
rect 0 104048 800 104168
rect 139200 104048 140000 104168
rect 0 102688 800 102808
rect 139200 102688 140000 102808
rect 0 101328 800 101448
rect 139200 101328 140000 101448
rect 0 99968 800 100088
rect 139200 99968 140000 100088
rect 0 98608 800 98728
rect 139200 98608 140000 98728
rect 0 97248 800 97368
rect 139200 97248 140000 97368
rect 0 95888 800 96008
rect 139200 95888 140000 96008
rect 0 94528 800 94648
rect 139200 94528 140000 94648
rect 0 93168 800 93288
rect 139200 93168 140000 93288
rect 0 91808 800 91928
rect 139200 91808 140000 91928
rect 0 90448 800 90568
rect 139200 90448 140000 90568
rect 0 89088 800 89208
rect 139200 89088 140000 89208
rect 0 87728 800 87848
rect 139200 87728 140000 87848
rect 0 86368 800 86488
rect 139200 86368 140000 86488
rect 0 85008 800 85128
rect 139200 85008 140000 85128
rect 0 83648 800 83768
rect 139200 83648 140000 83768
rect 0 82288 800 82408
rect 139200 82288 140000 82408
rect 0 80928 800 81048
rect 139200 80928 140000 81048
rect 0 79568 800 79688
rect 139200 79568 140000 79688
rect 0 78208 800 78328
rect 139200 78208 140000 78328
rect 0 76848 800 76968
rect 139200 76848 140000 76968
rect 0 75488 800 75608
rect 139200 75488 140000 75608
rect 0 74128 800 74248
rect 139200 74128 140000 74248
rect 0 72768 800 72888
rect 139200 72768 140000 72888
rect 139200 71408 140000 71528
rect 0 70728 800 70848
rect 139200 70048 140000 70168
rect 0 69368 800 69488
rect 139200 68688 140000 68808
rect 0 68008 800 68128
rect 0 66648 800 66768
rect 139200 66648 140000 66768
rect 0 65288 800 65408
rect 139200 65288 140000 65408
rect 0 63928 800 64048
rect 139200 63928 140000 64048
rect 0 62568 800 62688
rect 139200 62568 140000 62688
rect 0 61208 800 61328
rect 139200 61208 140000 61328
rect 0 59848 800 59968
rect 139200 59848 140000 59968
rect 0 58488 800 58608
rect 139200 58488 140000 58608
rect 0 57128 800 57248
rect 139200 57128 140000 57248
rect 0 55768 800 55888
rect 139200 55768 140000 55888
rect 0 54408 800 54528
rect 139200 54408 140000 54528
rect 0 53048 800 53168
rect 139200 53048 140000 53168
rect 0 51688 800 51808
rect 139200 51688 140000 51808
rect 0 50328 800 50448
rect 139200 50328 140000 50448
rect 0 48968 800 49088
rect 139200 48968 140000 49088
rect 0 47608 800 47728
rect 139200 47608 140000 47728
rect 0 46248 800 46368
rect 139200 46248 140000 46368
rect 0 44888 800 45008
rect 139200 44888 140000 45008
rect 0 43528 800 43648
rect 139200 43528 140000 43648
rect 0 42168 800 42288
rect 139200 42168 140000 42288
rect 0 40808 800 40928
rect 139200 40808 140000 40928
rect 0 39448 800 39568
rect 139200 39448 140000 39568
rect 0 38088 800 38208
rect 139200 38088 140000 38208
rect 0 36728 800 36848
rect 139200 36728 140000 36848
rect 0 35368 800 35488
rect 139200 35368 140000 35488
rect 0 34008 800 34128
rect 139200 34008 140000 34128
rect 0 32648 800 32768
rect 139200 32648 140000 32768
rect 0 31288 800 31408
rect 139200 31288 140000 31408
rect 0 29928 800 30048
rect 139200 29928 140000 30048
rect 0 28568 800 28688
rect 139200 28568 140000 28688
rect 0 27208 800 27328
rect 139200 27208 140000 27328
rect 0 25848 800 25968
rect 139200 25848 140000 25968
rect 0 24488 800 24608
rect 139200 24488 140000 24608
rect 0 23128 800 23248
rect 139200 23128 140000 23248
rect 0 21768 800 21888
rect 139200 21768 140000 21888
rect 0 20408 800 20528
rect 139200 20408 140000 20528
rect 0 19048 800 19168
rect 139200 19048 140000 19168
rect 0 17688 800 17808
rect 139200 17688 140000 17808
rect 0 16328 800 16448
rect 139200 16328 140000 16448
rect 0 14968 800 15088
rect 139200 14968 140000 15088
rect 0 13608 800 13728
rect 139200 13608 140000 13728
rect 0 12248 800 12368
rect 139200 12248 140000 12368
rect 0 10888 800 11008
rect 139200 10888 140000 11008
rect 0 9528 800 9648
rect 139200 9528 140000 9648
rect 0 8168 800 8288
rect 139200 8168 140000 8288
rect 0 6808 800 6928
rect 139200 6808 140000 6928
rect 0 5448 800 5568
rect 139200 5448 140000 5568
rect 0 4088 800 4208
rect 139200 4088 140000 4208
rect 0 2728 800 2848
rect 139200 2728 140000 2848
rect 0 1368 800 1488
rect 139200 1368 140000 1488
rect 139200 8 140000 128
<< obsm3 >>
rect 880 139328 139200 139501
rect 800 138248 139200 139328
rect 880 137968 139120 138248
rect 800 136888 139200 137968
rect 880 136608 139120 136888
rect 800 135528 139200 136608
rect 880 135248 139120 135528
rect 800 134168 139200 135248
rect 880 133888 139120 134168
rect 800 132808 139200 133888
rect 880 132528 139120 132808
rect 800 131448 139200 132528
rect 880 131168 139120 131448
rect 800 130088 139200 131168
rect 880 129808 139120 130088
rect 800 128728 139200 129808
rect 880 128448 139120 128728
rect 800 127368 139200 128448
rect 880 127088 139120 127368
rect 800 126008 139200 127088
rect 880 125728 139120 126008
rect 800 124648 139200 125728
rect 880 124368 139120 124648
rect 800 123288 139200 124368
rect 880 123008 139120 123288
rect 800 121928 139200 123008
rect 880 121648 139120 121928
rect 800 120568 139200 121648
rect 880 120288 139120 120568
rect 800 119208 139200 120288
rect 880 118928 139120 119208
rect 800 117848 139200 118928
rect 880 117568 139120 117848
rect 800 116488 139200 117568
rect 880 116208 139120 116488
rect 800 115128 139200 116208
rect 880 114848 139120 115128
rect 800 113768 139200 114848
rect 880 113488 139120 113768
rect 800 112408 139200 113488
rect 880 112128 139120 112408
rect 800 111048 139200 112128
rect 880 110768 139120 111048
rect 800 109688 139200 110768
rect 880 109408 139120 109688
rect 800 108328 139200 109408
rect 880 108048 139120 108328
rect 800 106968 139200 108048
rect 880 106688 139120 106968
rect 800 105608 139200 106688
rect 880 105328 139120 105608
rect 800 104248 139200 105328
rect 880 103968 139120 104248
rect 800 102888 139200 103968
rect 880 102608 139120 102888
rect 800 101528 139200 102608
rect 880 101248 139120 101528
rect 800 100168 139200 101248
rect 880 99888 139120 100168
rect 800 98808 139200 99888
rect 880 98528 139120 98808
rect 800 97448 139200 98528
rect 880 97168 139120 97448
rect 800 96088 139200 97168
rect 880 95808 139120 96088
rect 800 94728 139200 95808
rect 880 94448 139120 94728
rect 800 93368 139200 94448
rect 880 93088 139120 93368
rect 800 92008 139200 93088
rect 880 91728 139120 92008
rect 800 90648 139200 91728
rect 880 90368 139120 90648
rect 800 89288 139200 90368
rect 880 89008 139120 89288
rect 800 87928 139200 89008
rect 880 87648 139120 87928
rect 800 86568 139200 87648
rect 880 86288 139120 86568
rect 800 85208 139200 86288
rect 880 84928 139120 85208
rect 800 83848 139200 84928
rect 880 83568 139120 83848
rect 800 82488 139200 83568
rect 880 82208 139120 82488
rect 800 81128 139200 82208
rect 880 80848 139120 81128
rect 800 79768 139200 80848
rect 880 79488 139120 79768
rect 800 78408 139200 79488
rect 880 78128 139120 78408
rect 800 77048 139200 78128
rect 880 76768 139120 77048
rect 800 75688 139200 76768
rect 880 75408 139120 75688
rect 800 74328 139200 75408
rect 880 74048 139120 74328
rect 800 72968 139200 74048
rect 880 72688 139120 72968
rect 800 71608 139200 72688
rect 800 71328 139120 71608
rect 800 70928 139200 71328
rect 880 70648 139200 70928
rect 800 70248 139200 70648
rect 800 69968 139120 70248
rect 800 69568 139200 69968
rect 880 69288 139200 69568
rect 800 68888 139200 69288
rect 800 68608 139120 68888
rect 800 68208 139200 68608
rect 880 67928 139200 68208
rect 800 66848 139200 67928
rect 880 66568 139120 66848
rect 800 65488 139200 66568
rect 880 65208 139120 65488
rect 800 64128 139200 65208
rect 880 63848 139120 64128
rect 800 62768 139200 63848
rect 880 62488 139120 62768
rect 800 61408 139200 62488
rect 880 61128 139120 61408
rect 800 60048 139200 61128
rect 880 59768 139120 60048
rect 800 58688 139200 59768
rect 880 58408 139120 58688
rect 800 57328 139200 58408
rect 880 57048 139120 57328
rect 800 55968 139200 57048
rect 880 55688 139120 55968
rect 800 54608 139200 55688
rect 880 54328 139120 54608
rect 800 53248 139200 54328
rect 880 52968 139120 53248
rect 800 51888 139200 52968
rect 880 51608 139120 51888
rect 800 50528 139200 51608
rect 880 50248 139120 50528
rect 800 49168 139200 50248
rect 880 48888 139120 49168
rect 800 47808 139200 48888
rect 880 47528 139120 47808
rect 800 46448 139200 47528
rect 880 46168 139120 46448
rect 800 45088 139200 46168
rect 880 44808 139120 45088
rect 800 43728 139200 44808
rect 880 43448 139120 43728
rect 800 42368 139200 43448
rect 880 42088 139120 42368
rect 800 41008 139200 42088
rect 880 40728 139120 41008
rect 800 39648 139200 40728
rect 880 39368 139120 39648
rect 800 38288 139200 39368
rect 880 38008 139120 38288
rect 800 36928 139200 38008
rect 880 36648 139120 36928
rect 800 35568 139200 36648
rect 880 35288 139120 35568
rect 800 34208 139200 35288
rect 880 33928 139120 34208
rect 800 32848 139200 33928
rect 880 32568 139120 32848
rect 800 31488 139200 32568
rect 880 31208 139120 31488
rect 800 30128 139200 31208
rect 880 29848 139120 30128
rect 800 28768 139200 29848
rect 880 28488 139120 28768
rect 800 27408 139200 28488
rect 880 27128 139120 27408
rect 800 26048 139200 27128
rect 880 25768 139120 26048
rect 800 24688 139200 25768
rect 880 24408 139120 24688
rect 800 23328 139200 24408
rect 880 23048 139120 23328
rect 800 21968 139200 23048
rect 880 21688 139120 21968
rect 800 20608 139200 21688
rect 880 20328 139120 20608
rect 800 19248 139200 20328
rect 880 18968 139120 19248
rect 800 17888 139200 18968
rect 880 17608 139120 17888
rect 800 16528 139200 17608
rect 880 16248 139120 16528
rect 800 15168 139200 16248
rect 880 14888 139120 15168
rect 800 13808 139200 14888
rect 880 13528 139120 13808
rect 800 12448 139200 13528
rect 880 12168 139120 12448
rect 800 11088 139200 12168
rect 880 10808 139120 11088
rect 800 9728 139200 10808
rect 880 9448 139120 9728
rect 800 8368 139200 9448
rect 880 8088 139120 8368
rect 800 7008 139200 8088
rect 880 6728 139120 7008
rect 800 5648 139200 6728
rect 880 5368 139120 5648
rect 800 4288 139200 5368
rect 880 4008 139120 4288
rect 800 2928 139200 4008
rect 880 2648 139120 2928
rect 800 1568 139200 2648
rect 880 1288 139120 1568
rect 800 208 139200 1288
rect 800 35 139120 208
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< obsm4 >>
rect 54155 2619 65568 136781
rect 66048 2619 80928 136781
rect 81408 2619 87341 136781
<< labels >>
rlabel metal2 s 57978 0 58034 800 6 clock
port 1 nsew signal input
rlabel metal2 s 14186 139200 14242 140000 6 io_dbus_addr[0]
port 2 nsew signal input
rlabel metal2 s 57978 139200 58034 140000 6 io_dbus_addr[10]
port 3 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 io_dbus_addr[11]
port 4 nsew signal input
rlabel metal3 s 139200 19048 140000 19168 6 io_dbus_addr[12]
port 5 nsew signal input
rlabel metal2 s 11610 139200 11666 140000 6 io_dbus_addr[13]
port 6 nsew signal input
rlabel metal3 s 139200 53048 140000 53168 6 io_dbus_addr[14]
port 7 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 io_dbus_addr[15]
port 8 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 io_dbus_addr[16]
port 9 nsew signal input
rlabel metal3 s 139200 82288 140000 82408 6 io_dbus_addr[17]
port 10 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 io_dbus_addr[18]
port 11 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_dbus_addr[19]
port 12 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 io_dbus_addr[1]
port 13 nsew signal input
rlabel metal3 s 139200 32648 140000 32768 6 io_dbus_addr[20]
port 14 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 io_dbus_addr[21]
port 15 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 io_dbus_addr[22]
port 16 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_dbus_addr[23]
port 17 nsew signal input
rlabel metal3 s 139200 90448 140000 90568 6 io_dbus_addr[24]
port 18 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 io_dbus_addr[25]
port 19 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 io_dbus_addr[26]
port 20 nsew signal input
rlabel metal3 s 139200 132608 140000 132728 6 io_dbus_addr[27]
port 21 nsew signal input
rlabel metal3 s 139200 25848 140000 25968 6 io_dbus_addr[28]
port 22 nsew signal input
rlabel metal3 s 139200 110848 140000 110968 6 io_dbus_addr[29]
port 23 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 io_dbus_addr[2]
port 24 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 io_dbus_addr[30]
port 25 nsew signal input
rlabel metal3 s 139200 48968 140000 49088 6 io_dbus_addr[31]
port 26 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 io_dbus_addr[3]
port 27 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 io_dbus_addr[4]
port 28 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 io_dbus_addr[5]
port 29 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 io_dbus_addr[6]
port 30 nsew signal input
rlabel metal2 s 12898 139200 12954 140000 6 io_dbus_addr[7]
port 31 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 io_dbus_addr[8]
port 32 nsew signal input
rlabel metal2 s 138478 139200 138534 140000 6 io_dbus_addr[9]
port 33 nsew signal input
rlabel metal2 s 112718 139200 112774 140000 6 io_dbus_ld_type[0]
port 34 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 io_dbus_ld_type[1]
port 35 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 io_dbus_ld_type[2]
port 36 nsew signal input
rlabel metal3 s 139200 23128 140000 23248 6 io_dbus_rd_en
port 37 nsew signal input
rlabel metal3 s 139200 27208 140000 27328 6 io_dbus_rdata[0]
port 38 nsew signal output
rlabel metal2 s 70858 139200 70914 140000 6 io_dbus_rdata[10]
port 39 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_dbus_rdata[11]
port 40 nsew signal output
rlabel metal3 s 139200 34008 140000 34128 6 io_dbus_rdata[12]
port 41 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 io_dbus_rdata[13]
port 42 nsew signal output
rlabel metal2 s 85670 139200 85726 140000 6 io_dbus_rdata[14]
port 43 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 io_dbus_rdata[15]
port 44 nsew signal output
rlabel metal2 s 125598 139200 125654 140000 6 io_dbus_rdata[16]
port 45 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 io_dbus_rdata[17]
port 46 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 io_dbus_rdata[18]
port 47 nsew signal output
rlabel metal2 s 72790 139200 72846 140000 6 io_dbus_rdata[19]
port 48 nsew signal output
rlabel metal2 s 124310 139200 124366 140000 6 io_dbus_rdata[1]
port 49 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 io_dbus_rdata[20]
port 50 nsew signal output
rlabel metal2 s 72790 0 72846 800 6 io_dbus_rdata[21]
port 51 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 io_dbus_rdata[22]
port 52 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 io_dbus_rdata[23]
port 53 nsew signal output
rlabel metal3 s 139200 87728 140000 87848 6 io_dbus_rdata[24]
port 54 nsew signal output
rlabel metal2 s 139766 139200 139822 140000 6 io_dbus_rdata[25]
port 55 nsew signal output
rlabel metal3 s 139200 136688 140000 136808 6 io_dbus_rdata[26]
port 56 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 io_dbus_rdata[27]
port 57 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 io_dbus_rdata[28]
port 58 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 io_dbus_rdata[29]
port 59 nsew signal output
rlabel metal3 s 139200 112208 140000 112328 6 io_dbus_rdata[2]
port 60 nsew signal output
rlabel metal3 s 139200 125808 140000 125928 6 io_dbus_rdata[30]
port 61 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 io_dbus_rdata[31]
port 62 nsew signal output
rlabel metal3 s 139200 108128 140000 108248 6 io_dbus_rdata[3]
port 63 nsew signal output
rlabel metal2 s 81806 139200 81862 140000 6 io_dbus_rdata[4]
port 64 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 io_dbus_rdata[5]
port 65 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 io_dbus_rdata[6]
port 66 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 io_dbus_rdata[7]
port 67 nsew signal output
rlabel metal2 s 662 139200 718 140000 6 io_dbus_rdata[8]
port 68 nsew signal output
rlabel metal2 s 117870 139200 117926 140000 6 io_dbus_rdata[9]
port 69 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 io_dbus_st_type[0]
port 70 nsew signal input
rlabel metal3 s 139200 20408 140000 20528 6 io_dbus_st_type[1]
port 71 nsew signal input
rlabel metal3 s 139200 99968 140000 100088 6 io_dbus_valid
port 72 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 io_dbus_wdata[0]
port 73 nsew signal input
rlabel metal2 s 79230 139200 79286 140000 6 io_dbus_wdata[10]
port 74 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 io_dbus_wdata[11]
port 75 nsew signal input
rlabel metal2 s 32218 139200 32274 140000 6 io_dbus_wdata[12]
port 76 nsew signal input
rlabel metal2 s 24490 139200 24546 140000 6 io_dbus_wdata[13]
port 77 nsew signal input
rlabel metal3 s 139200 75488 140000 75608 6 io_dbus_wdata[14]
port 78 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 io_dbus_wdata[15]
port 79 nsew signal input
rlabel metal2 s 75366 139200 75422 140000 6 io_dbus_wdata[16]
port 80 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 io_dbus_wdata[17]
port 81 nsew signal input
rlabel metal3 s 139200 55768 140000 55888 6 io_dbus_wdata[18]
port 82 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 io_dbus_wdata[19]
port 83 nsew signal input
rlabel metal2 s 56690 139200 56746 140000 6 io_dbus_wdata[1]
port 84 nsew signal input
rlabel metal2 s 114006 139200 114062 140000 6 io_dbus_wdata[20]
port 85 nsew signal input
rlabel metal2 s 80518 139200 80574 140000 6 io_dbus_wdata[21]
port 86 nsew signal input
rlabel metal2 s 77942 139200 77998 140000 6 io_dbus_wdata[22]
port 87 nsew signal input
rlabel metal3 s 139200 12248 140000 12368 6 io_dbus_wdata[23]
port 88 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_dbus_wdata[24]
port 89 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 io_dbus_wdata[25]
port 90 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 io_dbus_wdata[26]
port 91 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 io_dbus_wdata[27]
port 92 nsew signal input
rlabel metal2 s 6458 139200 6514 140000 6 io_dbus_wdata[28]
port 93 nsew signal input
rlabel metal3 s 139200 5448 140000 5568 6 io_dbus_wdata[29]
port 94 nsew signal input
rlabel metal2 s 110142 139200 110198 140000 6 io_dbus_wdata[2]
port 95 nsew signal input
rlabel metal3 s 0 123088 800 123208 6 io_dbus_wdata[30]
port 96 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 io_dbus_wdata[31]
port 97 nsew signal input
rlabel metal2 s 65706 139200 65762 140000 6 io_dbus_wdata[3]
port 98 nsew signal input
rlabel metal3 s 139200 129888 140000 130008 6 io_dbus_wdata[4]
port 99 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 io_dbus_wdata[5]
port 100 nsew signal input
rlabel metal2 s 89534 139200 89590 140000 6 io_dbus_wdata[6]
port 101 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 io_dbus_wdata[7]
port 102 nsew signal input
rlabel metal2 s 97262 139200 97318 140000 6 io_dbus_wdata[8]
port 103 nsew signal input
rlabel metal2 s 76654 139200 76710 140000 6 io_dbus_wdata[9]
port 104 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 io_dbus_wr_en
port 105 nsew signal input
rlabel metal2 s 27066 139200 27122 140000 6 io_dmem_io_addr[0]
port 106 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 io_dmem_io_addr[1]
port 107 nsew signal output
rlabel metal2 s 108854 139200 108910 140000 6 io_dmem_io_addr[2]
port 108 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 io_dmem_io_addr[3]
port 109 nsew signal output
rlabel metal3 s 139200 74128 140000 74248 6 io_dmem_io_addr[4]
port 110 nsew signal output
rlabel metal2 s 99838 139200 99894 140000 6 io_dmem_io_addr[5]
port 111 nsew signal output
rlabel metal3 s 139200 85008 140000 85128 6 io_dmem_io_addr[6]
port 112 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 io_dmem_io_addr[7]
port 113 nsew signal output
rlabel metal2 s 15474 139200 15530 140000 6 io_dmem_io_cs
port 114 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 io_dmem_io_rdata[0]
port 115 nsew signal input
rlabel metal2 s 84382 139200 84438 140000 6 io_dmem_io_rdata[10]
port 116 nsew signal input
rlabel metal2 s 38658 139200 38714 140000 6 io_dmem_io_rdata[11]
port 117 nsew signal input
rlabel metal2 s 102414 139200 102470 140000 6 io_dmem_io_rdata[12]
port 118 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 io_dmem_io_rdata[13]
port 119 nsew signal input
rlabel metal3 s 139200 116288 140000 116408 6 io_dmem_io_rdata[14]
port 120 nsew signal input
rlabel metal3 s 139200 62568 140000 62688 6 io_dmem_io_rdata[15]
port 121 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 io_dmem_io_rdata[16]
port 122 nsew signal input
rlabel metal3 s 139200 28568 140000 28688 6 io_dmem_io_rdata[17]
port 123 nsew signal input
rlabel metal2 s 128174 139200 128230 140000 6 io_dmem_io_rdata[18]
port 124 nsew signal input
rlabel metal3 s 139200 61208 140000 61328 6 io_dmem_io_rdata[19]
port 125 nsew signal input
rlabel metal2 s 7746 139200 7802 140000 6 io_dmem_io_rdata[1]
port 126 nsew signal input
rlabel metal2 s 5170 139200 5226 140000 6 io_dmem_io_rdata[20]
port 127 nsew signal input
rlabel metal2 s 86958 139200 87014 140000 6 io_dmem_io_rdata[21]
port 128 nsew signal input
rlabel metal3 s 139200 44888 140000 45008 6 io_dmem_io_rdata[22]
port 129 nsew signal input
rlabel metal2 s 33506 139200 33562 140000 6 io_dmem_io_rdata[23]
port 130 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 io_dmem_io_rdata[24]
port 131 nsew signal input
rlabel metal3 s 139200 59848 140000 59968 6 io_dmem_io_rdata[25]
port 132 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 io_dmem_io_rdata[26]
port 133 nsew signal input
rlabel metal2 s 9034 139200 9090 140000 6 io_dmem_io_rdata[27]
port 134 nsew signal input
rlabel metal2 s 120446 139200 120502 140000 6 io_dmem_io_rdata[28]
port 135 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 io_dmem_io_rdata[29]
port 136 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 io_dmem_io_rdata[2]
port 137 nsew signal input
rlabel metal3 s 139200 123088 140000 123208 6 io_dmem_io_rdata[30]
port 138 nsew signal input
rlabel metal3 s 139200 105408 140000 105528 6 io_dmem_io_rdata[31]
port 139 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 io_dmem_io_rdata[3]
port 140 nsew signal input
rlabel metal2 s 37370 139200 37426 140000 6 io_dmem_io_rdata[4]
port 141 nsew signal input
rlabel metal2 s 88246 139200 88302 140000 6 io_dmem_io_rdata[5]
port 142 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 io_dmem_io_rdata[6]
port 143 nsew signal input
rlabel metal3 s 139200 138048 140000 138168 6 io_dmem_io_rdata[7]
port 144 nsew signal input
rlabel metal3 s 139200 79568 140000 79688 6 io_dmem_io_rdata[8]
port 145 nsew signal input
rlabel metal3 s 0 127168 800 127288 6 io_dmem_io_rdata[9]
port 146 nsew signal input
rlabel metal3 s 139200 119008 140000 119128 6 io_dmem_io_st_type[0]
port 147 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 io_dmem_io_st_type[1]
port 148 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 io_dmem_io_st_type[2]
port 149 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 io_dmem_io_st_type[3]
port 150 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 io_dmem_io_wdata[0]
port 151 nsew signal output
rlabel metal3 s 139200 47608 140000 47728 6 io_dmem_io_wdata[10]
port 152 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 io_dmem_io_wdata[11]
port 153 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 io_dmem_io_wdata[12]
port 154 nsew signal output
rlabel metal3 s 139200 131248 140000 131368 6 io_dmem_io_wdata[13]
port 155 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 io_dmem_io_wdata[14]
port 156 nsew signal output
rlabel metal2 s 135902 139200 135958 140000 6 io_dmem_io_wdata[15]
port 157 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 io_dmem_io_wdata[16]
port 158 nsew signal output
rlabel metal3 s 139200 104048 140000 104168 6 io_dmem_io_wdata[17]
port 159 nsew signal output
rlabel metal2 s 85670 0 85726 800 6 io_dmem_io_wdata[18]
port 160 nsew signal output
rlabel metal3 s 139200 135328 140000 135448 6 io_dmem_io_wdata[19]
port 161 nsew signal output
rlabel metal2 s 20626 139200 20682 140000 6 io_dmem_io_wdata[1]
port 162 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_dmem_io_wdata[20]
port 163 nsew signal output
rlabel metal2 s 55402 139200 55458 140000 6 io_dmem_io_wdata[21]
port 164 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 io_dmem_io_wdata[22]
port 165 nsew signal output
rlabel metal2 s 1950 139200 2006 140000 6 io_dmem_io_wdata[23]
port 166 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 io_dmem_io_wdata[24]
port 167 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 io_dmem_io_wdata[25]
port 168 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 io_dmem_io_wdata[26]
port 169 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 io_dmem_io_wdata[27]
port 170 nsew signal output
rlabel metal2 s 47674 139200 47730 140000 6 io_dmem_io_wdata[28]
port 171 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 io_dmem_io_wdata[29]
port 172 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 io_dmem_io_wdata[2]
port 173 nsew signal output
rlabel metal2 s 68282 139200 68338 140000 6 io_dmem_io_wdata[30]
port 174 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 io_dmem_io_wdata[31]
port 175 nsew signal output
rlabel metal2 s 52826 139200 52882 140000 6 io_dmem_io_wdata[3]
port 176 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 io_dmem_io_wdata[4]
port 177 nsew signal output
rlabel metal3 s 139200 70048 140000 70168 6 io_dmem_io_wdata[5]
port 178 nsew signal output
rlabel metal2 s 45098 139200 45154 140000 6 io_dmem_io_wdata[6]
port 179 nsew signal output
rlabel metal3 s 139200 50328 140000 50448 6 io_dmem_io_wdata[7]
port 180 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 io_dmem_io_wdata[8]
port 181 nsew signal output
rlabel metal2 s 21914 139200 21970 140000 6 io_dmem_io_wdata[9]
port 182 nsew signal output
rlabel metal3 s 0 138048 800 138168 6 io_dmem_io_wr_en
port 183 nsew signal output
rlabel metal3 s 139200 76848 140000 76968 6 io_ibus_addr[0]
port 184 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 io_ibus_addr[10]
port 185 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_ibus_addr[11]
port 186 nsew signal input
rlabel metal2 s 39946 139200 40002 140000 6 io_ibus_addr[12]
port 187 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 io_ibus_addr[13]
port 188 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 io_ibus_addr[14]
port 189 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 io_ibus_addr[15]
port 190 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 io_ibus_addr[16]
port 191 nsew signal input
rlabel metal3 s 139200 117648 140000 117768 6 io_ibus_addr[17]
port 192 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 io_ibus_addr[18]
port 193 nsew signal input
rlabel metal2 s 69570 139200 69626 140000 6 io_ibus_addr[19]
port 194 nsew signal input
rlabel metal2 s 134614 139200 134670 140000 6 io_ibus_addr[1]
port 195 nsew signal input
rlabel metal3 s 139200 101328 140000 101448 6 io_ibus_addr[20]
port 196 nsew signal input
rlabel metal2 s 30930 139200 30986 140000 6 io_ibus_addr[21]
port 197 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 io_ibus_addr[22]
port 198 nsew signal input
rlabel metal2 s 130750 139200 130806 140000 6 io_ibus_addr[23]
port 199 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_ibus_addr[24]
port 200 nsew signal input
rlabel metal3 s 139200 16328 140000 16448 6 io_ibus_addr[25]
port 201 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_ibus_addr[26]
port 202 nsew signal input
rlabel metal3 s 139200 113568 140000 113688 6 io_ibus_addr[27]
port 203 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 io_ibus_addr[28]
port 204 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_ibus_addr[29]
port 205 nsew signal input
rlabel metal3 s 139200 63928 140000 64048 6 io_ibus_addr[2]
port 206 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 io_ibus_addr[30]
port 207 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 io_ibus_addr[31]
port 208 nsew signal input
rlabel metal3 s 139200 24488 140000 24608 6 io_ibus_addr[3]
port 209 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 io_ibus_addr[4]
port 210 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 io_ibus_addr[5]
port 211 nsew signal input
rlabel metal2 s 61842 139200 61898 140000 6 io_ibus_addr[6]
port 212 nsew signal input
rlabel metal3 s 139200 54408 140000 54528 6 io_ibus_addr[7]
port 213 nsew signal input
rlabel metal3 s 139200 8 140000 128 6 io_ibus_addr[8]
port 214 nsew signal input
rlabel metal3 s 139200 17688 140000 17808 6 io_ibus_addr[9]
port 215 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 io_ibus_inst[0]
port 216 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 io_ibus_inst[10]
port 217 nsew signal output
rlabel metal3 s 139200 40808 140000 40928 6 io_ibus_inst[11]
port 218 nsew signal output
rlabel metal2 s 63130 139200 63186 140000 6 io_ibus_inst[12]
port 219 nsew signal output
rlabel metal2 s 7746 0 7802 800 6 io_ibus_inst[13]
port 220 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 io_ibus_inst[14]
port 221 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 io_ibus_inst[15]
port 222 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 io_ibus_inst[16]
port 223 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 io_ibus_inst[17]
port 224 nsew signal output
rlabel metal2 s 23202 139200 23258 140000 6 io_ibus_inst[18]
port 225 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 io_ibus_inst[19]
port 226 nsew signal output
rlabel metal2 s 66994 139200 67050 140000 6 io_ibus_inst[1]
port 227 nsew signal output
rlabel metal3 s 139200 14968 140000 15088 6 io_ibus_inst[20]
port 228 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 io_ibus_inst[21]
port 229 nsew signal output
rlabel metal3 s 139200 6808 140000 6928 6 io_ibus_inst[22]
port 230 nsew signal output
rlabel metal2 s 16762 139200 16818 140000 6 io_ibus_inst[23]
port 231 nsew signal output
rlabel metal3 s 139200 95888 140000 96008 6 io_ibus_inst[24]
port 232 nsew signal output
rlabel metal2 s 59266 139200 59322 140000 6 io_ibus_inst[25]
port 233 nsew signal output
rlabel metal3 s 139200 31288 140000 31408 6 io_ibus_inst[26]
port 234 nsew signal output
rlabel metal2 s 104990 139200 105046 140000 6 io_ibus_inst[27]
port 235 nsew signal output
rlabel metal3 s 139200 97248 140000 97368 6 io_ibus_inst[28]
port 236 nsew signal output
rlabel metal3 s 139200 127168 140000 127288 6 io_ibus_inst[29]
port 237 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 io_ibus_inst[2]
port 238 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 io_ibus_inst[30]
port 239 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 io_ibus_inst[31]
port 240 nsew signal output
rlabel metal2 s 119158 0 119214 800 6 io_ibus_inst[3]
port 241 nsew signal output
rlabel metal3 s 139200 8168 140000 8288 6 io_ibus_inst[4]
port 242 nsew signal output
rlabel metal3 s 139200 38088 140000 38208 6 io_ibus_inst[5]
port 243 nsew signal output
rlabel metal2 s 50250 139200 50306 140000 6 io_ibus_inst[6]
port 244 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 io_ibus_inst[7]
port 245 nsew signal output
rlabel metal3 s 139200 65288 140000 65408 6 io_ibus_inst[8]
port 246 nsew signal output
rlabel metal3 s 139200 51688 140000 51808 6 io_ibus_inst[9]
port 247 nsew signal output
rlabel metal3 s 139200 98608 140000 98728 6 io_ibus_valid
port 248 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 io_imem_io_addr[0]
port 249 nsew signal output
rlabel metal2 s 54114 139200 54170 140000 6 io_imem_io_addr[1]
port 250 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 io_imem_io_addr[2]
port 251 nsew signal output
rlabel metal2 s 101126 0 101182 800 6 io_imem_io_addr[3]
port 252 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 io_imem_io_addr[4]
port 253 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 io_imem_io_addr[5]
port 254 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 io_imem_io_addr[6]
port 255 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 io_imem_io_addr[7]
port 256 nsew signal output
rlabel metal3 s 139200 9528 140000 9648 6 io_imem_io_addr[8]
port 257 nsew signal output
rlabel metal2 s 3238 139200 3294 140000 6 io_imem_io_cs
port 258 nsew signal output
rlabel metal2 s 126886 139200 126942 140000 6 io_imem_io_rdata[0]
port 259 nsew signal input
rlabel metal2 s 121734 139200 121790 140000 6 io_imem_io_rdata[10]
port 260 nsew signal input
rlabel metal2 s 103702 139200 103758 140000 6 io_imem_io_rdata[11]
port 261 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 io_imem_io_rdata[12]
port 262 nsew signal input
rlabel metal3 s 139200 86368 140000 86488 6 io_imem_io_rdata[13]
port 263 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 io_imem_io_rdata[14]
port 264 nsew signal input
rlabel metal2 s 29642 139200 29698 140000 6 io_imem_io_rdata[15]
port 265 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 io_imem_io_rdata[16]
port 266 nsew signal input
rlabel metal3 s 139200 72768 140000 72888 6 io_imem_io_rdata[17]
port 267 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 io_imem_io_rdata[18]
port 268 nsew signal input
rlabel metal2 s 137190 139200 137246 140000 6 io_imem_io_rdata[19]
port 269 nsew signal input
rlabel metal3 s 139200 120368 140000 120488 6 io_imem_io_rdata[1]
port 270 nsew signal input
rlabel metal2 s 60554 139200 60610 140000 6 io_imem_io_rdata[20]
port 271 nsew signal input
rlabel metal3 s 139200 114928 140000 115048 6 io_imem_io_rdata[21]
port 272 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 io_imem_io_rdata[22]
port 273 nsew signal input
rlabel metal2 s 25778 139200 25834 140000 6 io_imem_io_rdata[23]
port 274 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 io_imem_io_rdata[24]
port 275 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 io_imem_io_rdata[25]
port 276 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 io_imem_io_rdata[26]
port 277 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 io_imem_io_rdata[27]
port 278 nsew signal input
rlabel metal3 s 139200 2728 140000 2848 6 io_imem_io_rdata[28]
port 279 nsew signal input
rlabel metal2 s 132038 139200 132094 140000 6 io_imem_io_rdata[29]
port 280 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 io_imem_io_rdata[2]
port 281 nsew signal input
rlabel metal2 s 51538 139200 51594 140000 6 io_imem_io_rdata[30]
port 282 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 io_imem_io_rdata[31]
port 283 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 io_imem_io_rdata[3]
port 284 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 io_imem_io_rdata[4]
port 285 nsew signal input
rlabel metal2 s 115294 139200 115350 140000 6 io_imem_io_rdata[5]
port 286 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 io_imem_io_rdata[6]
port 287 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 io_imem_io_rdata[7]
port 288 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 io_imem_io_rdata[8]
port 289 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_imem_io_rdata[9]
port 290 nsew signal input
rlabel metal3 s 139200 93168 140000 93288 6 io_imem_io_wdata[0]
port 291 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 io_imem_io_wdata[10]
port 292 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 io_imem_io_wdata[11]
port 293 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 io_imem_io_wdata[12]
port 294 nsew signal output
rlabel metal3 s 139200 89088 140000 89208 6 io_imem_io_wdata[13]
port 295 nsew signal output
rlabel metal2 s 94686 139200 94742 140000 6 io_imem_io_wdata[14]
port 296 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 io_imem_io_wdata[15]
port 297 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 io_imem_io_wdata[16]
port 298 nsew signal output
rlabel metal2 s 123022 139200 123078 140000 6 io_imem_io_wdata[17]
port 299 nsew signal output
rlabel metal3 s 139200 10888 140000 11008 6 io_imem_io_wdata[18]
port 300 nsew signal output
rlabel metal2 s 83094 139200 83150 140000 6 io_imem_io_wdata[19]
port 301 nsew signal output
rlabel metal2 s 126886 0 126942 800 6 io_imem_io_wdata[1]
port 302 nsew signal output
rlabel metal2 s 34794 139200 34850 140000 6 io_imem_io_wdata[20]
port 303 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 io_imem_io_wdata[21]
port 304 nsew signal output
rlabel metal3 s 139200 68688 140000 68808 6 io_imem_io_wdata[22]
port 305 nsew signal output
rlabel metal3 s 0 135328 800 135448 6 io_imem_io_wdata[23]
port 306 nsew signal output
rlabel metal3 s 139200 91808 140000 91928 6 io_imem_io_wdata[24]
port 307 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 io_imem_io_wdata[25]
port 308 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 io_imem_io_wdata[26]
port 309 nsew signal output
rlabel metal2 s 42522 139200 42578 140000 6 io_imem_io_wdata[27]
port 310 nsew signal output
rlabel metal2 s 119158 139200 119214 140000 6 io_imem_io_wdata[28]
port 311 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 io_imem_io_wdata[29]
port 312 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 io_imem_io_wdata[2]
port 313 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 io_imem_io_wdata[30]
port 314 nsew signal output
rlabel metal3 s 139200 21768 140000 21888 6 io_imem_io_wdata[31]
port 315 nsew signal output
rlabel metal2 s 28354 139200 28410 140000 6 io_imem_io_wdata[3]
port 316 nsew signal output
rlabel metal3 s 139200 46248 140000 46368 6 io_imem_io_wdata[4]
port 317 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_imem_io_wdata[5]
port 318 nsew signal output
rlabel metal2 s 64418 139200 64474 140000 6 io_imem_io_wdata[6]
port 319 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 io_imem_io_wdata[7]
port 320 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 io_imem_io_wdata[8]
port 321 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 io_imem_io_wdata[9]
port 322 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 io_imem_io_wr_en
port 323 nsew signal output
rlabel metal3 s 139200 94528 140000 94648 6 io_motor_ack_i
port 324 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 io_motor_addr_sel
port 325 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 io_motor_data_i[0]
port 326 nsew signal input
rlabel metal3 s 139200 42168 140000 42288 6 io_motor_data_i[10]
port 327 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 io_motor_data_i[11]
port 328 nsew signal input
rlabel metal2 s 90822 139200 90878 140000 6 io_motor_data_i[12]
port 329 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 io_motor_data_i[13]
port 330 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 io_motor_data_i[14]
port 331 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 io_motor_data_i[15]
port 332 nsew signal input
rlabel metal3 s 139200 29928 140000 30048 6 io_motor_data_i[16]
port 333 nsew signal input
rlabel metal2 s 19338 139200 19394 140000 6 io_motor_data_i[17]
port 334 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 io_motor_data_i[18]
port 335 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_motor_data_i[19]
port 336 nsew signal input
rlabel metal2 s 48962 139200 49018 140000 6 io_motor_data_i[1]
port 337 nsew signal input
rlabel metal3 s 139200 80928 140000 81048 6 io_motor_data_i[20]
port 338 nsew signal input
rlabel metal3 s 139200 133968 140000 134088 6 io_motor_data_i[21]
port 339 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 io_motor_data_i[22]
port 340 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 io_motor_data_i[23]
port 341 nsew signal input
rlabel metal3 s 139200 57128 140000 57248 6 io_motor_data_i[24]
port 342 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 io_motor_data_i[25]
port 343 nsew signal input
rlabel metal2 s 107566 139200 107622 140000 6 io_motor_data_i[26]
port 344 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 io_motor_data_i[27]
port 345 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 io_motor_data_i[28]
port 346 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_motor_data_i[29]
port 347 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 io_motor_data_i[2]
port 348 nsew signal input
rlabel metal3 s 139200 35368 140000 35488 6 io_motor_data_i[30]
port 349 nsew signal input
rlabel metal2 s 46386 139200 46442 140000 6 io_motor_data_i[31]
port 350 nsew signal input
rlabel metal3 s 139200 121728 140000 121848 6 io_motor_data_i[3]
port 351 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 io_motor_data_i[4]
port 352 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 io_motor_data_i[5]
port 353 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 io_motor_data_i[6]
port 354 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_motor_data_i[7]
port 355 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 io_motor_data_i[8]
port 356 nsew signal input
rlabel metal3 s 139200 71408 140000 71528 6 io_motor_data_i[9]
port 357 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 io_spi_clk
port 358 nsew signal output
rlabel metal2 s 95974 139200 96030 140000 6 io_spi_cs
port 359 nsew signal output
rlabel metal2 s 129462 139200 129518 140000 6 io_spi_irq
port 360 nsew signal output
rlabel metal2 s 10322 139200 10378 140000 6 io_spi_miso
port 361 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 io_spi_mosi
port 362 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 io_uart_irq
port 363 nsew signal output
rlabel metal2 s 133326 139200 133382 140000 6 io_uart_rx
port 364 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 io_uart_tx
port 365 nsew signal output
rlabel metal3 s 139200 109488 140000 109608 6 io_wbm_m2s_addr[0]
port 366 nsew signal output
rlabel metal3 s 139200 43528 140000 43648 6 io_wbm_m2s_addr[10]
port 367 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 io_wbm_m2s_addr[11]
port 368 nsew signal output
rlabel metal2 s 116582 139200 116638 140000 6 io_wbm_m2s_addr[12]
port 369 nsew signal output
rlabel metal2 s 36082 139200 36138 140000 6 io_wbm_m2s_addr[13]
port 370 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 io_wbm_m2s_addr[14]
port 371 nsew signal output
rlabel metal3 s 139200 83648 140000 83768 6 io_wbm_m2s_addr[15]
port 372 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 io_wbm_m2s_addr[1]
port 373 nsew signal output
rlabel metal3 s 139200 39448 140000 39568 6 io_wbm_m2s_addr[2]
port 374 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 io_wbm_m2s_addr[3]
port 375 nsew signal output
rlabel metal3 s 139200 1368 140000 1488 6 io_wbm_m2s_addr[4]
port 376 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_wbm_m2s_addr[5]
port 377 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 io_wbm_m2s_addr[6]
port 378 nsew signal output
rlabel metal3 s 139200 58488 140000 58608 6 io_wbm_m2s_addr[7]
port 379 nsew signal output
rlabel metal2 s 111430 139200 111486 140000 6 io_wbm_m2s_addr[8]
port 380 nsew signal output
rlabel metal3 s 139200 124448 140000 124568 6 io_wbm_m2s_addr[9]
port 381 nsew signal output
rlabel metal3 s 139200 4088 140000 4208 6 io_wbm_m2s_data[0]
port 382 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 io_wbm_m2s_data[10]
port 383 nsew signal output
rlabel metal3 s 139200 78208 140000 78328 6 io_wbm_m2s_data[11]
port 384 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 io_wbm_m2s_data[12]
port 385 nsew signal output
rlabel metal3 s 139200 128528 140000 128648 6 io_wbm_m2s_data[13]
port 386 nsew signal output
rlabel metal2 s 106278 139200 106334 140000 6 io_wbm_m2s_data[14]
port 387 nsew signal output
rlabel metal3 s 139200 13608 140000 13728 6 io_wbm_m2s_data[15]
port 388 nsew signal output
rlabel metal2 s 101126 139200 101182 140000 6 io_wbm_m2s_data[16]
port 389 nsew signal output
rlabel metal3 s 0 39448 800 39568 6 io_wbm_m2s_data[17]
port 390 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 io_wbm_m2s_data[18]
port 391 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 io_wbm_m2s_data[19]
port 392 nsew signal output
rlabel metal2 s 18 0 74 800 6 io_wbm_m2s_data[1]
port 393 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 io_wbm_m2s_data[20]
port 394 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 io_wbm_m2s_data[21]
port 395 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 io_wbm_m2s_data[22]
port 396 nsew signal output
rlabel metal2 s 41234 139200 41290 140000 6 io_wbm_m2s_data[23]
port 397 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 io_wbm_m2s_data[24]
port 398 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 io_wbm_m2s_data[25]
port 399 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 io_wbm_m2s_data[26]
port 400 nsew signal output
rlabel metal2 s 74078 139200 74134 140000 6 io_wbm_m2s_data[27]
port 401 nsew signal output
rlabel metal2 s 43810 139200 43866 140000 6 io_wbm_m2s_data[28]
port 402 nsew signal output
rlabel metal2 s 74078 0 74134 800 6 io_wbm_m2s_data[29]
port 403 nsew signal output
rlabel metal2 s 98550 139200 98606 140000 6 io_wbm_m2s_data[2]
port 404 nsew signal output
rlabel metal3 s 139200 36728 140000 36848 6 io_wbm_m2s_data[30]
port 405 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 io_wbm_m2s_data[31]
port 406 nsew signal output
rlabel metal3 s 139200 106768 140000 106888 6 io_wbm_m2s_data[3]
port 407 nsew signal output
rlabel metal2 s 29642 0 29698 800 6 io_wbm_m2s_data[4]
port 408 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 io_wbm_m2s_data[5]
port 409 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 io_wbm_m2s_data[6]
port 410 nsew signal output
rlabel metal3 s 139200 102688 140000 102808 6 io_wbm_m2s_data[7]
port 411 nsew signal output
rlabel metal2 s 83094 0 83150 800 6 io_wbm_m2s_data[8]
port 412 nsew signal output
rlabel metal2 s 93398 139200 93454 140000 6 io_wbm_m2s_data[9]
port 413 nsew signal output
rlabel metal2 s 92110 139200 92166 140000 6 io_wbm_m2s_sel[0]
port 414 nsew signal output
rlabel metal3 s 0 132608 800 132728 6 io_wbm_m2s_sel[1]
port 415 nsew signal output
rlabel metal2 s 18050 139200 18106 140000 6 io_wbm_m2s_sel[2]
port 416 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 io_wbm_m2s_sel[3]
port 417 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 io_wbm_m2s_stb
port 418 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 io_wbm_m2s_we
port 419 nsew signal output
rlabel metal3 s 139200 66648 140000 66768 6 reset
port 420 nsew signal input
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 421 nsew power input
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 422 nsew ground input
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 422 nsew ground input
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 422 nsew ground input
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 422 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 140000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11514086
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Wishbone_InterConnect/runs/Wishbone_InterConnect/results/finishing/WB_InterConnect.magic.gds
string GDS_START 843636
<< end >>

