VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WB_InterConnect
  CLASS BLOCK ;
  FOREIGN WB_InterConnect ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END clock
  PIN io_dbus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 68.040 1000.000 68.640 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 996.000 641.150 1000.000 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 853.440 1000.000 854.040 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 996.000 16.470 1000.000 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 0.000 934.170 4.000 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 996.000 280.510 1000.000 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 996.000 579.970 1000.000 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 469.240 1000.000 469.840 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 397.840 1000.000 398.440 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 965.640 1000.000 966.240 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 863.640 1000.000 864.240 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 996.000 792.490 1000.000 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 996.000 676.570 1000.000 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 574.640 1000.000 575.240 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 996.000 93.750 1000.000 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 996.000 995.350 1000.000 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 0.000 872.990 4.000 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 996.000 757.070 1000.000 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 996.000 950.270 1000.000 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 404.640 1000.000 405.240 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 996.000 22.910 1000.000 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 996.000 802.150 1000.000 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 996.000 473.710 1000.000 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 248.240 1000.000 248.840 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.840 4.000 942.440 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 996.000 377.110 1000.000 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 329.840 1000.000 330.440 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 714.040 1000.000 714.640 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 975.840 1000.000 976.440 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 0.000 908.410 4.000 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 996.000 87.310 1000.000 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 996.000 402.870 1000.000 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 996.000 174.250 1000.000 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 992.840 1000.000 993.440 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 115.640 1000.000 116.240 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 996.000 245.090 1000.000 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 996.000 853.670 1000.000 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 741.240 1000.000 741.840 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.570 996.000 914.850 1000.000 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 340.040 1000.000 340.640 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 996.000 396.430 1000.000 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 996.000 625.050 1000.000 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 489.640 1000.000 490.240 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 996.000 209.670 1000.000 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 996.000 77.650 1000.000 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 996.000 386.770 1000.000 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 996.000 879.430 1000.000 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 996.000 969.590 1000.000 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 955.440 1000.000 956.040 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 442.040 1000.000 442.640 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 826.240 1000.000 826.840 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 996.000 509.130 1000.000 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 996.000 361.010 1000.000 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 996.000 599.290 1000.000 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 778.640 1000.000 779.240 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 61.240 1000.000 61.840 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 996.000 534.890 1000.000 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 3.440 1000.000 4.040 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 996.000 544.550 1000.000 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 996.000 438.290 1000.000 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 142.840 1000.000 143.440 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 255.040 1000.000 255.640 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 367.240 1000.000 367.840 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 0.000 599.290 4.000 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 180.240 1000.000 180.840 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 387.640 1000.000 388.240 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 996.000 705.550 1000.000 ;
    END
  END io_dbus_wr_en
  PIN io_dmem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 302.640 1000.000 303.240 ;
    END
  END io_dmem_io_addr[0]
  PIN io_dmem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 210.840 1000.000 211.440 ;
    END
  END io_dmem_io_addr[1]
  PIN io_dmem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END io_dmem_io_addr[2]
  PIN io_dmem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END io_dmem_io_addr[3]
  PIN io_dmem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_dmem_io_addr[4]
  PIN io_dmem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END io_dmem_io_addr[5]
  PIN io_dmem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 78.240 1000.000 78.840 ;
    END
  END io_dmem_io_addr[6]
  PIN io_dmem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_dmem_io_addr[7]
  PIN io_dmem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 217.640 1000.000 218.240 ;
    END
  END io_dmem_io_rdata[0]
  PIN io_dmem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END io_dmem_io_rdata[10]
  PIN io_dmem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 105.440 1000.000 106.040 ;
    END
  END io_dmem_io_rdata[11]
  PIN io_dmem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 996.000 863.330 1000.000 ;
    END
  END io_dmem_io_rdata[12]
  PIN io_dmem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 23.840 1000.000 24.440 ;
    END
  END io_dmem_io_rdata[13]
  PIN io_dmem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 833.040 1000.000 833.640 ;
    END
  END io_dmem_io_rdata[14]
  PIN io_dmem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 996.000 164.590 1000.000 ;
    END
  END io_dmem_io_rdata[15]
  PIN io_dmem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END io_dmem_io_rdata[16]
  PIN io_dmem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 996.000 113.070 1000.000 ;
    END
  END io_dmem_io_rdata[17]
  PIN io_dmem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END io_dmem_io_rdata[18]
  PIN io_dmem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END io_dmem_io_rdata[19]
  PIN io_dmem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END io_dmem_io_rdata[1]
  PIN io_dmem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 676.640 1000.000 677.240 ;
    END
  END io_dmem_io_rdata[20]
  PIN io_dmem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END io_dmem_io_rdata[21]
  PIN io_dmem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 544.040 1000.000 544.640 ;
    END
  END io_dmem_io_rdata[22]
  PIN io_dmem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 996.000 138.830 1000.000 ;
    END
  END io_dmem_io_rdata[23]
  PIN io_dmem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END io_dmem_io_rdata[24]
  PIN io_dmem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_dmem_io_rdata[25]
  PIN io_dmem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 200.640 1000.000 201.240 ;
    END
  END io_dmem_io_rdata[26]
  PIN io_dmem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 163.240 1000.000 163.840 ;
    END
  END io_dmem_io_rdata[27]
  PIN io_dmem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 292.440 1000.000 293.040 ;
    END
  END io_dmem_io_rdata[28]
  PIN io_dmem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 996.000 58.330 1000.000 ;
    END
  END io_dmem_io_rdata[29]
  PIN io_dmem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END io_dmem_io_rdata[2]
  PIN io_dmem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_dmem_io_rdata[30]
  PIN io_dmem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 880.640 1000.000 881.240 ;
    END
  END io_dmem_io_rdata[31]
  PIN io_dmem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END io_dmem_io_rdata[3]
  PIN io_dmem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 996.000 563.870 1000.000 ;
    END
  END io_dmem_io_rdata[4]
  PIN io_dmem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 136.040 1000.000 136.640 ;
    END
  END io_dmem_io_rdata[5]
  PIN io_dmem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END io_dmem_io_rdata[6]
  PIN io_dmem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END io_dmem_io_rdata[7]
  PIN io_dmem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 996.000 341.690 1000.000 ;
    END
  END io_dmem_io_rdata[8]
  PIN io_dmem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 996.000 351.350 1000.000 ;
    END
  END io_dmem_io_rdata[9]
  PIN io_dmem_io_st_type[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END io_dmem_io_st_type[0]
  PIN io_dmem_io_st_type[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 996.000 605.730 1000.000 ;
    END
  END io_dmem_io_st_type[1]
  PIN io_dmem_io_st_type[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END io_dmem_io_st_type[2]
  PIN io_dmem_io_st_type[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END io_dmem_io_st_type[3]
  PIN io_dmem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 805.840 1000.000 806.440 ;
    END
  END io_dmem_io_wdata[0]
  PIN io_dmem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.240 4.000 690.840 ;
    END
  END io_dmem_io_wdata[10]
  PIN io_dmem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 350.240 1000.000 350.840 ;
    END
  END io_dmem_io_wdata[11]
  PIN io_dmem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_dmem_io_wdata[12]
  PIN io_dmem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 996.000 979.250 1000.000 ;
    END
  END io_dmem_io_wdata[13]
  PIN io_dmem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END io_dmem_io_wdata[14]
  PIN io_dmem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.970 0.000 979.250 4.000 ;
    END
  END io_dmem_io_wdata[15]
  PIN io_dmem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END io_dmem_io_wdata[16]
  PIN io_dmem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END io_dmem_io_wdata[17]
  PIN io_dmem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END io_dmem_io_wdata[18]
  PIN io_dmem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 788.840 1000.000 789.440 ;
    END
  END io_dmem_io_wdata[19]
  PIN io_dmem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END io_dmem_io_wdata[1]
  PIN io_dmem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END io_dmem_io_wdata[20]
  PIN io_dmem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 996.000 589.630 1000.000 ;
    END
  END io_dmem_io_wdata[21]
  PIN io_dmem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END io_dmem_io_wdata[22]
  PIN io_dmem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 996.000 412.530 1000.000 ;
    END
  END io_dmem_io_wdata[23]
  PIN io_dmem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_dmem_io_wdata[24]
  PIN io_dmem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END io_dmem_io_wdata[25]
  PIN io_dmem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 843.240 1000.000 843.840 ;
    END
  END io_dmem_io_wdata[26]
  PIN io_dmem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 996.000 570.310 1000.000 ;
    END
  END io_dmem_io_wdata[27]
  PIN io_dmem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END io_dmem_io_wdata[28]
  PIN io_dmem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END io_dmem_io_wdata[29]
  PIN io_dmem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END io_dmem_io_wdata[2]
  PIN io_dmem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 462.440 1000.000 463.040 ;
    END
  END io_dmem_io_wdata[30]
  PIN io_dmem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_dmem_io_wdata[31]
  PIN io_dmem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END io_dmem_io_wdata[3]
  PIN io_dmem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END io_dmem_io_wdata[4]
  PIN io_dmem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 751.440 1000.000 752.040 ;
    END
  END io_dmem_io_wdata[5]
  PIN io_dmem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 996.000 943.830 1000.000 ;
    END
  END io_dmem_io_wdata[6]
  PIN io_dmem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END io_dmem_io_wdata[7]
  PIN io_dmem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 996.000 325.590 1000.000 ;
    END
  END io_dmem_io_wdata[8]
  PIN io_dmem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END io_dmem_io_wdata[9]
  PIN io_dmem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 0.000 856.890 4.000 ;
    END
  END io_dmem_io_wr_en
  PIN io_ibus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END io_ibus_addr[0]
  PIN io_ibus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END io_ibus_addr[10]
  PIN io_ibus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 996.000 332.030 1000.000 ;
    END
  END io_ibus_addr[11]
  PIN io_ibus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 0.000 493.030 4.000 ;
    END
  END io_ibus_addr[12]
  PIN io_ibus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 435.240 1000.000 435.840 ;
    END
  END io_ibus_addr[13]
  PIN io_ibus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END io_ibus_addr[14]
  PIN io_ibus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 377.440 1000.000 378.040 ;
    END
  END io_ibus_addr[15]
  PIN io_ibus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_ibus_addr[16]
  PIN io_ibus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END io_ibus_addr[17]
  PIN io_ibus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END io_ibus_addr[18]
  PIN io_ibus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 996.000 225.770 1000.000 ;
    END
  END io_ibus_addr[19]
  PIN io_ibus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END io_ibus_addr[1]
  PIN io_ibus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_ibus_addr[20]
  PIN io_ibus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END io_ibus_addr[21]
  PIN io_ibus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END io_ibus_addr[22]
  PIN io_ibus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END io_ibus_addr[23]
  PIN io_ibus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 601.840 1000.000 602.440 ;
    END
  END io_ibus_addr[24]
  PIN io_ibus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END io_ibus_addr[25]
  PIN io_ibus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 996.000 889.090 1000.000 ;
    END
  END io_ibus_addr[26]
  PIN io_ibus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END io_ibus_addr[27]
  PIN io_ibus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 0.000 963.150 4.000 ;
    END
  END io_ibus_addr[28]
  PIN io_ibus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END io_ibus_addr[29]
  PIN io_ibus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 639.240 1000.000 639.840 ;
    END
  END io_ibus_addr[2]
  PIN io_ibus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 996.000 6.810 1000.000 ;
    END
  END io_ibus_addr[30]
  PIN io_ibus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END io_ibus_addr[31]
  PIN io_ibus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.650 996.000 959.930 1000.000 ;
    END
  END io_ibus_addr[3]
  PIN io_ibus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 499.840 1000.000 500.440 ;
    END
  END io_ibus_addr[4]
  PIN io_ibus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 4.000 ;
    END
  END io_ibus_addr[5]
  PIN io_ibus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 649.440 1000.000 650.040 ;
    END
  END io_ibus_addr[6]
  PIN io_ibus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 996.000 261.190 1000.000 ;
    END
  END io_ibus_addr[7]
  PIN io_ibus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 945.240 1000.000 945.840 ;
    END
  END io_ibus_addr[8]
  PIN io_ibus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END io_ibus_addr[9]
  PIN io_ibus_inst[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 996.000 493.030 1000.000 ;
    END
  END io_ibus_inst[0]
  PIN io_ibus_inst[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 190.440 1000.000 191.040 ;
    END
  END io_ibus_inst[10]
  PIN io_ibus_inst[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 816.040 1000.000 816.640 ;
    END
  END io_ibus_inst[11]
  PIN io_ibus_inst[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 724.240 1000.000 724.840 ;
    END
  END io_ibus_inst[12]
  PIN io_ibus_inst[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END io_ibus_inst[13]
  PIN io_ibus_inst[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 996.000 483.370 1000.000 ;
    END
  END io_ibus_inst[14]
  PIN io_ibus_inst[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 996.000 731.310 1000.000 ;
    END
  END io_ibus_inst[15]
  PIN io_ibus_inst[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 996.000 431.850 1000.000 ;
    END
  END io_ibus_inst[16]
  PIN io_ibus_inst[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_ibus_inst[17]
  PIN io_ibus_inst[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 996.000 296.610 1000.000 ;
    END
  END io_ibus_inst[18]
  PIN io_ibus_inst[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END io_ibus_inst[19]
  PIN io_ibus_inst[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END io_ibus_inst[1]
  PIN io_ibus_inst[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 996.000 148.490 1000.000 ;
    END
  END io_ibus_inst[20]
  PIN io_ibus_inst[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 996.000 740.970 1000.000 ;
    END
  END io_ibus_inst[21]
  PIN io_ibus_inst[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END io_ibus_inst[22]
  PIN io_ibus_inst[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 238.040 1000.000 238.640 ;
    END
  END io_ibus_inst[23]
  PIN io_ibus_inst[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END io_ibus_inst[24]
  PIN io_ibus_inst[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 996.000 457.610 1000.000 ;
    END
  END io_ibus_inst[25]
  PIN io_ibus_inst[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 907.840 1000.000 908.440 ;
    END
  END io_ibus_inst[26]
  PIN io_ibus_inst[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 452.240 1000.000 452.840 ;
    END
  END io_ibus_inst[27]
  PIN io_ibus_inst[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 51.040 1000.000 51.640 ;
    END
  END io_ibus_inst[28]
  PIN io_ibus_inst[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END io_ibus_inst[29]
  PIN io_ibus_inst[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END io_ibus_inst[2]
  PIN io_ibus_inst[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.290 0.000 998.570 4.000 ;
    END
  END io_ibus_inst[30]
  PIN io_ibus_inst[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.040 4.000 969.640 ;
    END
  END io_ibus_inst[31]
  PIN io_ibus_inst[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 938.440 1000.000 939.040 ;
    END
  END io_ibus_inst[3]
  PIN io_ibus_inst[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_ibus_inst[4]
  PIN io_ibus_inst[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END io_ibus_inst[5]
  PIN io_ibus_inst[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 996.000 518.790 1000.000 ;
    END
  END io_ibus_inst[6]
  PIN io_ibus_inst[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 996.000 42.230 1000.000 ;
    END
  END io_ibus_inst[7]
  PIN io_ibus_inst[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END io_ibus_inst[8]
  PIN io_ibus_inst[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END io_ibus_inst[9]
  PIN io_ibus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END io_ibus_valid
  PIN io_imem_io_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 581.440 1000.000 582.040 ;
    END
  END io_imem_io_addr[0]
  PIN io_imem_io_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 153.040 1000.000 153.640 ;
    END
  END io_imem_io_addr[10]
  PIN io_imem_io_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END io_imem_io_addr[11]
  PIN io_imem_io_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 88.440 1000.000 89.040 ;
    END
  END io_imem_io_addr[12]
  PIN io_imem_io_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 996.000 67.990 1000.000 ;
    END
  END io_imem_io_addr[13]
  PIN io_imem_io_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 996.000 686.230 1000.000 ;
    END
  END io_imem_io_addr[14]
  PIN io_imem_io_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END io_imem_io_addr[15]
  PIN io_imem_io_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 275.440 1000.000 276.040 ;
    END
  END io_imem_io_addr[16]
  PIN io_imem_io_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 996.000 467.270 1000.000 ;
    END
  END io_imem_io_addr[17]
  PIN io_imem_io_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END io_imem_io_addr[18]
  PIN io_imem_io_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END io_imem_io_addr[19]
  PIN io_imem_io_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 996.000 447.950 1000.000 ;
    END
  END io_imem_io_addr[1]
  PIN io_imem_io_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 996.000 721.650 1000.000 ;
    END
  END io_imem_io_addr[20]
  PIN io_imem_io_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END io_imem_io_addr[21]
  PIN io_imem_io_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END io_imem_io_addr[22]
  PIN io_imem_io_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 996.000 499.470 1000.000 ;
    END
  END io_imem_io_addr[23]
  PIN io_imem_io_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END io_imem_io_addr[24]
  PIN io_imem_io_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 996.000 872.990 1000.000 ;
    END
  END io_imem_io_addr[25]
  PIN io_imem_io_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END io_imem_io_addr[26]
  PIN io_imem_io_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END io_imem_io_addr[27]
  PIN io_imem_io_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 414.840 1000.000 415.440 ;
    END
  END io_imem_io_addr[28]
  PIN io_imem_io_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_imem_io_addr[29]
  PIN io_imem_io_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END io_imem_io_addr[2]
  PIN io_imem_io_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END io_imem_io_addr[30]
  PIN io_imem_io_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 629.040 1000.000 629.640 ;
    END
  END io_imem_io_addr[31]
  PIN io_imem_io_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END io_imem_io_addr[3]
  PIN io_imem_io_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END io_imem_io_addr[4]
  PIN io_imem_io_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END io_imem_io_addr[5]
  PIN io_imem_io_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END io_imem_io_addr[6]
  PIN io_imem_io_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_imem_io_addr[7]
  PIN io_imem_io_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 996.000 119.510 1000.000 ;
    END
  END io_imem_io_addr[8]
  PIN io_imem_io_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 554.240 1000.000 554.840 ;
    END
  END io_imem_io_addr[9]
  PIN io_imem_io_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 996.000 844.010 1000.000 ;
    END
  END io_imem_io_rdata[0]
  PIN io_imem_io_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 996.000 811.810 1000.000 ;
    END
  END io_imem_io_rdata[10]
  PIN io_imem_io_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_imem_io_rdata[11]
  PIN io_imem_io_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END io_imem_io_rdata[12]
  PIN io_imem_io_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 656.240 1000.000 656.840 ;
    END
  END io_imem_io_rdata[13]
  PIN io_imem_io_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 0.000 898.750 4.000 ;
    END
  END io_imem_io_rdata[14]
  PIN io_imem_io_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END io_imem_io_rdata[15]
  PIN io_imem_io_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END io_imem_io_rdata[16]
  PIN io_imem_io_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END io_imem_io_rdata[17]
  PIN io_imem_io_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 985.410 996.000 985.690 1000.000 ;
    END
  END io_imem_io_rdata[18]
  PIN io_imem_io_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.230 996.000 924.510 1000.000 ;
    END
  END io_imem_io_rdata[19]
  PIN io_imem_io_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 918.040 1000.000 918.640 ;
    END
  END io_imem_io_rdata[1]
  PIN io_imem_io_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 996.000 367.450 1000.000 ;
    END
  END io_imem_io_rdata[20]
  PIN io_imem_io_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 870.440 1000.000 871.040 ;
    END
  END io_imem_io_rdata[21]
  PIN io_imem_io_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END io_imem_io_rdata[22]
  PIN io_imem_io_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 996.000 827.910 1000.000 ;
    END
  END io_imem_io_rdata[23]
  PIN io_imem_io_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 996.000 183.910 1000.000 ;
    END
  END io_imem_io_rdata[24]
  PIN io_imem_io_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END io_imem_io_rdata[25]
  PIN io_imem_io_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 996.000 190.350 1000.000 ;
    END
  END io_imem_io_rdata[26]
  PIN io_imem_io_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END io_imem_io_rdata[27]
  PIN io_imem_io_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 40.840 1000.000 41.440 ;
    END
  END io_imem_io_rdata[28]
  PIN io_imem_io_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_imem_io_rdata[29]
  PIN io_imem_io_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 125.840 1000.000 126.440 ;
    END
  END io_imem_io_rdata[2]
  PIN io_imem_io_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.240 4.000 996.840 ;
    END
  END io_imem_io_rdata[30]
  PIN io_imem_io_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 615.440 4.000 616.040 ;
    END
  END io_imem_io_rdata[31]
  PIN io_imem_io_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END io_imem_io_rdata[3]
  PIN io_imem_io_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END io_imem_io_rdata[4]
  PIN io_imem_io_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 996.000 776.390 1000.000 ;
    END
  END io_imem_io_rdata[5]
  PIN io_imem_io_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END io_imem_io_rdata[6]
  PIN io_imem_io_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END io_imem_io_rdata[7]
  PIN io_imem_io_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END io_imem_io_rdata[8]
  PIN io_imem_io_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 506.640 1000.000 507.240 ;
    END
  END io_imem_io_rdata[9]
  PIN io_imem_io_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 703.840 1000.000 704.440 ;
    END
  END io_imem_io_wdata[0]
  PIN io_imem_io_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END io_imem_io_wdata[10]
  PIN io_imem_io_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 996.000 270.850 1000.000 ;
    END
  END io_imem_io_wdata[11]
  PIN io_imem_io_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io_imem_io_wdata[12]
  PIN io_imem_io_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 666.440 1000.000 667.040 ;
    END
  END io_imem_io_wdata[13]
  PIN io_imem_io_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END io_imem_io_wdata[14]
  PIN io_imem_io_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 537.240 1000.000 537.840 ;
    END
  END io_imem_io_wdata[15]
  PIN io_imem_io_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END io_imem_io_wdata[16]
  PIN io_imem_io_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 996.000 837.570 1000.000 ;
    END
  END io_imem_io_wdata[17]
  PIN io_imem_io_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END io_imem_io_wdata[18]
  PIN io_imem_io_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 996.000 554.210 1000.000 ;
    END
  END io_imem_io_wdata[19]
  PIN io_imem_io_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END io_imem_io_wdata[1]
  PIN io_imem_io_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 996.000 200.010 1000.000 ;
    END
  END io_imem_io_wdata[20]
  PIN io_imem_io_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_imem_io_wdata[21]
  PIN io_imem_io_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 516.840 1000.000 517.440 ;
    END
  END io_imem_io_wdata[22]
  PIN io_imem_io_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END io_imem_io_wdata[23]
  PIN io_imem_io_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 686.840 1000.000 687.440 ;
    END
  END io_imem_io_wdata[24]
  PIN io_imem_io_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END io_imem_io_wdata[25]
  PIN io_imem_io_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.550 0.000 943.830 4.000 ;
    END
  END io_imem_io_wdata[26]
  PIN io_imem_io_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 996.000 254.750 1000.000 ;
    END
  END io_imem_io_wdata[27]
  PIN io_imem_io_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END io_imem_io_wdata[28]
  PIN io_imem_io_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END io_imem_io_wdata[29]
  PIN io_imem_io_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 996.000 219.330 1000.000 ;
    END
  END io_imem_io_wdata[2]
  PIN io_imem_io_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_imem_io_wdata[30]
  PIN io_imem_io_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 173.440 1000.000 174.040 ;
    END
  END io_imem_io_wdata[31]
  PIN io_imem_io_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 996.000 154.930 1000.000 ;
    END
  END io_imem_io_wdata[3]
  PIN io_imem_io_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 360.440 1000.000 361.040 ;
    END
  END io_imem_io_wdata[4]
  PIN io_imem_io_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 996.000 634.710 1000.000 ;
    END
  END io_imem_io_wdata[5]
  PIN io_imem_io_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 996.000 422.190 1000.000 ;
    END
  END io_imem_io_wdata[6]
  PIN io_imem_io_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 996.000 32.570 1000.000 ;
    END
  END io_imem_io_wdata[7]
  PIN io_imem_io_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END io_imem_io_wdata[8]
  PIN io_imem_io_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END io_imem_io_wdata[9]
  PIN io_imem_io_wr_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 761.640 1000.000 762.240 ;
    END
  END io_imem_io_wr_en
  PIN io_motor_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 693.640 1000.000 694.240 ;
    END
  END io_motor_ack_i
  PIN io_motor_addr_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END io_motor_addr_sel
  PIN io_motor_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 618.840 1000.000 619.440 ;
    END
  END io_motor_data_i[0]
  PIN io_motor_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 312.840 1000.000 313.440 ;
    END
  END io_motor_data_i[10]
  PIN io_motor_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END io_motor_data_i[11]
  PIN io_motor_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 996.000 615.390 1000.000 ;
    END
  END io_motor_data_i[12]
  PIN io_motor_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.470 996.000 898.750 1000.000 ;
    END
  END io_motor_data_i[13]
  PIN io_motor_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END io_motor_data_i[14]
  PIN io_motor_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END io_motor_data_i[15]
  PIN io_motor_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 227.840 1000.000 228.440 ;
    END
  END io_motor_data_i[16]
  PIN io_motor_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 996.000 103.410 1000.000 ;
    END
  END io_motor_data_i[17]
  PIN io_motor_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END io_motor_data_i[18]
  PIN io_motor_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END io_motor_data_i[19]
  PIN io_motor_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 996.000 315.930 1000.000 ;
    END
  END io_motor_data_i[1]
  PIN io_motor_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 591.640 1000.000 592.240 ;
    END
  END io_motor_data_i[20]
  PIN io_motor_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 982.640 1000.000 983.240 ;
    END
  END io_motor_data_i[21]
  PIN io_motor_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END io_motor_data_i[22]
  PIN io_motor_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 996.000 766.730 1000.000 ;
    END
  END io_motor_data_i[23]
  PIN io_motor_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END io_motor_data_i[24]
  PIN io_motor_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END io_motor_data_i[25]
  PIN io_motor_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END io_motor_data_i[26]
  PIN io_motor_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END io_motor_data_i[27]
  PIN io_motor_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END io_motor_data_i[28]
  PIN io_motor_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_motor_data_i[29]
  PIN io_motor_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 0.000 988.910 4.000 ;
    END
  END io_motor_data_i[2]
  PIN io_motor_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_motor_data_i[30]
  PIN io_motor_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_motor_data_i[31]
  PIN io_motor_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 890.840 1000.000 891.440 ;
    END
  END io_motor_data_i[3]
  PIN io_motor_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END io_motor_data_i[4]
  PIN io_motor_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END io_motor_data_i[5]
  PIN io_motor_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END io_motor_data_i[6]
  PIN io_motor_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_motor_data_i[7]
  PIN io_motor_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_motor_data_i[8]
  PIN io_motor_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 527.040 1000.000 527.640 ;
    END
  END io_motor_data_i[9]
  PIN io_spi_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END io_spi_clk
  PIN io_spi_cs
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 996.000 670.130 1000.000 ;
    END
  END io_spi_cs
  PIN io_spi_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 996.000 908.410 1000.000 ;
    END
  END io_spi_irq
  PIN io_spi_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 996.000 51.890 1000.000 ;
    END
  END io_spi_miso
  PIN io_spi_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_spi_mosi
  PIN io_uart_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END io_uart_irq
  PIN io_uart_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.890 996.000 934.170 1000.000 ;
    END
  END io_uart_rx
  PIN io_uart_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END io_uart_tx
  PIN io_wbm_m2s_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 799.040 1000.000 799.640 ;
    END
  END io_wbm_m2s_addr[0]
  PIN io_wbm_m2s_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 323.040 1000.000 323.640 ;
    END
  END io_wbm_m2s_addr[10]
  PIN io_wbm_m2s_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END io_wbm_m2s_addr[11]
  PIN io_wbm_m2s_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 996.000 818.250 1000.000 ;
    END
  END io_wbm_m2s_addr[12]
  PIN io_wbm_m2s_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 996.000 235.430 1000.000 ;
    END
  END io_wbm_m2s_addr[13]
  PIN io_wbm_m2s_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_wbm_m2s_addr[14]
  PIN io_wbm_m2s_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 612.040 1000.000 612.640 ;
    END
  END io_wbm_m2s_addr[15]
  PIN io_wbm_m2s_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END io_wbm_m2s_addr[1]
  PIN io_wbm_m2s_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 285.640 1000.000 286.240 ;
    END
  END io_wbm_m2s_addr[2]
  PIN io_wbm_m2s_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_wbm_m2s_addr[3]
  PIN io_wbm_m2s_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 13.640 1000.000 14.240 ;
    END
  END io_wbm_m2s_addr[4]
  PIN io_wbm_m2s_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_wbm_m2s_addr[5]
  PIN io_wbm_m2s_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END io_wbm_m2s_addr[6]
  PIN io_wbm_m2s_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 425.040 1000.000 425.640 ;
    END
  END io_wbm_m2s_addr[7]
  PIN io_wbm_m2s_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 996.000 782.830 1000.000 ;
    END
  END io_wbm_m2s_addr[8]
  PIN io_wbm_m2s_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 901.040 1000.000 901.640 ;
    END
  END io_wbm_m2s_addr[9]
  PIN io_wbm_m2s_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 34.040 1000.000 34.640 ;
    END
  END io_wbm_m2s_data[0]
  PIN io_wbm_m2s_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END io_wbm_m2s_data[10]
  PIN io_wbm_m2s_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 564.440 1000.000 565.040 ;
    END
  END io_wbm_m2s_data[11]
  PIN io_wbm_m2s_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_wbm_m2s_data[12]
  PIN io_wbm_m2s_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 928.240 1000.000 928.840 ;
    END
  END io_wbm_m2s_data[13]
  PIN io_wbm_m2s_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 996.000 747.410 1000.000 ;
    END
  END io_wbm_m2s_data[14]
  PIN io_wbm_m2s_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 98.640 1000.000 99.240 ;
    END
  END io_wbm_m2s_data[15]
  PIN io_wbm_m2s_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 996.000 711.990 1000.000 ;
    END
  END io_wbm_m2s_data[16]
  PIN io_wbm_m2s_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END io_wbm_m2s_data[17]
  PIN io_wbm_m2s_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_wbm_m2s_data[18]
  PIN io_wbm_m2s_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 0.000 660.470 4.000 ;
    END
  END io_wbm_m2s_data[19]
  PIN io_wbm_m2s_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_wbm_m2s_data[1]
  PIN io_wbm_m2s_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END io_wbm_m2s_data[20]
  PIN io_wbm_m2s_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END io_wbm_m2s_data[21]
  PIN io_wbm_m2s_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END io_wbm_m2s_data[22]
  PIN io_wbm_m2s_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 996.000 290.170 1000.000 ;
    END
  END io_wbm_m2s_data[23]
  PIN io_wbm_m2s_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END io_wbm_m2s_data[24]
  PIN io_wbm_m2s_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END io_wbm_m2s_data[25]
  PIN io_wbm_m2s_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_wbm_m2s_data[26]
  PIN io_wbm_m2s_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 996.000 528.450 1000.000 ;
    END
  END io_wbm_m2s_data[27]
  PIN io_wbm_m2s_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 996.000 306.270 1000.000 ;
    END
  END io_wbm_m2s_data[28]
  PIN io_wbm_m2s_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END io_wbm_m2s_data[29]
  PIN io_wbm_m2s_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 996.000 695.890 1000.000 ;
    END
  END io_wbm_m2s_data[2]
  PIN io_wbm_m2s_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 265.240 1000.000 265.840 ;
    END
  END io_wbm_m2s_data[30]
  PIN io_wbm_m2s_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 669.840 4.000 670.440 ;
    END
  END io_wbm_m2s_data[31]
  PIN io_wbm_m2s_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 768.440 1000.000 769.040 ;
    END
  END io_wbm_m2s_data[3]
  PIN io_wbm_m2s_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END io_wbm_m2s_data[4]
  PIN io_wbm_m2s_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END io_wbm_m2s_data[5]
  PIN io_wbm_m2s_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_wbm_m2s_data[6]
  PIN io_wbm_m2s_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 731.040 1000.000 731.640 ;
    END
  END io_wbm_m2s_data[7]
  PIN io_wbm_m2s_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END io_wbm_m2s_data[8]
  PIN io_wbm_m2s_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 996.000 660.470 1000.000 ;
    END
  END io_wbm_m2s_data[9]
  PIN io_wbm_m2s_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 996.000 650.810 1000.000 ;
    END
  END io_wbm_m2s_sel[0]
  PIN io_wbm_m2s_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 948.640 4.000 949.240 ;
    END
  END io_wbm_m2s_sel[1]
  PIN io_wbm_m2s_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 996.000 129.170 1000.000 ;
    END
  END io_wbm_m2s_sel[2]
  PIN io_wbm_m2s_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END io_wbm_m2s_sel[3]
  PIN io_wbm_m2s_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END io_wbm_m2s_stb
  PIN io_wbm_m2s_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END io_wbm_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 479.440 1000.000 480.040 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 987.600 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 987.445 ;
      LAYER met1 ;
        RECT 0.070 9.220 998.590 988.340 ;
      LAYER met2 ;
        RECT 0.100 995.720 6.250 996.725 ;
        RECT 7.090 995.720 15.910 996.725 ;
        RECT 16.750 995.720 22.350 996.725 ;
        RECT 23.190 995.720 32.010 996.725 ;
        RECT 32.850 995.720 41.670 996.725 ;
        RECT 42.510 995.720 51.330 996.725 ;
        RECT 52.170 995.720 57.770 996.725 ;
        RECT 58.610 995.720 67.430 996.725 ;
        RECT 68.270 995.720 77.090 996.725 ;
        RECT 77.930 995.720 86.750 996.725 ;
        RECT 87.590 995.720 93.190 996.725 ;
        RECT 94.030 995.720 102.850 996.725 ;
        RECT 103.690 995.720 112.510 996.725 ;
        RECT 113.350 995.720 118.950 996.725 ;
        RECT 119.790 995.720 128.610 996.725 ;
        RECT 129.450 995.720 138.270 996.725 ;
        RECT 139.110 995.720 147.930 996.725 ;
        RECT 148.770 995.720 154.370 996.725 ;
        RECT 155.210 995.720 164.030 996.725 ;
        RECT 164.870 995.720 173.690 996.725 ;
        RECT 174.530 995.720 183.350 996.725 ;
        RECT 184.190 995.720 189.790 996.725 ;
        RECT 190.630 995.720 199.450 996.725 ;
        RECT 200.290 995.720 209.110 996.725 ;
        RECT 209.950 995.720 218.770 996.725 ;
        RECT 219.610 995.720 225.210 996.725 ;
        RECT 226.050 995.720 234.870 996.725 ;
        RECT 235.710 995.720 244.530 996.725 ;
        RECT 245.370 995.720 254.190 996.725 ;
        RECT 255.030 995.720 260.630 996.725 ;
        RECT 261.470 995.720 270.290 996.725 ;
        RECT 271.130 995.720 279.950 996.725 ;
        RECT 280.790 995.720 289.610 996.725 ;
        RECT 290.450 995.720 296.050 996.725 ;
        RECT 296.890 995.720 305.710 996.725 ;
        RECT 306.550 995.720 315.370 996.725 ;
        RECT 316.210 995.720 325.030 996.725 ;
        RECT 325.870 995.720 331.470 996.725 ;
        RECT 332.310 995.720 341.130 996.725 ;
        RECT 341.970 995.720 350.790 996.725 ;
        RECT 351.630 995.720 360.450 996.725 ;
        RECT 361.290 995.720 366.890 996.725 ;
        RECT 367.730 995.720 376.550 996.725 ;
        RECT 377.390 995.720 386.210 996.725 ;
        RECT 387.050 995.720 395.870 996.725 ;
        RECT 396.710 995.720 402.310 996.725 ;
        RECT 403.150 995.720 411.970 996.725 ;
        RECT 412.810 995.720 421.630 996.725 ;
        RECT 422.470 995.720 431.290 996.725 ;
        RECT 432.130 995.720 437.730 996.725 ;
        RECT 438.570 995.720 447.390 996.725 ;
        RECT 448.230 995.720 457.050 996.725 ;
        RECT 457.890 995.720 466.710 996.725 ;
        RECT 467.550 995.720 473.150 996.725 ;
        RECT 473.990 995.720 482.810 996.725 ;
        RECT 483.650 995.720 492.470 996.725 ;
        RECT 493.310 995.720 498.910 996.725 ;
        RECT 499.750 995.720 508.570 996.725 ;
        RECT 509.410 995.720 518.230 996.725 ;
        RECT 519.070 995.720 527.890 996.725 ;
        RECT 528.730 995.720 534.330 996.725 ;
        RECT 535.170 995.720 543.990 996.725 ;
        RECT 544.830 995.720 553.650 996.725 ;
        RECT 554.490 995.720 563.310 996.725 ;
        RECT 564.150 995.720 569.750 996.725 ;
        RECT 570.590 995.720 579.410 996.725 ;
        RECT 580.250 995.720 589.070 996.725 ;
        RECT 589.910 995.720 598.730 996.725 ;
        RECT 599.570 995.720 605.170 996.725 ;
        RECT 606.010 995.720 614.830 996.725 ;
        RECT 615.670 995.720 624.490 996.725 ;
        RECT 625.330 995.720 634.150 996.725 ;
        RECT 634.990 995.720 640.590 996.725 ;
        RECT 641.430 995.720 650.250 996.725 ;
        RECT 651.090 995.720 659.910 996.725 ;
        RECT 660.750 995.720 669.570 996.725 ;
        RECT 670.410 995.720 676.010 996.725 ;
        RECT 676.850 995.720 685.670 996.725 ;
        RECT 686.510 995.720 695.330 996.725 ;
        RECT 696.170 995.720 704.990 996.725 ;
        RECT 705.830 995.720 711.430 996.725 ;
        RECT 712.270 995.720 721.090 996.725 ;
        RECT 721.930 995.720 730.750 996.725 ;
        RECT 731.590 995.720 740.410 996.725 ;
        RECT 741.250 995.720 746.850 996.725 ;
        RECT 747.690 995.720 756.510 996.725 ;
        RECT 757.350 995.720 766.170 996.725 ;
        RECT 767.010 995.720 775.830 996.725 ;
        RECT 776.670 995.720 782.270 996.725 ;
        RECT 783.110 995.720 791.930 996.725 ;
        RECT 792.770 995.720 801.590 996.725 ;
        RECT 802.430 995.720 811.250 996.725 ;
        RECT 812.090 995.720 817.690 996.725 ;
        RECT 818.530 995.720 827.350 996.725 ;
        RECT 828.190 995.720 837.010 996.725 ;
        RECT 837.850 995.720 843.450 996.725 ;
        RECT 844.290 995.720 853.110 996.725 ;
        RECT 853.950 995.720 862.770 996.725 ;
        RECT 863.610 995.720 872.430 996.725 ;
        RECT 873.270 995.720 878.870 996.725 ;
        RECT 879.710 995.720 888.530 996.725 ;
        RECT 889.370 995.720 898.190 996.725 ;
        RECT 899.030 995.720 907.850 996.725 ;
        RECT 908.690 995.720 914.290 996.725 ;
        RECT 915.130 995.720 923.950 996.725 ;
        RECT 924.790 995.720 933.610 996.725 ;
        RECT 934.450 995.720 943.270 996.725 ;
        RECT 944.110 995.720 949.710 996.725 ;
        RECT 950.550 995.720 959.370 996.725 ;
        RECT 960.210 995.720 969.030 996.725 ;
        RECT 969.870 995.720 978.690 996.725 ;
        RECT 979.530 995.720 985.130 996.725 ;
        RECT 985.970 995.720 994.790 996.725 ;
        RECT 995.630 995.720 998.560 996.725 ;
        RECT 0.100 4.280 998.560 995.720 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 15.910 4.280 ;
        RECT 16.750 3.555 25.570 4.280 ;
        RECT 26.410 3.555 32.010 4.280 ;
        RECT 32.850 3.555 41.670 4.280 ;
        RECT 42.510 3.555 51.330 4.280 ;
        RECT 52.170 3.555 60.990 4.280 ;
        RECT 61.830 3.555 67.430 4.280 ;
        RECT 68.270 3.555 77.090 4.280 ;
        RECT 77.930 3.555 86.750 4.280 ;
        RECT 87.590 3.555 96.410 4.280 ;
        RECT 97.250 3.555 102.850 4.280 ;
        RECT 103.690 3.555 112.510 4.280 ;
        RECT 113.350 3.555 122.170 4.280 ;
        RECT 123.010 3.555 131.830 4.280 ;
        RECT 132.670 3.555 138.270 4.280 ;
        RECT 139.110 3.555 147.930 4.280 ;
        RECT 148.770 3.555 157.590 4.280 ;
        RECT 158.430 3.555 167.250 4.280 ;
        RECT 168.090 3.555 173.690 4.280 ;
        RECT 174.530 3.555 183.350 4.280 ;
        RECT 184.190 3.555 193.010 4.280 ;
        RECT 193.850 3.555 202.670 4.280 ;
        RECT 203.510 3.555 209.110 4.280 ;
        RECT 209.950 3.555 218.770 4.280 ;
        RECT 219.610 3.555 228.430 4.280 ;
        RECT 229.270 3.555 238.090 4.280 ;
        RECT 238.930 3.555 244.530 4.280 ;
        RECT 245.370 3.555 254.190 4.280 ;
        RECT 255.030 3.555 263.850 4.280 ;
        RECT 264.690 3.555 273.510 4.280 ;
        RECT 274.350 3.555 279.950 4.280 ;
        RECT 280.790 3.555 289.610 4.280 ;
        RECT 290.450 3.555 299.270 4.280 ;
        RECT 300.110 3.555 308.930 4.280 ;
        RECT 309.770 3.555 315.370 4.280 ;
        RECT 316.210 3.555 325.030 4.280 ;
        RECT 325.870 3.555 334.690 4.280 ;
        RECT 335.530 3.555 344.350 4.280 ;
        RECT 345.190 3.555 350.790 4.280 ;
        RECT 351.630 3.555 360.450 4.280 ;
        RECT 361.290 3.555 370.110 4.280 ;
        RECT 370.950 3.555 376.550 4.280 ;
        RECT 377.390 3.555 386.210 4.280 ;
        RECT 387.050 3.555 395.870 4.280 ;
        RECT 396.710 3.555 405.530 4.280 ;
        RECT 406.370 3.555 411.970 4.280 ;
        RECT 412.810 3.555 421.630 4.280 ;
        RECT 422.470 3.555 431.290 4.280 ;
        RECT 432.130 3.555 440.950 4.280 ;
        RECT 441.790 3.555 447.390 4.280 ;
        RECT 448.230 3.555 457.050 4.280 ;
        RECT 457.890 3.555 466.710 4.280 ;
        RECT 467.550 3.555 476.370 4.280 ;
        RECT 477.210 3.555 482.810 4.280 ;
        RECT 483.650 3.555 492.470 4.280 ;
        RECT 493.310 3.555 502.130 4.280 ;
        RECT 502.970 3.555 511.790 4.280 ;
        RECT 512.630 3.555 518.230 4.280 ;
        RECT 519.070 3.555 527.890 4.280 ;
        RECT 528.730 3.555 537.550 4.280 ;
        RECT 538.390 3.555 547.210 4.280 ;
        RECT 548.050 3.555 553.650 4.280 ;
        RECT 554.490 3.555 563.310 4.280 ;
        RECT 564.150 3.555 572.970 4.280 ;
        RECT 573.810 3.555 582.630 4.280 ;
        RECT 583.470 3.555 589.070 4.280 ;
        RECT 589.910 3.555 598.730 4.280 ;
        RECT 599.570 3.555 608.390 4.280 ;
        RECT 609.230 3.555 618.050 4.280 ;
        RECT 618.890 3.555 624.490 4.280 ;
        RECT 625.330 3.555 634.150 4.280 ;
        RECT 634.990 3.555 643.810 4.280 ;
        RECT 644.650 3.555 653.470 4.280 ;
        RECT 654.310 3.555 659.910 4.280 ;
        RECT 660.750 3.555 669.570 4.280 ;
        RECT 670.410 3.555 679.230 4.280 ;
        RECT 680.070 3.555 688.890 4.280 ;
        RECT 689.730 3.555 695.330 4.280 ;
        RECT 696.170 3.555 704.990 4.280 ;
        RECT 705.830 3.555 714.650 4.280 ;
        RECT 715.490 3.555 721.090 4.280 ;
        RECT 721.930 3.555 730.750 4.280 ;
        RECT 731.590 3.555 740.410 4.280 ;
        RECT 741.250 3.555 750.070 4.280 ;
        RECT 750.910 3.555 756.510 4.280 ;
        RECT 757.350 3.555 766.170 4.280 ;
        RECT 767.010 3.555 775.830 4.280 ;
        RECT 776.670 3.555 785.490 4.280 ;
        RECT 786.330 3.555 791.930 4.280 ;
        RECT 792.770 3.555 801.590 4.280 ;
        RECT 802.430 3.555 811.250 4.280 ;
        RECT 812.090 3.555 820.910 4.280 ;
        RECT 821.750 3.555 827.350 4.280 ;
        RECT 828.190 3.555 837.010 4.280 ;
        RECT 837.850 3.555 846.670 4.280 ;
        RECT 847.510 3.555 856.330 4.280 ;
        RECT 857.170 3.555 862.770 4.280 ;
        RECT 863.610 3.555 872.430 4.280 ;
        RECT 873.270 3.555 882.090 4.280 ;
        RECT 882.930 3.555 891.750 4.280 ;
        RECT 892.590 3.555 898.190 4.280 ;
        RECT 899.030 3.555 907.850 4.280 ;
        RECT 908.690 3.555 917.510 4.280 ;
        RECT 918.350 3.555 927.170 4.280 ;
        RECT 928.010 3.555 933.610 4.280 ;
        RECT 934.450 3.555 943.270 4.280 ;
        RECT 944.110 3.555 952.930 4.280 ;
        RECT 953.770 3.555 962.590 4.280 ;
        RECT 963.430 3.555 969.030 4.280 ;
        RECT 969.870 3.555 978.690 4.280 ;
        RECT 979.530 3.555 988.350 4.280 ;
        RECT 989.190 3.555 998.010 4.280 ;
      LAYER met3 ;
        RECT 4.400 995.840 996.000 996.705 ;
        RECT 4.000 993.840 996.000 995.840 ;
        RECT 4.000 992.440 995.600 993.840 ;
        RECT 4.000 987.040 996.000 992.440 ;
        RECT 4.400 985.640 996.000 987.040 ;
        RECT 4.000 983.640 996.000 985.640 ;
        RECT 4.000 982.240 995.600 983.640 ;
        RECT 4.000 980.240 996.000 982.240 ;
        RECT 4.400 978.840 996.000 980.240 ;
        RECT 4.000 976.840 996.000 978.840 ;
        RECT 4.000 975.440 995.600 976.840 ;
        RECT 4.000 970.040 996.000 975.440 ;
        RECT 4.400 968.640 996.000 970.040 ;
        RECT 4.000 966.640 996.000 968.640 ;
        RECT 4.000 965.240 995.600 966.640 ;
        RECT 4.000 959.840 996.000 965.240 ;
        RECT 4.400 958.440 996.000 959.840 ;
        RECT 4.000 956.440 996.000 958.440 ;
        RECT 4.000 955.040 995.600 956.440 ;
        RECT 4.000 949.640 996.000 955.040 ;
        RECT 4.400 948.240 996.000 949.640 ;
        RECT 4.000 946.240 996.000 948.240 ;
        RECT 4.000 944.840 995.600 946.240 ;
        RECT 4.000 942.840 996.000 944.840 ;
        RECT 4.400 941.440 996.000 942.840 ;
        RECT 4.000 939.440 996.000 941.440 ;
        RECT 4.000 938.040 995.600 939.440 ;
        RECT 4.000 932.640 996.000 938.040 ;
        RECT 4.400 931.240 996.000 932.640 ;
        RECT 4.000 929.240 996.000 931.240 ;
        RECT 4.000 927.840 995.600 929.240 ;
        RECT 4.000 922.440 996.000 927.840 ;
        RECT 4.400 921.040 996.000 922.440 ;
        RECT 4.000 919.040 996.000 921.040 ;
        RECT 4.000 917.640 995.600 919.040 ;
        RECT 4.000 912.240 996.000 917.640 ;
        RECT 4.400 910.840 996.000 912.240 ;
        RECT 4.000 908.840 996.000 910.840 ;
        RECT 4.000 907.440 995.600 908.840 ;
        RECT 4.000 905.440 996.000 907.440 ;
        RECT 4.400 904.040 996.000 905.440 ;
        RECT 4.000 902.040 996.000 904.040 ;
        RECT 4.000 900.640 995.600 902.040 ;
        RECT 4.000 895.240 996.000 900.640 ;
        RECT 4.400 893.840 996.000 895.240 ;
        RECT 4.000 891.840 996.000 893.840 ;
        RECT 4.000 890.440 995.600 891.840 ;
        RECT 4.000 885.040 996.000 890.440 ;
        RECT 4.400 883.640 996.000 885.040 ;
        RECT 4.000 881.640 996.000 883.640 ;
        RECT 4.000 880.240 995.600 881.640 ;
        RECT 4.000 874.840 996.000 880.240 ;
        RECT 4.400 873.440 996.000 874.840 ;
        RECT 4.000 871.440 996.000 873.440 ;
        RECT 4.000 870.040 995.600 871.440 ;
        RECT 4.000 868.040 996.000 870.040 ;
        RECT 4.400 866.640 996.000 868.040 ;
        RECT 4.000 864.640 996.000 866.640 ;
        RECT 4.000 863.240 995.600 864.640 ;
        RECT 4.000 857.840 996.000 863.240 ;
        RECT 4.400 856.440 996.000 857.840 ;
        RECT 4.000 854.440 996.000 856.440 ;
        RECT 4.000 853.040 995.600 854.440 ;
        RECT 4.000 847.640 996.000 853.040 ;
        RECT 4.400 846.240 996.000 847.640 ;
        RECT 4.000 844.240 996.000 846.240 ;
        RECT 4.000 842.840 995.600 844.240 ;
        RECT 4.000 837.440 996.000 842.840 ;
        RECT 4.400 836.040 996.000 837.440 ;
        RECT 4.000 834.040 996.000 836.040 ;
        RECT 4.000 832.640 995.600 834.040 ;
        RECT 4.000 830.640 996.000 832.640 ;
        RECT 4.400 829.240 996.000 830.640 ;
        RECT 4.000 827.240 996.000 829.240 ;
        RECT 4.000 825.840 995.600 827.240 ;
        RECT 4.000 820.440 996.000 825.840 ;
        RECT 4.400 819.040 996.000 820.440 ;
        RECT 4.000 817.040 996.000 819.040 ;
        RECT 4.000 815.640 995.600 817.040 ;
        RECT 4.000 810.240 996.000 815.640 ;
        RECT 4.400 808.840 996.000 810.240 ;
        RECT 4.000 806.840 996.000 808.840 ;
        RECT 4.000 805.440 995.600 806.840 ;
        RECT 4.000 800.040 996.000 805.440 ;
        RECT 4.400 798.640 995.600 800.040 ;
        RECT 4.000 793.240 996.000 798.640 ;
        RECT 4.400 791.840 996.000 793.240 ;
        RECT 4.000 789.840 996.000 791.840 ;
        RECT 4.000 788.440 995.600 789.840 ;
        RECT 4.000 783.040 996.000 788.440 ;
        RECT 4.400 781.640 996.000 783.040 ;
        RECT 4.000 779.640 996.000 781.640 ;
        RECT 4.000 778.240 995.600 779.640 ;
        RECT 4.000 772.840 996.000 778.240 ;
        RECT 4.400 771.440 996.000 772.840 ;
        RECT 4.000 769.440 996.000 771.440 ;
        RECT 4.000 768.040 995.600 769.440 ;
        RECT 4.000 762.640 996.000 768.040 ;
        RECT 4.400 761.240 995.600 762.640 ;
        RECT 4.000 755.840 996.000 761.240 ;
        RECT 4.400 754.440 996.000 755.840 ;
        RECT 4.000 752.440 996.000 754.440 ;
        RECT 4.000 751.040 995.600 752.440 ;
        RECT 4.000 745.640 996.000 751.040 ;
        RECT 4.400 744.240 996.000 745.640 ;
        RECT 4.000 742.240 996.000 744.240 ;
        RECT 4.000 740.840 995.600 742.240 ;
        RECT 4.000 735.440 996.000 740.840 ;
        RECT 4.400 734.040 996.000 735.440 ;
        RECT 4.000 732.040 996.000 734.040 ;
        RECT 4.000 730.640 995.600 732.040 ;
        RECT 4.000 728.640 996.000 730.640 ;
        RECT 4.400 727.240 996.000 728.640 ;
        RECT 4.000 725.240 996.000 727.240 ;
        RECT 4.000 723.840 995.600 725.240 ;
        RECT 4.000 718.440 996.000 723.840 ;
        RECT 4.400 717.040 996.000 718.440 ;
        RECT 4.000 715.040 996.000 717.040 ;
        RECT 4.000 713.640 995.600 715.040 ;
        RECT 4.000 708.240 996.000 713.640 ;
        RECT 4.400 706.840 996.000 708.240 ;
        RECT 4.000 704.840 996.000 706.840 ;
        RECT 4.000 703.440 995.600 704.840 ;
        RECT 4.000 698.040 996.000 703.440 ;
        RECT 4.400 696.640 996.000 698.040 ;
        RECT 4.000 694.640 996.000 696.640 ;
        RECT 4.000 693.240 995.600 694.640 ;
        RECT 4.000 691.240 996.000 693.240 ;
        RECT 4.400 689.840 996.000 691.240 ;
        RECT 4.000 687.840 996.000 689.840 ;
        RECT 4.000 686.440 995.600 687.840 ;
        RECT 4.000 681.040 996.000 686.440 ;
        RECT 4.400 679.640 996.000 681.040 ;
        RECT 4.000 677.640 996.000 679.640 ;
        RECT 4.000 676.240 995.600 677.640 ;
        RECT 4.000 670.840 996.000 676.240 ;
        RECT 4.400 669.440 996.000 670.840 ;
        RECT 4.000 667.440 996.000 669.440 ;
        RECT 4.000 666.040 995.600 667.440 ;
        RECT 4.000 660.640 996.000 666.040 ;
        RECT 4.400 659.240 996.000 660.640 ;
        RECT 4.000 657.240 996.000 659.240 ;
        RECT 4.000 655.840 995.600 657.240 ;
        RECT 4.000 653.840 996.000 655.840 ;
        RECT 4.400 652.440 996.000 653.840 ;
        RECT 4.000 650.440 996.000 652.440 ;
        RECT 4.000 649.040 995.600 650.440 ;
        RECT 4.000 643.640 996.000 649.040 ;
        RECT 4.400 642.240 996.000 643.640 ;
        RECT 4.000 640.240 996.000 642.240 ;
        RECT 4.000 638.840 995.600 640.240 ;
        RECT 4.000 633.440 996.000 638.840 ;
        RECT 4.400 632.040 996.000 633.440 ;
        RECT 4.000 630.040 996.000 632.040 ;
        RECT 4.000 628.640 995.600 630.040 ;
        RECT 4.000 623.240 996.000 628.640 ;
        RECT 4.400 621.840 996.000 623.240 ;
        RECT 4.000 619.840 996.000 621.840 ;
        RECT 4.000 618.440 995.600 619.840 ;
        RECT 4.000 616.440 996.000 618.440 ;
        RECT 4.400 615.040 996.000 616.440 ;
        RECT 4.000 613.040 996.000 615.040 ;
        RECT 4.000 611.640 995.600 613.040 ;
        RECT 4.000 606.240 996.000 611.640 ;
        RECT 4.400 604.840 996.000 606.240 ;
        RECT 4.000 602.840 996.000 604.840 ;
        RECT 4.000 601.440 995.600 602.840 ;
        RECT 4.000 596.040 996.000 601.440 ;
        RECT 4.400 594.640 996.000 596.040 ;
        RECT 4.000 592.640 996.000 594.640 ;
        RECT 4.000 591.240 995.600 592.640 ;
        RECT 4.000 585.840 996.000 591.240 ;
        RECT 4.400 584.440 996.000 585.840 ;
        RECT 4.000 582.440 996.000 584.440 ;
        RECT 4.000 581.040 995.600 582.440 ;
        RECT 4.000 579.040 996.000 581.040 ;
        RECT 4.400 577.640 996.000 579.040 ;
        RECT 4.000 575.640 996.000 577.640 ;
        RECT 4.000 574.240 995.600 575.640 ;
        RECT 4.000 568.840 996.000 574.240 ;
        RECT 4.400 567.440 996.000 568.840 ;
        RECT 4.000 565.440 996.000 567.440 ;
        RECT 4.000 564.040 995.600 565.440 ;
        RECT 4.000 558.640 996.000 564.040 ;
        RECT 4.400 557.240 996.000 558.640 ;
        RECT 4.000 555.240 996.000 557.240 ;
        RECT 4.000 553.840 995.600 555.240 ;
        RECT 4.000 548.440 996.000 553.840 ;
        RECT 4.400 547.040 996.000 548.440 ;
        RECT 4.000 545.040 996.000 547.040 ;
        RECT 4.000 543.640 995.600 545.040 ;
        RECT 4.000 541.640 996.000 543.640 ;
        RECT 4.400 540.240 996.000 541.640 ;
        RECT 4.000 538.240 996.000 540.240 ;
        RECT 4.000 536.840 995.600 538.240 ;
        RECT 4.000 531.440 996.000 536.840 ;
        RECT 4.400 530.040 996.000 531.440 ;
        RECT 4.000 528.040 996.000 530.040 ;
        RECT 4.000 526.640 995.600 528.040 ;
        RECT 4.000 521.240 996.000 526.640 ;
        RECT 4.400 519.840 996.000 521.240 ;
        RECT 4.000 517.840 996.000 519.840 ;
        RECT 4.000 516.440 995.600 517.840 ;
        RECT 4.000 511.040 996.000 516.440 ;
        RECT 4.400 509.640 996.000 511.040 ;
        RECT 4.000 507.640 996.000 509.640 ;
        RECT 4.000 506.240 995.600 507.640 ;
        RECT 4.000 504.240 996.000 506.240 ;
        RECT 4.400 502.840 996.000 504.240 ;
        RECT 4.000 500.840 996.000 502.840 ;
        RECT 4.000 499.440 995.600 500.840 ;
        RECT 4.000 494.040 996.000 499.440 ;
        RECT 4.400 492.640 996.000 494.040 ;
        RECT 4.000 490.640 996.000 492.640 ;
        RECT 4.000 489.240 995.600 490.640 ;
        RECT 4.000 483.840 996.000 489.240 ;
        RECT 4.400 482.440 996.000 483.840 ;
        RECT 4.000 480.440 996.000 482.440 ;
        RECT 4.000 479.040 995.600 480.440 ;
        RECT 4.000 473.640 996.000 479.040 ;
        RECT 4.400 472.240 996.000 473.640 ;
        RECT 4.000 470.240 996.000 472.240 ;
        RECT 4.000 468.840 995.600 470.240 ;
        RECT 4.000 466.840 996.000 468.840 ;
        RECT 4.400 465.440 996.000 466.840 ;
        RECT 4.000 463.440 996.000 465.440 ;
        RECT 4.000 462.040 995.600 463.440 ;
        RECT 4.000 456.640 996.000 462.040 ;
        RECT 4.400 455.240 996.000 456.640 ;
        RECT 4.000 453.240 996.000 455.240 ;
        RECT 4.000 451.840 995.600 453.240 ;
        RECT 4.000 446.440 996.000 451.840 ;
        RECT 4.400 445.040 996.000 446.440 ;
        RECT 4.000 443.040 996.000 445.040 ;
        RECT 4.000 441.640 995.600 443.040 ;
        RECT 4.000 436.240 996.000 441.640 ;
        RECT 4.400 434.840 995.600 436.240 ;
        RECT 4.000 429.440 996.000 434.840 ;
        RECT 4.400 428.040 996.000 429.440 ;
        RECT 4.000 426.040 996.000 428.040 ;
        RECT 4.000 424.640 995.600 426.040 ;
        RECT 4.000 419.240 996.000 424.640 ;
        RECT 4.400 417.840 996.000 419.240 ;
        RECT 4.000 415.840 996.000 417.840 ;
        RECT 4.000 414.440 995.600 415.840 ;
        RECT 4.000 409.040 996.000 414.440 ;
        RECT 4.400 407.640 996.000 409.040 ;
        RECT 4.000 405.640 996.000 407.640 ;
        RECT 4.000 404.240 995.600 405.640 ;
        RECT 4.000 398.840 996.000 404.240 ;
        RECT 4.400 397.440 995.600 398.840 ;
        RECT 4.000 392.040 996.000 397.440 ;
        RECT 4.400 390.640 996.000 392.040 ;
        RECT 4.000 388.640 996.000 390.640 ;
        RECT 4.000 387.240 995.600 388.640 ;
        RECT 4.000 381.840 996.000 387.240 ;
        RECT 4.400 380.440 996.000 381.840 ;
        RECT 4.000 378.440 996.000 380.440 ;
        RECT 4.000 377.040 995.600 378.440 ;
        RECT 4.000 371.640 996.000 377.040 ;
        RECT 4.400 370.240 996.000 371.640 ;
        RECT 4.000 368.240 996.000 370.240 ;
        RECT 4.000 366.840 995.600 368.240 ;
        RECT 4.000 364.840 996.000 366.840 ;
        RECT 4.400 363.440 996.000 364.840 ;
        RECT 4.000 361.440 996.000 363.440 ;
        RECT 4.000 360.040 995.600 361.440 ;
        RECT 4.000 354.640 996.000 360.040 ;
        RECT 4.400 353.240 996.000 354.640 ;
        RECT 4.000 351.240 996.000 353.240 ;
        RECT 4.000 349.840 995.600 351.240 ;
        RECT 4.000 344.440 996.000 349.840 ;
        RECT 4.400 343.040 996.000 344.440 ;
        RECT 4.000 341.040 996.000 343.040 ;
        RECT 4.000 339.640 995.600 341.040 ;
        RECT 4.000 334.240 996.000 339.640 ;
        RECT 4.400 332.840 996.000 334.240 ;
        RECT 4.000 330.840 996.000 332.840 ;
        RECT 4.000 329.440 995.600 330.840 ;
        RECT 4.000 327.440 996.000 329.440 ;
        RECT 4.400 326.040 996.000 327.440 ;
        RECT 4.000 324.040 996.000 326.040 ;
        RECT 4.000 322.640 995.600 324.040 ;
        RECT 4.000 317.240 996.000 322.640 ;
        RECT 4.400 315.840 996.000 317.240 ;
        RECT 4.000 313.840 996.000 315.840 ;
        RECT 4.000 312.440 995.600 313.840 ;
        RECT 4.000 307.040 996.000 312.440 ;
        RECT 4.400 305.640 996.000 307.040 ;
        RECT 4.000 303.640 996.000 305.640 ;
        RECT 4.000 302.240 995.600 303.640 ;
        RECT 4.000 296.840 996.000 302.240 ;
        RECT 4.400 295.440 996.000 296.840 ;
        RECT 4.000 293.440 996.000 295.440 ;
        RECT 4.000 292.040 995.600 293.440 ;
        RECT 4.000 290.040 996.000 292.040 ;
        RECT 4.400 288.640 996.000 290.040 ;
        RECT 4.000 286.640 996.000 288.640 ;
        RECT 4.000 285.240 995.600 286.640 ;
        RECT 4.000 279.840 996.000 285.240 ;
        RECT 4.400 278.440 996.000 279.840 ;
        RECT 4.000 276.440 996.000 278.440 ;
        RECT 4.000 275.040 995.600 276.440 ;
        RECT 4.000 269.640 996.000 275.040 ;
        RECT 4.400 268.240 996.000 269.640 ;
        RECT 4.000 266.240 996.000 268.240 ;
        RECT 4.000 264.840 995.600 266.240 ;
        RECT 4.000 259.440 996.000 264.840 ;
        RECT 4.400 258.040 996.000 259.440 ;
        RECT 4.000 256.040 996.000 258.040 ;
        RECT 4.000 254.640 995.600 256.040 ;
        RECT 4.000 252.640 996.000 254.640 ;
        RECT 4.400 251.240 996.000 252.640 ;
        RECT 4.000 249.240 996.000 251.240 ;
        RECT 4.000 247.840 995.600 249.240 ;
        RECT 4.000 242.440 996.000 247.840 ;
        RECT 4.400 241.040 996.000 242.440 ;
        RECT 4.000 239.040 996.000 241.040 ;
        RECT 4.000 237.640 995.600 239.040 ;
        RECT 4.000 232.240 996.000 237.640 ;
        RECT 4.400 230.840 996.000 232.240 ;
        RECT 4.000 228.840 996.000 230.840 ;
        RECT 4.000 227.440 995.600 228.840 ;
        RECT 4.000 222.040 996.000 227.440 ;
        RECT 4.400 220.640 996.000 222.040 ;
        RECT 4.000 218.640 996.000 220.640 ;
        RECT 4.000 217.240 995.600 218.640 ;
        RECT 4.000 215.240 996.000 217.240 ;
        RECT 4.400 213.840 996.000 215.240 ;
        RECT 4.000 211.840 996.000 213.840 ;
        RECT 4.000 210.440 995.600 211.840 ;
        RECT 4.000 205.040 996.000 210.440 ;
        RECT 4.400 203.640 996.000 205.040 ;
        RECT 4.000 201.640 996.000 203.640 ;
        RECT 4.000 200.240 995.600 201.640 ;
        RECT 4.000 194.840 996.000 200.240 ;
        RECT 4.400 193.440 996.000 194.840 ;
        RECT 4.000 191.440 996.000 193.440 ;
        RECT 4.000 190.040 995.600 191.440 ;
        RECT 4.000 184.640 996.000 190.040 ;
        RECT 4.400 183.240 996.000 184.640 ;
        RECT 4.000 181.240 996.000 183.240 ;
        RECT 4.000 179.840 995.600 181.240 ;
        RECT 4.000 177.840 996.000 179.840 ;
        RECT 4.400 176.440 996.000 177.840 ;
        RECT 4.000 174.440 996.000 176.440 ;
        RECT 4.000 173.040 995.600 174.440 ;
        RECT 4.000 167.640 996.000 173.040 ;
        RECT 4.400 166.240 996.000 167.640 ;
        RECT 4.000 164.240 996.000 166.240 ;
        RECT 4.000 162.840 995.600 164.240 ;
        RECT 4.000 157.440 996.000 162.840 ;
        RECT 4.400 156.040 996.000 157.440 ;
        RECT 4.000 154.040 996.000 156.040 ;
        RECT 4.000 152.640 995.600 154.040 ;
        RECT 4.000 147.240 996.000 152.640 ;
        RECT 4.400 145.840 996.000 147.240 ;
        RECT 4.000 143.840 996.000 145.840 ;
        RECT 4.000 142.440 995.600 143.840 ;
        RECT 4.000 140.440 996.000 142.440 ;
        RECT 4.400 139.040 996.000 140.440 ;
        RECT 4.000 137.040 996.000 139.040 ;
        RECT 4.000 135.640 995.600 137.040 ;
        RECT 4.000 130.240 996.000 135.640 ;
        RECT 4.400 128.840 996.000 130.240 ;
        RECT 4.000 126.840 996.000 128.840 ;
        RECT 4.000 125.440 995.600 126.840 ;
        RECT 4.000 120.040 996.000 125.440 ;
        RECT 4.400 118.640 996.000 120.040 ;
        RECT 4.000 116.640 996.000 118.640 ;
        RECT 4.000 115.240 995.600 116.640 ;
        RECT 4.000 109.840 996.000 115.240 ;
        RECT 4.400 108.440 996.000 109.840 ;
        RECT 4.000 106.440 996.000 108.440 ;
        RECT 4.000 105.040 995.600 106.440 ;
        RECT 4.000 103.040 996.000 105.040 ;
        RECT 4.400 101.640 996.000 103.040 ;
        RECT 4.000 99.640 996.000 101.640 ;
        RECT 4.000 98.240 995.600 99.640 ;
        RECT 4.000 92.840 996.000 98.240 ;
        RECT 4.400 91.440 996.000 92.840 ;
        RECT 4.000 89.440 996.000 91.440 ;
        RECT 4.000 88.040 995.600 89.440 ;
        RECT 4.000 82.640 996.000 88.040 ;
        RECT 4.400 81.240 996.000 82.640 ;
        RECT 4.000 79.240 996.000 81.240 ;
        RECT 4.000 77.840 995.600 79.240 ;
        RECT 4.000 72.440 996.000 77.840 ;
        RECT 4.400 71.040 996.000 72.440 ;
        RECT 4.000 69.040 996.000 71.040 ;
        RECT 4.000 67.640 995.600 69.040 ;
        RECT 4.000 65.640 996.000 67.640 ;
        RECT 4.400 64.240 996.000 65.640 ;
        RECT 4.000 62.240 996.000 64.240 ;
        RECT 4.000 60.840 995.600 62.240 ;
        RECT 4.000 55.440 996.000 60.840 ;
        RECT 4.400 54.040 996.000 55.440 ;
        RECT 4.000 52.040 996.000 54.040 ;
        RECT 4.000 50.640 995.600 52.040 ;
        RECT 4.000 45.240 996.000 50.640 ;
        RECT 4.400 43.840 996.000 45.240 ;
        RECT 4.000 41.840 996.000 43.840 ;
        RECT 4.000 40.440 995.600 41.840 ;
        RECT 4.000 35.040 996.000 40.440 ;
        RECT 4.400 33.640 995.600 35.040 ;
        RECT 4.000 28.240 996.000 33.640 ;
        RECT 4.400 26.840 996.000 28.240 ;
        RECT 4.000 24.840 996.000 26.840 ;
        RECT 4.000 23.440 995.600 24.840 ;
        RECT 4.000 18.040 996.000 23.440 ;
        RECT 4.400 16.640 996.000 18.040 ;
        RECT 4.000 14.640 996.000 16.640 ;
        RECT 4.000 13.240 995.600 14.640 ;
        RECT 4.000 7.840 996.000 13.240 ;
        RECT 4.400 6.440 996.000 7.840 ;
        RECT 4.000 4.440 996.000 6.440 ;
        RECT 4.000 3.575 995.600 4.440 ;
      LAYER met4 ;
        RECT 402.335 12.415 404.640 985.825 ;
        RECT 407.040 12.415 481.440 985.825 ;
        RECT 483.840 12.415 558.240 985.825 ;
        RECT 560.640 12.415 635.040 985.825 ;
        RECT 637.440 12.415 685.105 985.825 ;
  END
END WB_InterConnect
END LIBRARY

