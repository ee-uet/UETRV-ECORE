magic
tech sky130A
magscale 1 2
timestamp 1647604982
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 14 1980 18860 17456
<< metal2 >>
rect 18 19200 74 20000
rect 1306 19200 1362 20000
rect 1950 19200 2006 20000
rect 2594 19200 2650 20000
rect 3882 19200 3938 20000
rect 4526 19200 4582 20000
rect 5170 19200 5226 20000
rect 6458 19200 6514 20000
rect 7102 19200 7158 20000
rect 7746 19200 7802 20000
rect 9034 19200 9090 20000
rect 9678 19200 9734 20000
rect 10322 19200 10378 20000
rect 11610 19200 11666 20000
rect 12254 19200 12310 20000
rect 12898 19200 12954 20000
rect 14186 19200 14242 20000
rect 14830 19200 14886 20000
rect 15474 19200 15530 20000
rect 16762 19200 16818 20000
rect 17406 19200 17462 20000
rect 18050 19200 18106 20000
rect 19338 19200 19394 20000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
<< obsm2 >>
rect 130 19144 1250 19258
rect 1418 19144 1894 19258
rect 2062 19144 2538 19258
rect 2706 19144 3826 19258
rect 3994 19144 4470 19258
rect 4638 19144 5114 19258
rect 5282 19144 6402 19258
rect 6570 19144 7046 19258
rect 7214 19144 7690 19258
rect 7858 19144 8978 19258
rect 9146 19144 9622 19258
rect 9790 19144 10266 19258
rect 10434 19144 11554 19258
rect 11722 19144 12198 19258
rect 12366 19144 12842 19258
rect 13010 19144 14130 19258
rect 14298 19144 14774 19258
rect 14942 19144 15418 19258
rect 15586 19144 16706 19258
rect 16874 19144 17350 19258
rect 17518 19144 17994 19258
rect 18162 19144 18748 19258
rect 20 856 18748 19144
rect 130 711 606 856
rect 774 711 1250 856
rect 1418 711 2538 856
rect 2706 711 3182 856
rect 3350 711 3826 856
rect 3994 711 5114 856
rect 5282 711 5758 856
rect 5926 711 6402 856
rect 6570 711 7690 856
rect 7858 711 8334 856
rect 8502 711 8978 856
rect 9146 711 10266 856
rect 10434 711 10910 856
rect 11078 711 11554 856
rect 11722 711 12842 856
rect 13010 711 13486 856
rect 13654 711 14130 856
rect 14298 711 15418 856
rect 15586 711 16062 856
rect 16230 711 16706 856
rect 16874 711 17994 856
rect 18162 711 18638 856
<< metal3 >>
rect 0 19728 800 19848
rect 19200 19728 20000 19848
rect 0 19048 800 19168
rect 19200 18368 20000 18488
rect 0 17688 800 17808
rect 19200 17688 20000 17808
rect 0 17008 800 17128
rect 19200 17008 20000 17128
rect 0 16328 800 16448
rect 19200 15648 20000 15768
rect 0 14968 800 15088
rect 19200 14968 20000 15088
rect 0 14288 800 14408
rect 19200 14288 20000 14408
rect 0 13608 800 13728
rect 19200 12928 20000 13048
rect 0 12248 800 12368
rect 19200 12248 20000 12368
rect 0 11568 800 11688
rect 19200 11568 20000 11688
rect 0 10888 800 11008
rect 19200 10208 20000 10328
rect 0 9528 800 9648
rect 19200 9528 20000 9648
rect 0 8848 800 8968
rect 19200 8848 20000 8968
rect 0 8168 800 8288
rect 19200 7488 20000 7608
rect 0 6808 800 6928
rect 19200 6808 20000 6928
rect 0 6128 800 6248
rect 19200 6128 20000 6248
rect 0 5448 800 5568
rect 19200 4768 20000 4888
rect 0 4088 800 4208
rect 19200 4088 20000 4208
rect 0 3408 800 3528
rect 19200 3408 20000 3528
rect 0 2728 800 2848
rect 19200 2048 20000 2168
rect 0 1368 800 1488
rect 19200 1368 20000 1488
rect 0 688 800 808
rect 19200 688 20000 808
<< obsm3 >>
rect 880 18968 19200 19141
rect 800 18568 19200 18968
rect 800 18288 19120 18568
rect 800 17888 19200 18288
rect 880 17608 19120 17888
rect 800 17208 19200 17608
rect 880 16928 19120 17208
rect 800 16528 19200 16928
rect 880 16248 19200 16528
rect 800 15848 19200 16248
rect 800 15568 19120 15848
rect 800 15168 19200 15568
rect 880 14888 19120 15168
rect 800 14488 19200 14888
rect 880 14208 19120 14488
rect 800 13808 19200 14208
rect 880 13528 19200 13808
rect 800 13128 19200 13528
rect 800 12848 19120 13128
rect 800 12448 19200 12848
rect 880 12168 19120 12448
rect 800 11768 19200 12168
rect 880 11488 19120 11768
rect 800 11088 19200 11488
rect 880 10808 19200 11088
rect 800 10408 19200 10808
rect 800 10128 19120 10408
rect 800 9728 19200 10128
rect 880 9448 19120 9728
rect 800 9048 19200 9448
rect 880 8768 19120 9048
rect 800 8368 19200 8768
rect 880 8088 19200 8368
rect 800 7688 19200 8088
rect 800 7408 19120 7688
rect 800 7008 19200 7408
rect 880 6728 19120 7008
rect 800 6328 19200 6728
rect 880 6048 19120 6328
rect 800 5648 19200 6048
rect 880 5368 19200 5648
rect 800 4968 19200 5368
rect 800 4688 19120 4968
rect 800 4288 19200 4688
rect 880 4008 19120 4288
rect 800 3608 19200 4008
rect 880 3328 19120 3608
rect 800 2928 19200 3328
rect 880 2648 19200 2928
rect 800 2248 19200 2648
rect 800 1968 19120 2248
rect 800 1568 19200 1968
rect 880 1288 19120 1568
rect 800 888 19200 1288
rect 880 715 19120 888
<< metal4 >>
rect 3910 2128 4230 17456
rect 6874 2128 7194 17456
rect 9840 2128 10160 17456
rect 12805 2128 13125 17456
rect 15771 2128 16091 17456
<< obsm4 >>
rect 4310 2128 6794 17456
rect 7274 2128 9760 17456
rect 10240 2128 12725 17456
rect 13205 2128 15691 17456
<< labels >>
rlabel metal3 s 0 1368 800 1488 6 clock
port 1 nsew signal input
rlabel metal2 s 18050 19200 18106 20000 6 io_spi_clk
port 2 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 io_spi_cs
port 3 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 io_spi_intr
port 4 nsew signal output
rlabel metal2 s 7102 19200 7158 20000 6 io_spi_miso
port 5 nsew signal input
rlabel metal2 s 7746 19200 7802 20000 6 io_spi_mosi
port 6 nsew signal output
rlabel metal2 s 9034 19200 9090 20000 6 io_spi_select
port 7 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 io_wbs_ack_o
port 8 nsew signal output
rlabel metal3 s 19200 4088 20000 4208 6 io_wbs_data_o[0]
port 9 nsew signal output
rlabel metal2 s 17406 19200 17462 20000 6 io_wbs_data_o[10]
port 10 nsew signal output
rlabel metal2 s 10322 19200 10378 20000 6 io_wbs_data_o[11]
port 11 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 io_wbs_data_o[12]
port 12 nsew signal output
rlabel metal3 s 19200 6128 20000 6248 6 io_wbs_data_o[13]
port 13 nsew signal output
rlabel metal3 s 19200 8848 20000 8968 6 io_wbs_data_o[14]
port 14 nsew signal output
rlabel metal3 s 19200 17688 20000 17808 6 io_wbs_data_o[15]
port 15 nsew signal output
rlabel metal3 s 19200 15648 20000 15768 6 io_wbs_data_o[16]
port 16 nsew signal output
rlabel metal3 s 19200 2048 20000 2168 6 io_wbs_data_o[17]
port 17 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 io_wbs_data_o[18]
port 18 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 io_wbs_data_o[19]
port 19 nsew signal output
rlabel metal3 s 19200 12928 20000 13048 6 io_wbs_data_o[1]
port 20 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 io_wbs_data_o[20]
port 21 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 io_wbs_data_o[21]
port 22 nsew signal output
rlabel metal3 s 19200 14288 20000 14408 6 io_wbs_data_o[22]
port 23 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 io_wbs_data_o[23]
port 24 nsew signal output
rlabel metal2 s 12254 19200 12310 20000 6 io_wbs_data_o[24]
port 25 nsew signal output
rlabel metal2 s 18 19200 74 20000 6 io_wbs_data_o[25]
port 26 nsew signal output
rlabel metal3 s 19200 14968 20000 15088 6 io_wbs_data_o[26]
port 27 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 io_wbs_data_o[27]
port 28 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_wbs_data_o[28]
port 29 nsew signal output
rlabel metal3 s 0 688 800 808 6 io_wbs_data_o[29]
port 30 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 io_wbs_data_o[2]
port 31 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 io_wbs_data_o[30]
port 32 nsew signal output
rlabel metal2 s 12898 19200 12954 20000 6 io_wbs_data_o[31]
port 33 nsew signal output
rlabel metal2 s 14186 19200 14242 20000 6 io_wbs_data_o[3]
port 34 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 io_wbs_data_o[4]
port 35 nsew signal output
rlabel metal2 s 9678 19200 9734 20000 6 io_wbs_data_o[5]
port 36 nsew signal output
rlabel metal3 s 19200 17008 20000 17128 6 io_wbs_data_o[6]
port 37 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 io_wbs_data_o[7]
port 38 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_wbs_data_o[8]
port 39 nsew signal output
rlabel metal3 s 19200 688 20000 808 6 io_wbs_data_o[9]
port 40 nsew signal output
rlabel metal3 s 19200 7488 20000 7608 6 io_wbs_m2s_addr[0]
port 41 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 io_wbs_m2s_addr[10]
port 42 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 io_wbs_m2s_addr[11]
port 43 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 io_wbs_m2s_addr[12]
port 44 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 io_wbs_m2s_addr[13]
port 45 nsew signal input
rlabel metal3 s 19200 18368 20000 18488 6 io_wbs_m2s_addr[14]
port 46 nsew signal input
rlabel metal2 s 3882 19200 3938 20000 6 io_wbs_m2s_addr[15]
port 47 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 io_wbs_m2s_addr[1]
port 48 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 io_wbs_m2s_addr[2]
port 49 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_wbs_m2s_addr[3]
port 50 nsew signal input
rlabel metal3 s 19200 6808 20000 6928 6 io_wbs_m2s_addr[4]
port 51 nsew signal input
rlabel metal3 s 19200 3408 20000 3528 6 io_wbs_m2s_addr[5]
port 52 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 io_wbs_m2s_addr[6]
port 53 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_wbs_m2s_addr[7]
port 54 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_wbs_m2s_addr[8]
port 55 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 io_wbs_m2s_addr[9]
port 56 nsew signal input
rlabel metal3 s 19200 4768 20000 4888 6 io_wbs_m2s_data[0]
port 57 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 io_wbs_m2s_data[10]
port 58 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 io_wbs_m2s_data[11]
port 59 nsew signal input
rlabel metal3 s 19200 12248 20000 12368 6 io_wbs_m2s_data[12]
port 60 nsew signal input
rlabel metal2 s 5170 19200 5226 20000 6 io_wbs_m2s_data[13]
port 61 nsew signal input
rlabel metal2 s 2594 19200 2650 20000 6 io_wbs_m2s_data[14]
port 62 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 io_wbs_m2s_data[15]
port 63 nsew signal input
rlabel metal2 s 18 0 74 800 6 io_wbs_m2s_data[16]
port 64 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 io_wbs_m2s_data[17]
port 65 nsew signal input
rlabel metal2 s 6458 19200 6514 20000 6 io_wbs_m2s_data[18]
port 66 nsew signal input
rlabel metal2 s 11610 19200 11666 20000 6 io_wbs_m2s_data[19]
port 67 nsew signal input
rlabel metal2 s 16762 19200 16818 20000 6 io_wbs_m2s_data[1]
port 68 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 io_wbs_m2s_data[20]
port 69 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 io_wbs_m2s_data[21]
port 70 nsew signal input
rlabel metal2 s 662 0 718 800 6 io_wbs_m2s_data[22]
port 71 nsew signal input
rlabel metal2 s 19338 19200 19394 20000 6 io_wbs_m2s_data[23]
port 72 nsew signal input
rlabel metal2 s 14830 19200 14886 20000 6 io_wbs_m2s_data[24]
port 73 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 io_wbs_m2s_data[25]
port 74 nsew signal input
rlabel metal3 s 19200 19728 20000 19848 6 io_wbs_m2s_data[26]
port 75 nsew signal input
rlabel metal3 s 19200 1368 20000 1488 6 io_wbs_m2s_data[27]
port 76 nsew signal input
rlabel metal2 s 1950 19200 2006 20000 6 io_wbs_m2s_data[28]
port 77 nsew signal input
rlabel metal3 s 19200 10208 20000 10328 6 io_wbs_m2s_data[29]
port 78 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 io_wbs_m2s_data[2]
port 79 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 io_wbs_m2s_data[30]
port 80 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 io_wbs_m2s_data[31]
port 81 nsew signal input
rlabel metal3 s 19200 11568 20000 11688 6 io_wbs_m2s_data[3]
port 82 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 io_wbs_m2s_data[4]
port 83 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_wbs_m2s_data[5]
port 84 nsew signal input
rlabel metal2 s 15474 19200 15530 20000 6 io_wbs_m2s_data[6]
port 85 nsew signal input
rlabel metal2 s 1306 19200 1362 20000 6 io_wbs_m2s_data[7]
port 86 nsew signal input
rlabel metal2 s 4526 19200 4582 20000 6 io_wbs_m2s_data[8]
port 87 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 io_wbs_m2s_data[9]
port 88 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 io_wbs_m2s_stb
port 89 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 io_wbs_m2s_we
port 90 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 reset
port 91 nsew signal input
rlabel metal4 s 3910 2128 4230 17456 6 vccd1
port 92 nsew power input
rlabel metal4 s 9840 2128 10160 17456 6 vccd1
port 92 nsew power input
rlabel metal4 s 15771 2128 16091 17456 6 vccd1
port 92 nsew power input
rlabel metal4 s 6874 2128 7194 17456 6 vssd1
port 93 nsew ground input
rlabel metal4 s 12805 2128 13125 17456 6 vssd1
port 93 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1421962
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/SPI/runs/SPI/results/finishing/SPI.magic.gds
string GDS_START 332394
<< end >>

