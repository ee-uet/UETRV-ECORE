magic
tech sky130A
magscale 1 2
timestamp 1649148650
<< metal1 >>
rect 242894 536800 242900 536852
rect 242952 536840 242958 536852
rect 396626 536840 396632 536852
rect 242952 536812 396632 536840
rect 242952 536800 242958 536812
rect 396626 536800 396632 536812
rect 396684 536800 396690 536852
rect 237374 535440 237380 535492
rect 237432 535480 237438 535492
rect 396626 535480 396632 535492
rect 237432 535452 396632 535480
rect 237432 535440 237438 535452
rect 396626 535440 396632 535452
rect 396684 535440 396690 535492
rect 231854 532788 231860 532840
rect 231912 532828 231918 532840
rect 396718 532828 396724 532840
rect 231912 532800 396724 532828
rect 231912 532788 231918 532800
rect 396718 532788 396724 532800
rect 396776 532788 396782 532840
rect 226334 532720 226340 532772
rect 226392 532760 226398 532772
rect 396626 532760 396632 532772
rect 226392 532732 396632 532760
rect 226392 532720 226398 532732
rect 396626 532720 396632 532732
rect 396684 532720 396690 532772
rect 222194 530000 222200 530052
rect 222252 530040 222258 530052
rect 396718 530040 396724 530052
rect 222252 530012 396724 530040
rect 222252 530000 222258 530012
rect 396718 530000 396724 530012
rect 396776 530000 396782 530052
rect 213914 529932 213920 529984
rect 213972 529972 213978 529984
rect 396626 529972 396632 529984
rect 213972 529944 396632 529972
rect 213972 529932 213978 529944
rect 396626 529932 396632 529944
rect 396684 529932 396690 529984
rect 207014 527144 207020 527196
rect 207072 527184 207078 527196
rect 396626 527184 396632 527196
rect 207072 527156 396632 527184
rect 207072 527144 207078 527156
rect 396626 527144 396632 527156
rect 396684 527144 396690 527196
rect 191834 509260 191840 509312
rect 191892 509300 191898 509312
rect 396350 509300 396356 509312
rect 191892 509272 396356 509300
rect 191892 509260 191898 509272
rect 396350 509260 396356 509272
rect 396408 509260 396414 509312
rect 190454 507832 190460 507884
rect 190512 507872 190518 507884
rect 396626 507872 396632 507884
rect 190512 507844 396632 507872
rect 190512 507832 190518 507844
rect 396626 507832 396632 507844
rect 396684 507832 396690 507884
rect 48130 498856 48136 498908
rect 48188 498896 48194 498908
rect 177298 498896 177304 498908
rect 48188 498868 177304 498896
rect 48188 498856 48194 498868
rect 177298 498856 177304 498868
rect 177356 498856 177362 498908
rect 49418 498788 49424 498840
rect 49476 498828 49482 498840
rect 338114 498828 338120 498840
rect 49476 498800 338120 498828
rect 49476 498788 49482 498800
rect 338114 498788 338120 498800
rect 338172 498788 338178 498840
rect 457438 498040 457444 498092
rect 457496 498080 457502 498092
rect 462314 498080 462320 498092
rect 457496 498052 462320 498080
rect 457496 498040 457502 498052
rect 462314 498040 462320 498052
rect 462372 498040 462378 498092
rect 49326 497768 49332 497820
rect 49384 497808 49390 497820
rect 53834 497808 53840 497820
rect 49384 497780 53840 497808
rect 49384 497768 49390 497780
rect 53834 497768 53840 497780
rect 53892 497768 53898 497820
rect 116854 497428 116860 497480
rect 116912 497468 116918 497480
rect 133138 497468 133144 497480
rect 116912 497440 133144 497468
rect 116912 497428 116918 497440
rect 133138 497428 133144 497440
rect 133196 497428 133202 497480
rect 113542 497360 113548 497412
rect 113600 497400 113606 497412
rect 131850 497400 131856 497412
rect 113600 497372 131856 497400
rect 113600 497360 113606 497372
rect 131850 497360 131856 497372
rect 131908 497360 131914 497412
rect 92290 497292 92296 497344
rect 92348 497332 92354 497344
rect 131758 497332 131764 497344
rect 92348 497304 131764 497332
rect 92348 497292 92354 497304
rect 131758 497292 131764 497304
rect 131816 497292 131822 497344
rect 89530 497224 89536 497276
rect 89588 497264 89594 497276
rect 130470 497264 130476 497276
rect 89588 497236 130476 497264
rect 89588 497224 89594 497236
rect 130470 497224 130476 497236
rect 130528 497224 130534 497276
rect 85942 497156 85948 497208
rect 86000 497196 86006 497208
rect 130378 497196 130384 497208
rect 86000 497168 130384 497196
rect 86000 497156 86006 497168
rect 130378 497156 130384 497168
rect 130436 497156 130442 497208
rect 118602 497088 118608 497140
rect 118660 497128 118666 497140
rect 189810 497128 189816 497140
rect 118660 497100 189816 497128
rect 118660 497088 118666 497100
rect 189810 497088 189816 497100
rect 189868 497088 189874 497140
rect 86494 497020 86500 497072
rect 86552 497060 86558 497072
rect 189718 497060 189724 497072
rect 86552 497032 189724 497060
rect 86552 497020 86558 497032
rect 189718 497020 189724 497032
rect 189776 497020 189782 497072
rect 410518 497020 410524 497072
rect 410576 497060 410582 497072
rect 432138 497060 432144 497072
rect 410576 497032 432144 497060
rect 410576 497020 410582 497032
rect 432138 497020 432144 497032
rect 432196 497020 432202 497072
rect 81250 496952 81256 497004
rect 81308 496992 81314 497004
rect 185578 496992 185584 497004
rect 81308 496964 185584 496992
rect 81308 496952 81314 496964
rect 185578 496952 185584 496964
rect 185636 496952 185642 497004
rect 432598 496952 432604 497004
rect 432656 496992 432662 497004
rect 456794 496992 456800 497004
rect 432656 496964 456800 496992
rect 432656 496952 432662 496964
rect 456794 496952 456800 496964
rect 456852 496952 456858 497004
rect 79870 496884 79876 496936
rect 79928 496924 79934 496936
rect 188338 496924 188344 496936
rect 79928 496896 188344 496924
rect 79928 496884 79934 496896
rect 188338 496884 188344 496896
rect 188396 496884 188402 496936
rect 284938 496884 284944 496936
rect 284996 496924 285002 496936
rect 426434 496924 426440 496936
rect 284996 496896 426440 496924
rect 284996 496884 285002 496896
rect 426434 496884 426440 496896
rect 426492 496884 426498 496936
rect 427078 496884 427084 496936
rect 427136 496924 427142 496936
rect 430574 496924 430580 496936
rect 427136 496896 430580 496924
rect 427136 496884 427142 496896
rect 430574 496884 430580 496896
rect 430632 496884 430638 496936
rect 494698 496884 494704 496936
rect 494756 496924 494762 496936
rect 498194 496924 498200 496936
rect 494756 496896 498200 496924
rect 494756 496884 494762 496896
rect 498194 496884 498200 496896
rect 498252 496884 498258 496936
rect 73338 496816 73344 496868
rect 73396 496856 73402 496868
rect 75178 496856 75184 496868
rect 73396 496828 75184 496856
rect 73396 496816 73402 496828
rect 75178 496816 75184 496828
rect 75236 496816 75242 496868
rect 78306 496816 78312 496868
rect 78364 496856 78370 496868
rect 79318 496856 79324 496868
rect 78364 496828 79324 496856
rect 78364 496816 78370 496828
rect 79318 496816 79324 496828
rect 79376 496816 79382 496868
rect 103422 496816 103428 496868
rect 103480 496856 103486 496868
rect 150894 496856 150900 496868
rect 103480 496828 150900 496856
rect 103480 496816 103486 496828
rect 150894 496816 150900 496828
rect 150952 496816 150958 496868
rect 150986 496816 150992 496868
rect 151044 496856 151050 496868
rect 359458 496856 359464 496868
rect 151044 496828 359464 496856
rect 151044 496816 151050 496828
rect 359458 496816 359464 496828
rect 359516 496816 359522 496868
rect 424318 496816 424324 496868
rect 424376 496856 424382 496868
rect 426526 496856 426532 496868
rect 424376 496828 426532 496856
rect 424376 496816 424382 496828
rect 426526 496816 426532 496828
rect 426584 496816 426590 496868
rect 428458 496816 428464 496868
rect 428516 496856 428522 496868
rect 433334 496856 433340 496868
rect 428516 496828 433340 496856
rect 428516 496816 428522 496828
rect 433334 496816 433340 496828
rect 433392 496816 433398 496868
rect 479518 496816 479524 496868
rect 479576 496856 479582 496868
rect 495434 496856 495440 496868
rect 479576 496828 495440 496856
rect 479576 496816 479582 496828
rect 495434 496816 495440 496828
rect 495492 496816 495498 496868
rect 497458 496816 497464 496868
rect 497516 496856 497522 496868
rect 505094 496856 505100 496868
rect 497516 496828 505100 496856
rect 497516 496816 497522 496828
rect 505094 496816 505100 496828
rect 505152 496816 505158 496868
rect 96338 496136 96344 496188
rect 96396 496176 96402 496188
rect 184198 496176 184204 496188
rect 96396 496148 184204 496176
rect 96396 496136 96402 496148
rect 184198 496136 184204 496148
rect 184256 496136 184262 496188
rect 47946 496068 47952 496120
rect 48004 496108 48010 496120
rect 163498 496108 163504 496120
rect 48004 496080 163504 496108
rect 48004 496068 48010 496080
rect 163498 496068 163504 496080
rect 163556 496068 163562 496120
rect 193214 496068 193220 496120
rect 193272 496108 193278 496120
rect 415394 496108 415400 496120
rect 193272 496080 415400 496108
rect 193272 496068 193278 496080
rect 415394 496068 415400 496080
rect 415452 496068 415458 496120
rect 255314 494776 255320 494828
rect 255372 494816 255378 494828
rect 455782 494816 455788 494828
rect 255372 494788 455788 494816
rect 255372 494776 255378 494788
rect 455782 494776 455788 494788
rect 455840 494776 455846 494828
rect 49510 494708 49516 494760
rect 49568 494748 49574 494760
rect 340874 494748 340880 494760
rect 49568 494720 340880 494748
rect 49568 494708 49574 494720
rect 340874 494708 340880 494720
rect 340932 494708 340938 494760
rect 106090 493348 106096 493400
rect 106148 493388 106154 493400
rect 177390 493388 177396 493400
rect 106148 493360 177396 493388
rect 106148 493348 106154 493360
rect 177390 493348 177396 493360
rect 177448 493348 177454 493400
rect 47854 493280 47860 493332
rect 47912 493320 47918 493332
rect 175918 493320 175924 493332
rect 47912 493292 175924 493320
rect 47912 493280 47918 493292
rect 175918 493280 175924 493292
rect 175976 493280 175982 493332
rect 209774 493280 209780 493332
rect 209832 493320 209838 493332
rect 433426 493320 433432 493332
rect 209832 493292 433432 493320
rect 209832 493280 209838 493292
rect 433426 493280 433432 493292
rect 433484 493280 433490 493332
rect 89162 491920 89168 491972
rect 89220 491960 89226 491972
rect 166258 491960 166264 491972
rect 89220 491932 166264 491960
rect 89220 491920 89226 491932
rect 166258 491920 166264 491932
rect 166316 491920 166322 491972
rect 195974 491920 195980 491972
rect 196032 491960 196038 491972
rect 427906 491960 427912 491972
rect 196032 491932 427912 491960
rect 196032 491920 196038 491932
rect 427906 491920 427912 491932
rect 427964 491920 427970 491972
rect 91186 490560 91192 490612
rect 91244 490600 91250 490612
rect 170398 490600 170404 490612
rect 91244 490572 170404 490600
rect 91244 490560 91250 490572
rect 170398 490560 170404 490572
rect 170456 490560 170462 490612
rect 204898 490560 204904 490612
rect 204956 490600 204962 490612
rect 419626 490600 419632 490612
rect 204956 490572 419632 490600
rect 204956 490560 204962 490572
rect 419626 490560 419632 490572
rect 419684 490560 419690 490612
rect 88150 489132 88156 489184
rect 88208 489172 88214 489184
rect 162118 489172 162124 489184
rect 88208 489144 162124 489172
rect 88208 489132 88214 489144
rect 162118 489132 162124 489144
rect 162176 489132 162182 489184
rect 216674 489132 216680 489184
rect 216732 489172 216738 489184
rect 434806 489172 434812 489184
rect 216732 489144 434812 489172
rect 216732 489132 216738 489144
rect 434806 489132 434812 489144
rect 434864 489132 434870 489184
rect 74350 487772 74356 487824
rect 74408 487812 74414 487824
rect 155218 487812 155224 487824
rect 74408 487784 155224 487812
rect 74408 487772 74414 487784
rect 155218 487772 155224 487784
rect 155276 487772 155282 487824
rect 211798 487772 211804 487824
rect 211856 487812 211862 487824
rect 419534 487812 419540 487824
rect 211856 487784 419540 487812
rect 211856 487772 211862 487784
rect 419534 487772 419540 487784
rect 419592 487772 419598 487824
rect 101950 486480 101956 486532
rect 102008 486520 102014 486532
rect 176010 486520 176016 486532
rect 102008 486492 176016 486520
rect 102008 486480 102014 486492
rect 176010 486480 176016 486492
rect 176068 486480 176074 486532
rect 198734 486480 198740 486532
rect 198792 486520 198798 486532
rect 422294 486520 422300 486532
rect 198792 486492 422300 486520
rect 198792 486480 198798 486492
rect 422294 486480 422300 486492
rect 422352 486480 422358 486532
rect 48038 486412 48044 486464
rect 48096 486452 48102 486464
rect 409874 486452 409880 486464
rect 48096 486424 409880 486452
rect 48096 486412 48102 486424
rect 409874 486412 409880 486424
rect 409932 486412 409938 486464
rect 252554 485120 252560 485172
rect 252612 485160 252618 485172
rect 433518 485160 433524 485172
rect 252612 485132 433524 485160
rect 252612 485120 252618 485132
rect 433518 485120 433524 485132
rect 433576 485120 433582 485172
rect 96430 485052 96436 485104
rect 96488 485092 96494 485104
rect 383654 485092 383660 485104
rect 96488 485064 383660 485092
rect 96488 485052 96494 485064
rect 383654 485052 383660 485064
rect 383712 485052 383718 485104
rect 263594 483624 263600 483676
rect 263652 483664 263658 483676
rect 437566 483664 437572 483676
rect 263652 483636 437572 483664
rect 263652 483624 263658 483636
rect 437566 483624 437572 483636
rect 437624 483624 437630 483676
rect 281534 482332 281540 482384
rect 281592 482372 281598 482384
rect 443086 482372 443092 482384
rect 281592 482344 443092 482372
rect 281592 482332 281598 482344
rect 443086 482332 443092 482344
rect 443144 482332 443150 482384
rect 75178 482264 75184 482316
rect 75236 482304 75242 482316
rect 331214 482304 331220 482316
rect 75236 482276 331220 482304
rect 75236 482264 75242 482276
rect 331214 482264 331220 482276
rect 331272 482264 331278 482316
rect 104710 480904 104716 480956
rect 104768 480944 104774 480956
rect 182818 480944 182824 480956
rect 104768 480916 182824 480944
rect 104768 480904 104774 480916
rect 182818 480904 182824 480916
rect 182876 480904 182882 480956
rect 205634 480904 205640 480956
rect 205692 480944 205698 480956
rect 423674 480944 423680 480956
rect 205692 480916 423680 480944
rect 205692 480904 205698 480916
rect 423674 480904 423680 480916
rect 423732 480904 423738 480956
rect 302234 479544 302240 479596
rect 302292 479584 302298 479596
rect 449986 479584 449992 479596
rect 302292 479556 449992 479584
rect 302292 479544 302298 479556
rect 449986 479544 449992 479556
rect 450044 479544 450050 479596
rect 133782 479476 133788 479528
rect 133840 479516 133846 479528
rect 389174 479516 389180 479528
rect 133840 479488 389180 479516
rect 133840 479476 133846 479488
rect 389174 479476 389180 479488
rect 389232 479476 389238 479528
rect 110322 478116 110328 478168
rect 110380 478156 110386 478168
rect 181438 478156 181444 478168
rect 110380 478128 181444 478156
rect 110380 478116 110386 478128
rect 181438 478116 181444 478128
rect 181496 478116 181502 478168
rect 273254 478116 273260 478168
rect 273312 478156 273318 478168
rect 441706 478156 441712 478168
rect 273312 478128 441712 478156
rect 273312 478116 273318 478128
rect 441706 478116 441712 478128
rect 441764 478116 441770 478168
rect 288434 476824 288440 476876
rect 288492 476864 288498 476876
rect 445846 476864 445852 476876
rect 288492 476836 445852 476864
rect 288492 476824 288498 476836
rect 445846 476824 445852 476836
rect 445904 476824 445910 476876
rect 108850 476756 108856 476808
rect 108908 476796 108914 476808
rect 407758 476796 407764 476808
rect 108908 476768 407764 476796
rect 108908 476756 108914 476768
rect 407758 476756 407764 476768
rect 407816 476756 407822 476808
rect 298094 475328 298100 475380
rect 298152 475368 298158 475380
rect 448606 475368 448612 475380
rect 298152 475340 448612 475368
rect 298152 475328 298158 475340
rect 448606 475328 448612 475340
rect 448664 475328 448670 475380
rect 304994 474036 305000 474088
rect 305052 474076 305058 474088
rect 451274 474076 451280 474088
rect 305052 474048 451280 474076
rect 305052 474036 305058 474048
rect 451274 474036 451280 474048
rect 451332 474036 451338 474088
rect 77202 473968 77208 474020
rect 77260 474008 77266 474020
rect 342898 474008 342904 474020
rect 77260 473980 342904 474008
rect 77260 473968 77266 473980
rect 342898 473968 342904 473980
rect 342956 473968 342962 474020
rect 291194 472676 291200 472728
rect 291252 472716 291258 472728
rect 447226 472716 447232 472728
rect 291252 472688 447232 472716
rect 291252 472676 291258 472688
rect 447226 472676 447232 472688
rect 447284 472676 447290 472728
rect 81250 472608 81256 472660
rect 81308 472648 81314 472660
rect 356054 472648 356060 472660
rect 81308 472620 356060 472648
rect 81308 472608 81314 472620
rect 356054 472608 356060 472620
rect 356112 472608 356118 472660
rect 212534 471248 212540 471300
rect 212592 471288 212598 471300
rect 425054 471288 425060 471300
rect 212592 471260 425060 471288
rect 212592 471248 212598 471260
rect 425054 471248 425060 471260
rect 425112 471248 425118 471300
rect 309134 469820 309140 469872
rect 309192 469860 309198 469872
rect 452746 469860 452752 469872
rect 309192 469832 452752 469860
rect 309192 469820 309198 469832
rect 452746 469820 452752 469832
rect 452804 469820 452810 469872
rect 230474 467100 230480 467152
rect 230532 467140 230538 467152
rect 427814 467140 427820 467152
rect 230532 467112 427820 467140
rect 230532 467100 230538 467112
rect 427814 467100 427820 467112
rect 427872 467100 427878 467152
rect 316034 465672 316040 465724
rect 316092 465712 316098 465724
rect 454678 465712 454684 465724
rect 316092 465684 454684 465712
rect 316092 465672 316098 465684
rect 454678 465672 454684 465684
rect 454736 465672 454742 465724
rect 245654 457444 245660 457496
rect 245712 457484 245718 457496
rect 410518 457484 410524 457496
rect 245712 457456 410524 457484
rect 245712 457444 245718 457456
rect 410518 457444 410524 457456
rect 410576 457444 410582 457496
rect 235994 454656 236000 454708
rect 236052 454696 236058 454708
rect 429194 454696 429200 454708
rect 236052 454668 429200 454696
rect 236052 454656 236058 454668
rect 429194 454656 429200 454668
rect 429252 454656 429258 454708
rect 224954 453296 224960 453348
rect 225012 453336 225018 453348
rect 424318 453336 424324 453348
rect 225012 453308 424324 453336
rect 225012 453296 225018 453308
rect 424318 453296 424324 453308
rect 424376 453296 424382 453348
rect 325694 451936 325700 451988
rect 325752 451976 325758 451988
rect 458266 451976 458272 451988
rect 325752 451948 458272 451976
rect 325752 451936 325758 451948
rect 458266 451936 458272 451948
rect 458324 451936 458330 451988
rect 157242 451868 157248 451920
rect 157300 451908 157306 451920
rect 410702 451908 410708 451920
rect 157300 451880 410708 451908
rect 157300 451868 157306 451880
rect 410702 451868 410708 451880
rect 410760 451868 410766 451920
rect 219434 450576 219440 450628
rect 219492 450616 219498 450628
rect 284938 450616 284944 450628
rect 219492 450588 284944 450616
rect 219492 450576 219498 450588
rect 284938 450576 284944 450588
rect 284996 450576 285002 450628
rect 322934 450576 322940 450628
rect 322992 450616 322998 450628
rect 432598 450616 432604 450628
rect 322992 450588 432604 450616
rect 322992 450576 322998 450588
rect 432598 450576 432604 450588
rect 432656 450576 432662 450628
rect 154482 450508 154488 450560
rect 154540 450548 154546 450560
rect 409230 450548 409236 450560
rect 154540 450520 409236 450548
rect 154540 450508 154546 450520
rect 409230 450508 409236 450520
rect 409288 450508 409294 450560
rect 318794 449216 318800 449268
rect 318852 449256 318858 449268
rect 456886 449256 456892 449268
rect 318852 449228 456892 449256
rect 318852 449216 318858 449228
rect 456886 449216 456892 449228
rect 456944 449216 456950 449268
rect 103330 449148 103336 449200
rect 103388 449188 103394 449200
rect 410610 449188 410616 449200
rect 103388 449160 410616 449188
rect 103388 449148 103394 449160
rect 410610 449148 410616 449160
rect 410668 449148 410674 449200
rect 311894 447856 311900 447908
rect 311952 447896 311958 447908
rect 454034 447896 454040 447908
rect 311952 447868 454040 447896
rect 311952 447856 311958 447868
rect 454034 447856 454040 447868
rect 454092 447856 454098 447908
rect 102042 447788 102048 447840
rect 102100 447828 102106 447840
rect 411990 447828 411996 447840
rect 102100 447800 411996 447828
rect 102100 447788 102106 447800
rect 411990 447788 411996 447800
rect 412048 447788 412054 447840
rect 295334 446428 295340 446480
rect 295392 446468 295398 446480
rect 448514 446468 448520 446480
rect 295392 446440 448520 446468
rect 295392 446428 295398 446440
rect 448514 446428 448520 446440
rect 448572 446428 448578 446480
rect 100662 446360 100668 446412
rect 100720 446400 100726 446412
rect 410426 446400 410432 446412
rect 100720 446372 410432 446400
rect 100720 446360 100726 446372
rect 410426 446360 410432 446372
rect 410484 446360 410490 446412
rect 324314 445068 324320 445120
rect 324372 445108 324378 445120
rect 497458 445108 497464 445120
rect 324372 445080 497464 445108
rect 324372 445068 324378 445080
rect 497458 445068 497464 445080
rect 497516 445068 497522 445120
rect 93670 445000 93676 445052
rect 93728 445040 93734 445052
rect 378134 445040 378140 445052
rect 93728 445012 378140 445040
rect 93728 445000 93734 445012
rect 378134 445000 378140 445012
rect 378192 445000 378198 445052
rect 321554 443708 321560 443760
rect 321612 443748 321618 443760
rect 502334 443748 502340 443760
rect 321612 443720 502340 443748
rect 321612 443708 321618 443720
rect 502334 443708 502340 443720
rect 502392 443708 502398 443760
rect 99190 443640 99196 443692
rect 99248 443680 99254 443692
rect 411898 443680 411904 443692
rect 99248 443652 411904 443680
rect 99248 443640 99254 443652
rect 411898 443640 411904 443652
rect 411956 443640 411962 443692
rect 317414 442280 317420 442332
rect 317472 442320 317478 442332
rect 500954 442320 500960 442332
rect 317472 442292 500960 442320
rect 317472 442280 317478 442292
rect 500954 442280 500960 442292
rect 501012 442280 501018 442332
rect 97902 442212 97908 442264
rect 97960 442252 97966 442264
rect 411806 442252 411812 442264
rect 97960 442224 411812 442252
rect 97960 442212 97966 442224
rect 411806 442212 411812 442224
rect 411864 442212 411870 442264
rect 310882 440920 310888 440972
rect 310940 440960 310946 440972
rect 479518 440960 479524 440972
rect 310940 440932 479524 440960
rect 310940 440920 310946 440932
rect 479518 440920 479524 440932
rect 479576 440920 479582 440972
rect 99282 440852 99288 440904
rect 99340 440892 99346 440904
rect 357986 440892 357992 440904
rect 99340 440864 357992 440892
rect 99340 440852 99346 440864
rect 357986 440852 357992 440864
rect 358044 440852 358050 440904
rect 314654 439560 314660 439612
rect 314712 439600 314718 439612
rect 494698 439600 494704 439612
rect 314712 439572 494704 439600
rect 314712 439560 314718 439572
rect 494698 439560 494704 439572
rect 494756 439560 494762 439612
rect 104802 439492 104808 439544
rect 104860 439532 104866 439544
rect 410150 439532 410156 439544
rect 104860 439504 410156 439532
rect 104860 439492 104866 439504
rect 410150 439492 410156 439504
rect 410208 439492 410214 439544
rect 307846 438200 307852 438252
rect 307904 438240 307910 438252
rect 492674 438240 492680 438252
rect 307904 438212 492680 438240
rect 307904 438200 307910 438212
rect 492674 438200 492680 438212
rect 492732 438200 492738 438252
rect 143442 438132 143448 438184
rect 143500 438172 143506 438184
rect 394694 438172 394700 438184
rect 143500 438144 394700 438172
rect 143500 438132 143506 438144
rect 394694 438132 394700 438144
rect 394752 438132 394758 438184
rect 303890 436840 303896 436892
rect 303948 436880 303954 436892
rect 489914 436880 489920 436892
rect 303948 436852 489920 436880
rect 303948 436840 303954 436852
rect 489914 436840 489920 436852
rect 489972 436840 489978 436892
rect 142062 436772 142068 436824
rect 142120 436812 142126 436824
rect 409414 436812 409420 436824
rect 142120 436784 409420 436812
rect 142120 436772 142126 436784
rect 409414 436772 409420 436784
rect 409472 436772 409478 436824
rect 88242 436704 88248 436756
rect 88300 436744 88306 436756
rect 411714 436744 411720 436756
rect 88300 436716 411720 436744
rect 88300 436704 88306 436716
rect 411714 436704 411720 436716
rect 411772 436704 411778 436756
rect 269114 435412 269120 435464
rect 269172 435452 269178 435464
rect 465074 435452 465080 435464
rect 269172 435424 465080 435452
rect 269172 435412 269178 435424
rect 465074 435412 465080 435424
rect 465132 435412 465138 435464
rect 85482 435344 85488 435396
rect 85540 435384 85546 435396
rect 411254 435384 411260 435396
rect 85540 435356 411260 435384
rect 85540 435344 85546 435356
rect 411254 435344 411260 435356
rect 411312 435344 411318 435396
rect 262214 434052 262220 434104
rect 262272 434092 262278 434104
rect 460934 434092 460940 434104
rect 262272 434064 460940 434092
rect 262272 434052 262278 434064
rect 460934 434052 460940 434064
rect 460992 434052 460998 434104
rect 81158 433984 81164 434036
rect 81216 434024 81222 434036
rect 335354 434024 335360 434036
rect 81216 433996 335360 434024
rect 81216 433984 81222 433996
rect 335354 433984 335360 433996
rect 335412 433984 335418 434036
rect 265434 432692 265440 432744
rect 265492 432732 265498 432744
rect 457438 432732 457444 432744
rect 265492 432704 457444 432732
rect 265492 432692 265498 432704
rect 457438 432692 457444 432704
rect 457496 432692 457502 432744
rect 111702 432624 111708 432676
rect 111760 432664 111766 432676
rect 410518 432664 410524 432676
rect 111760 432636 410524 432664
rect 111760 432624 111766 432636
rect 410518 432624 410524 432636
rect 410576 432624 410582 432676
rect 82722 432556 82728 432608
rect 82780 432596 82786 432608
rect 411346 432596 411352 432608
rect 82780 432568 411352 432596
rect 82780 432556 82786 432568
rect 411346 432556 411352 432568
rect 411404 432556 411410 432608
rect 258442 431332 258448 431384
rect 258500 431372 258506 431384
rect 458174 431372 458180 431384
rect 258500 431344 458180 431372
rect 258500 431332 258506 431344
rect 458174 431332 458180 431344
rect 458232 431332 458238 431384
rect 108942 431264 108948 431316
rect 109000 431304 109006 431316
rect 410242 431304 410248 431316
rect 109000 431276 410248 431304
rect 109000 431264 109006 431276
rect 410242 431264 410248 431276
rect 410300 431264 410306 431316
rect 96522 431196 96528 431248
rect 96580 431236 96586 431248
rect 411622 431236 411628 431248
rect 96580 431208 411628 431236
rect 96580 431196 96586 431208
rect 411622 431196 411628 431208
rect 411680 431196 411686 431248
rect 560938 430584 560944 430636
rect 560996 430624 561002 430636
rect 580166 430624 580172 430636
rect 560996 430596 580172 430624
rect 560996 430584 561002 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 251450 429972 251456 430024
rect 251508 430012 251514 430024
rect 452654 430012 452660 430024
rect 251508 429984 452660 430012
rect 251508 429972 251514 429984
rect 452654 429972 452660 429984
rect 452712 429972 452718 430024
rect 93762 429904 93768 429956
rect 93820 429944 93826 429956
rect 411438 429944 411444 429956
rect 93820 429916 411444 429944
rect 93820 429904 93826 429916
rect 411438 429904 411444 429916
rect 411496 429904 411502 429956
rect 47762 429836 47768 429888
rect 47820 429876 47826 429888
rect 409966 429876 409972 429888
rect 47820 429848 409972 429876
rect 47820 429836 47826 429848
rect 409966 429836 409972 429848
rect 410024 429836 410030 429888
rect 397362 428612 397368 428664
rect 397420 428652 397426 428664
rect 445754 428652 445760 428664
rect 397420 428624 445760 428652
rect 397420 428612 397426 428624
rect 445754 428612 445760 428624
rect 445812 428612 445818 428664
rect 200850 428544 200856 428596
rect 200908 428584 200914 428596
rect 416774 428584 416780 428596
rect 200908 428556 416780 428584
rect 200908 428544 200914 428556
rect 416774 428544 416780 428556
rect 416832 428544 416838 428596
rect 67542 428476 67548 428528
rect 67600 428516 67606 428528
rect 410058 428516 410064 428528
rect 67600 428488 410064 428516
rect 67600 428476 67606 428488
rect 410058 428476 410064 428488
rect 410116 428476 410122 428528
rect 49602 428408 49608 428460
rect 49660 428448 49666 428460
rect 411530 428448 411536 428460
rect 49660 428420 411536 428448
rect 49660 428408 49666 428420
rect 411530 428408 411536 428420
rect 411588 428408 411594 428460
rect 284570 427388 284576 427440
rect 284628 427428 284634 427440
rect 444374 427428 444380 427440
rect 284628 427400 444380 427428
rect 284628 427388 284634 427400
rect 444374 427388 444380 427400
rect 444432 427388 444438 427440
rect 277578 427320 277584 427372
rect 277636 427360 277642 427372
rect 441614 427360 441620 427372
rect 277636 427332 441620 427360
rect 277636 427320 277642 427332
rect 441614 427320 441620 427332
rect 441672 427320 441678 427372
rect 270586 427252 270592 427304
rect 270644 427292 270650 427304
rect 440326 427292 440332 427304
rect 270644 427264 440332 427292
rect 270644 427252 270650 427264
rect 440326 427252 440332 427264
rect 440384 427252 440390 427304
rect 267090 427184 267096 427236
rect 267148 427224 267154 427236
rect 438854 427224 438860 427236
rect 267148 427196 438860 427224
rect 267148 427184 267154 427196
rect 438854 427184 438860 427196
rect 438912 427184 438918 427236
rect 260282 427116 260288 427168
rect 260340 427156 260346 427168
rect 436094 427156 436100 427168
rect 260340 427128 436100 427156
rect 260340 427116 260346 427128
rect 436094 427116 436100 427128
rect 436152 427116 436158 427168
rect 84010 427048 84016 427100
rect 84068 427088 84074 427100
rect 359366 427088 359372 427100
rect 84068 427060 359372 427088
rect 84068 427048 84074 427060
rect 359366 427048 359372 427060
rect 359424 427048 359430 427100
rect 256786 426232 256792 426284
rect 256844 426272 256850 426284
rect 434714 426272 434720 426284
rect 256844 426244 434720 426272
rect 256844 426232 256850 426244
rect 434714 426232 434720 426244
rect 434772 426232 434778 426284
rect 248506 426164 248512 426216
rect 248564 426204 248570 426216
rect 449894 426204 449900 426216
rect 248564 426176 449900 426204
rect 248564 426164 248570 426176
rect 449894 426164 449900 426176
rect 449952 426164 449958 426216
rect 218606 426096 218612 426148
rect 218664 426136 218670 426148
rect 420914 426136 420920 426148
rect 218664 426108 420920 426136
rect 218664 426096 218670 426108
rect 420914 426096 420920 426108
rect 420972 426096 420978 426148
rect 244458 426028 244464 426080
rect 244516 426068 244522 426080
rect 447134 426068 447140 426080
rect 244516 426040 447140 426068
rect 244516 426028 244522 426040
rect 447134 426028 447140 426040
rect 447192 426028 447198 426080
rect 239306 425960 239312 426012
rect 239364 426000 239370 426012
rect 445938 426000 445944 426012
rect 239364 425972 445944 426000
rect 239364 425960 239370 425972
rect 445938 425960 445944 425972
rect 445996 425960 446002 426012
rect 233970 425892 233976 425944
rect 234028 425932 234034 425944
rect 442994 425932 443000 425944
rect 234028 425904 443000 425932
rect 234028 425892 234034 425904
rect 442994 425892 443000 425904
rect 443052 425892 443058 425944
rect 229094 425824 229100 425876
rect 229152 425864 229158 425876
rect 440234 425864 440240 425876
rect 229152 425836 440240 425864
rect 229152 425824 229158 425836
rect 440234 425824 440240 425836
rect 440292 425824 440298 425876
rect 223574 425756 223580 425808
rect 223632 425796 223638 425808
rect 437474 425796 437480 425808
rect 223632 425768 437480 425796
rect 223632 425756 223638 425768
rect 437474 425756 437480 425768
rect 437532 425756 437538 425808
rect 197998 425688 198004 425740
rect 198056 425728 198062 425740
rect 418154 425728 418160 425740
rect 198056 425700 418160 425728
rect 198056 425688 198062 425700
rect 418154 425688 418160 425700
rect 418212 425688 418218 425740
rect 300670 424940 300676 424992
rect 300728 424980 300734 424992
rect 488534 424980 488540 424992
rect 300728 424952 488540 424980
rect 300728 424940 300734 424952
rect 488534 424940 488540 424952
rect 488592 424940 488598 424992
rect 297634 424872 297640 424924
rect 297692 424912 297698 424924
rect 485774 424912 485780 424924
rect 297692 424884 485780 424912
rect 297692 424872 297698 424884
rect 485774 424872 485780 424884
rect 485832 424872 485838 424924
rect 290642 424804 290648 424856
rect 290700 424844 290706 424856
rect 480254 424844 480260 424856
rect 290700 424816 480260 424844
rect 290700 424804 290706 424816
rect 480254 424804 480260 424816
rect 480312 424804 480318 424856
rect 293862 424736 293868 424788
rect 293920 424776 293926 424788
rect 483014 424776 483020 424788
rect 293920 424748 483020 424776
rect 293920 424736 293926 424748
rect 483014 424736 483020 424748
rect 483072 424736 483078 424788
rect 283650 424668 283656 424720
rect 283708 424708 283714 424720
rect 474734 424708 474740 424720
rect 283708 424680 474740 424708
rect 283708 424668 283714 424680
rect 474734 424668 474740 424680
rect 474792 424668 474798 424720
rect 286962 424600 286968 424652
rect 287020 424640 287026 424652
rect 477494 424640 477500 424652
rect 287020 424612 477500 424640
rect 287020 424600 287026 424612
rect 477494 424600 477500 424612
rect 477552 424600 477558 424652
rect 276658 424532 276664 424584
rect 276716 424572 276722 424584
rect 470594 424572 470600 424584
rect 276716 424544 470600 424572
rect 276716 424532 276722 424544
rect 470594 424532 470600 424544
rect 470652 424532 470658 424584
rect 279970 424464 279976 424516
rect 280028 424504 280034 424516
rect 473354 424504 473360 424516
rect 280028 424476 473360 424504
rect 280028 424464 280034 424476
rect 473354 424464 473360 424476
rect 473412 424464 473418 424516
rect 273162 424396 273168 424448
rect 273220 424436 273226 424448
rect 467834 424436 467840 424448
rect 273220 424408 467840 424436
rect 273220 424396 273226 424408
rect 467834 424396 467840 424408
rect 467892 424396 467898 424448
rect 78582 424328 78588 424380
rect 78640 424368 78646 424380
rect 185670 424368 185676 424380
rect 78640 424340 185676 424368
rect 78640 424328 78646 424340
rect 185670 424328 185676 424340
rect 185728 424328 185734 424380
rect 203242 424328 203248 424380
rect 203300 424368 203306 424380
rect 430666 424368 430672 424380
rect 203300 424340 430672 424368
rect 203300 424328 203306 424340
rect 430666 424328 430672 424340
rect 430724 424328 430730 424380
rect 73062 423580 73068 423632
rect 73120 423620 73126 423632
rect 218606 423620 218612 423632
rect 73120 423592 218612 423620
rect 73120 423580 73126 423592
rect 218606 423580 218612 423592
rect 218664 423580 218670 423632
rect 342898 423580 342904 423632
rect 342956 423620 342962 423632
rect 344094 423620 344100 423632
rect 342956 423592 344100 423620
rect 342956 423580 342962 423592
rect 344094 423580 344100 423592
rect 344152 423580 344158 423632
rect 407758 423580 407764 423632
rect 407816 423620 407822 423632
rect 408678 423620 408684 423632
rect 407816 423592 408684 423620
rect 407816 423580 407822 423592
rect 408678 423580 408684 423592
rect 408736 423580 408742 423632
rect 71682 423512 71688 423564
rect 71740 423552 71746 423564
rect 211798 423552 211804 423564
rect 71740 423524 211804 423552
rect 71740 423512 71746 423524
rect 211798 423512 211804 423524
rect 211856 423512 211862 423564
rect 70302 423444 70308 423496
rect 70360 423484 70366 423496
rect 204898 423484 204904 423496
rect 70360 423456 204904 423484
rect 70360 423444 70366 423456
rect 204898 423444 204904 423456
rect 204956 423444 204962 423496
rect 68922 423376 68928 423428
rect 68980 423416 68986 423428
rect 197998 423416 198004 423428
rect 68980 423388 198004 423416
rect 68980 423376 68986 423388
rect 197998 423376 198004 423388
rect 198056 423376 198062 423428
rect 363874 423240 363880 423292
rect 363932 423280 363938 423292
rect 410334 423280 410340 423292
rect 363932 423252 410340 423280
rect 363932 423240 363938 423252
rect 410334 423240 410340 423252
rect 410392 423240 410398 423292
rect 250530 423172 250536 423224
rect 250588 423212 250594 423224
rect 428458 423212 428464 423224
rect 250588 423184 428464 423212
rect 250588 423172 250594 423184
rect 428458 423172 428464 423184
rect 428516 423172 428522 423224
rect 241330 423104 241336 423156
rect 241388 423144 241394 423156
rect 427078 423144 427084 423156
rect 241388 423116 427084 423144
rect 241388 423104 241394 423116
rect 427078 423104 427084 423116
rect 427136 423104 427142 423156
rect 146202 423036 146208 423088
rect 146260 423076 146266 423088
rect 396534 423076 396540 423088
rect 146260 423048 396540 423076
rect 146260 423036 146266 423048
rect 396534 423036 396540 423048
rect 396592 423036 396598 423088
rect 79318 422968 79324 423020
rect 79376 423008 79382 423020
rect 330110 423008 330116 423020
rect 79376 422980 330116 423008
rect 79376 422968 79382 422980
rect 330110 422968 330116 422980
rect 330168 422968 330174 423020
rect 359458 422968 359464 423020
rect 359516 423008 359522 423020
rect 403526 423008 403532 423020
rect 359516 422980 403532 423008
rect 359516 422968 359522 422980
rect 403526 422968 403532 422980
rect 403584 422968 403590 423020
rect 126882 422900 126888 422952
rect 126940 422940 126946 422952
rect 382550 422940 382556 422952
rect 126940 422912 382556 422940
rect 126940 422900 126946 422912
rect 382550 422900 382556 422912
rect 382608 422900 382614 422952
rect 365622 422832 365628 422884
rect 365680 422872 365686 422884
rect 419534 422872 419540 422884
rect 365680 422844 419540 422872
rect 365680 422832 365686 422844
rect 419534 422832 419540 422844
rect 419592 422832 419598 422884
rect 398742 422764 398748 422816
rect 398800 422804 398806 422816
rect 412726 422804 412732 422816
rect 398800 422776 412732 422804
rect 398800 422764 398806 422776
rect 412726 422764 412732 422776
rect 412784 422764 412790 422816
rect 386230 422696 386236 422748
rect 386288 422736 386294 422748
rect 412634 422736 412640 422748
rect 386288 422708 412640 422736
rect 386288 422696 386294 422708
rect 412634 422696 412640 422708
rect 412692 422696 412698 422748
rect 374362 422628 374368 422680
rect 374420 422668 374426 422680
rect 416130 422668 416136 422680
rect 374420 422640 416136 422668
rect 374420 422628 374426 422640
rect 416130 422628 416136 422640
rect 416188 422628 416194 422680
rect 405642 422560 405648 422612
rect 405700 422600 405706 422612
rect 418982 422600 418988 422612
rect 405700 422572 418988 422600
rect 405700 422560 405706 422572
rect 418982 422560 418988 422572
rect 419040 422560 419046 422612
rect 334250 422492 334256 422544
rect 334308 422532 334314 422544
rect 351086 422532 351092 422544
rect 334308 422504 351092 422532
rect 334308 422492 334314 422504
rect 351086 422492 351092 422504
rect 351144 422492 351150 422544
rect 362218 422492 362224 422544
rect 362276 422532 362282 422544
rect 416038 422532 416044 422544
rect 362276 422504 416044 422532
rect 362276 422492 362282 422504
rect 416038 422492 416044 422504
rect 416096 422492 416102 422544
rect 351730 422424 351736 422476
rect 351788 422464 351794 422476
rect 360102 422464 360108 422476
rect 351788 422436 360108 422464
rect 351788 422424 351794 422436
rect 360102 422424 360108 422436
rect 360160 422424 360166 422476
rect 377858 422424 377864 422476
rect 377916 422464 377922 422476
rect 431310 422464 431316 422476
rect 377916 422436 431316 422464
rect 377916 422424 377922 422436
rect 431310 422424 431316 422436
rect 431368 422424 431374 422476
rect 186222 422356 186228 422408
rect 186280 422396 186286 422408
rect 347774 422396 347780 422408
rect 186280 422368 347780 422396
rect 186280 422356 186286 422368
rect 347774 422356 347780 422368
rect 347832 422356 347838 422408
rect 353202 422356 353208 422408
rect 353260 422396 353266 422408
rect 420178 422396 420184 422408
rect 353260 422368 420184 422396
rect 353260 422356 353266 422368
rect 420178 422356 420184 422368
rect 420236 422356 420242 422408
rect 188890 422288 188896 422340
rect 188948 422328 188954 422340
rect 368566 422328 368572 422340
rect 188948 422300 368572 422328
rect 188948 422288 188954 422300
rect 368566 422288 368572 422300
rect 368624 422288 368630 422340
rect 435358 422328 435364 422340
rect 408788 422300 435364 422328
rect 407666 422220 407672 422272
rect 407724 422260 407730 422272
rect 408788 422260 408816 422300
rect 435358 422288 435364 422300
rect 435416 422288 435422 422340
rect 407724 422232 408816 422260
rect 407724 422220 407730 422232
rect 360102 421540 360108 421592
rect 360160 421580 360166 421592
rect 552014 421580 552020 421592
rect 360160 421552 552020 421580
rect 360160 421540 360166 421552
rect 552014 421540 552020 421552
rect 552072 421540 552078 421592
rect 186958 421472 186964 421524
rect 187016 421512 187022 421524
rect 552198 421512 552204 421524
rect 187016 421484 552204 421512
rect 187016 421472 187022 421484
rect 552198 421472 552204 421484
rect 552256 421472 552262 421524
rect 388346 421404 388352 421456
rect 388404 421444 388410 421456
rect 418798 421444 418804 421456
rect 388404 421416 418804 421444
rect 388404 421404 388410 421416
rect 418798 421404 418804 421416
rect 418856 421404 418862 421456
rect 376202 421336 376208 421388
rect 376260 421376 376266 421388
rect 417418 421376 417424 421388
rect 376260 421348 417424 421376
rect 376260 421336 376266 421348
rect 417418 421336 417424 421348
rect 417476 421336 417482 421388
rect 355226 421268 355232 421320
rect 355284 421308 355290 421320
rect 413278 421308 413284 421320
rect 355284 421280 413284 421308
rect 355284 421268 355290 421280
rect 413278 421268 413284 421280
rect 413336 421268 413342 421320
rect 346302 421200 346308 421252
rect 346360 421240 346366 421252
rect 413554 421240 413560 421252
rect 346360 421212 413560 421240
rect 346360 421200 346366 421212
rect 413554 421200 413560 421212
rect 413612 421200 413618 421252
rect 349890 421132 349896 421184
rect 349948 421172 349954 421184
rect 429194 421172 429200 421184
rect 349948 421144 429200 421172
rect 349948 421132 349954 421144
rect 429194 421132 429200 421144
rect 429252 421132 429258 421184
rect 169754 421064 169760 421116
rect 169812 421104 169818 421116
rect 391198 421104 391204 421116
rect 169812 421076 391204 421104
rect 169812 421064 169818 421076
rect 391198 421064 391204 421076
rect 391256 421064 391262 421116
rect 393682 421064 393688 421116
rect 393740 421104 393746 421116
rect 438118 421104 438124 421116
rect 393740 421076 438124 421104
rect 393740 421064 393746 421076
rect 438118 421064 438124 421076
rect 438176 421064 438182 421116
rect 329098 420996 329104 421048
rect 329156 421036 329162 421048
rect 551278 421036 551284 421048
rect 329156 421008 551284 421036
rect 329156 420996 329162 421008
rect 551278 420996 551284 421008
rect 551336 420996 551342 421048
rect 402330 420928 402336 420980
rect 402388 420968 402394 420980
rect 414750 420968 414756 420980
rect 402388 420940 414756 420968
rect 402388 420928 402394 420940
rect 414750 420928 414756 420940
rect 414808 420928 414814 420980
rect 367370 420316 367376 420368
rect 367428 420356 367434 420368
rect 482278 420356 482284 420368
rect 367428 420328 482284 420356
rect 367428 420316 367434 420328
rect 482278 420316 482284 420328
rect 482336 420316 482342 420368
rect 187510 420248 187516 420300
rect 187568 420288 187574 420300
rect 413370 420288 413376 420300
rect 187568 420260 413376 420288
rect 187568 420248 187574 420260
rect 413370 420248 413376 420260
rect 413428 420248 413434 420300
rect 190362 420180 190368 420232
rect 190420 420220 190426 420232
rect 413462 420220 413468 420232
rect 190420 420192 413468 420220
rect 190420 420180 190426 420192
rect 413462 420180 413468 420192
rect 413520 420180 413526 420232
rect 187050 420112 187056 420164
rect 187108 420152 187114 420164
rect 414658 420152 414664 420164
rect 187108 420124 414664 420152
rect 187108 420112 187114 420124
rect 414658 420112 414664 420124
rect 414716 420112 414722 420164
rect 190730 420044 190736 420096
rect 190788 420084 190794 420096
rect 414842 420084 414848 420096
rect 190788 420056 414848 420084
rect 190788 420044 190794 420056
rect 414842 420044 414848 420056
rect 414900 420044 414906 420096
rect 187326 419976 187332 420028
rect 187384 420016 187390 420028
rect 421650 420016 421656 420028
rect 187384 419988 421656 420016
rect 187384 419976 187390 419988
rect 421650 419976 421656 419988
rect 421708 419976 421714 420028
rect 187142 419908 187148 419960
rect 187200 419948 187206 419960
rect 424410 419948 424416 419960
rect 187200 419920 424416 419948
rect 187200 419908 187206 419920
rect 424410 419908 424416 419920
rect 424468 419908 424474 419960
rect 187234 419840 187240 419892
rect 187292 419880 187298 419892
rect 428550 419880 428556 419892
rect 187292 419852 428556 419880
rect 187292 419840 187298 419852
rect 428550 419840 428556 419852
rect 428608 419840 428614 419892
rect 372522 419772 372528 419824
rect 372580 419812 372586 419824
rect 550634 419812 550640 419824
rect 372580 419784 550640 419812
rect 372580 419772 372586 419784
rect 550634 419772 550640 419784
rect 550692 419772 550698 419824
rect 131942 419704 131948 419756
rect 132000 419744 132006 419756
rect 425882 419744 425888 419756
rect 132000 419716 425888 419744
rect 132000 419704 132006 419716
rect 425882 419704 425888 419716
rect 425940 419704 425946 419756
rect 189350 419636 189356 419688
rect 189408 419676 189414 419688
rect 494514 419676 494520 419688
rect 189408 419648 494520 419676
rect 189408 419636 189414 419648
rect 494514 419636 494520 419648
rect 494572 419636 494578 419688
rect 189074 419568 189080 419620
rect 189132 419608 189138 419620
rect 552290 419608 552296 419620
rect 189132 419580 552296 419608
rect 189132 419568 189138 419580
rect 552290 419568 552296 419580
rect 552348 419568 552354 419620
rect 187418 419500 187424 419552
rect 187476 419540 187482 419552
rect 552106 419540 552112 419552
rect 187476 419512 552112 419540
rect 187476 419500 187482 419512
rect 552106 419500 552112 419512
rect 552164 419500 552170 419552
rect 107562 419432 107568 419484
rect 107620 419472 107626 419484
rect 186314 419472 186320 419484
rect 107620 419444 186320 419472
rect 107620 419432 107626 419444
rect 186314 419432 186320 419444
rect 186372 419432 186378 419484
rect 412082 418888 412088 418940
rect 412140 418928 412146 418940
rect 413830 418928 413836 418940
rect 412140 418900 413836 418928
rect 412140 418888 412146 418900
rect 413830 418888 413836 418900
rect 413888 418888 413894 418940
rect 412634 418752 412640 418804
rect 412692 418792 412698 418804
rect 506750 418792 506756 418804
rect 412692 418764 506756 418792
rect 412692 418752 412698 418764
rect 506750 418752 506756 418764
rect 506808 418752 506814 418804
rect 549898 418140 549904 418192
rect 549956 418180 549962 418192
rect 580166 418180 580172 418192
rect 549956 418152 580172 418180
rect 549956 418140 549962 418152
rect 580166 418140 580172 418152
rect 580224 418140 580230 418192
rect 412726 417392 412732 417444
rect 412784 417432 412790 417444
rect 531314 417432 531320 417444
rect 412784 417404 531320 417432
rect 412784 417392 412790 417404
rect 531314 417392 531320 417404
rect 531372 417392 531378 417444
rect 412082 416848 412088 416900
rect 412140 416888 412146 416900
rect 413646 416888 413652 416900
rect 412140 416860 413652 416888
rect 412140 416848 412146 416860
rect 413646 416848 413652 416860
rect 413704 416848 413710 416900
rect 75822 416032 75828 416084
rect 75880 416072 75886 416084
rect 178678 416072 178684 416084
rect 75880 416044 178684 416072
rect 75880 416032 75886 416044
rect 178678 416032 178684 416044
rect 178736 416032 178742 416084
rect 187418 414128 187424 414180
rect 187476 414128 187482 414180
rect 173158 413992 173164 414044
rect 173216 414032 173222 414044
rect 186314 414032 186320 414044
rect 173216 414004 186320 414032
rect 173216 413992 173222 414004
rect 186314 413992 186320 414004
rect 186372 413992 186378 414044
rect 187436 413976 187464 414128
rect 187418 413924 187424 413976
rect 187476 413924 187482 413976
rect 186958 413788 186964 413840
rect 187016 413828 187022 413840
rect 187234 413828 187240 413840
rect 187016 413800 187240 413828
rect 187016 413788 187022 413800
rect 187234 413788 187240 413800
rect 187292 413788 187298 413840
rect 106182 413244 106188 413296
rect 106240 413284 106246 413296
rect 180058 413284 180064 413296
rect 106240 413256 180064 413284
rect 106240 413244 106246 413256
rect 180058 413244 180064 413256
rect 180116 413244 180122 413296
rect 139302 412564 139308 412616
rect 139360 412604 139366 412616
rect 186314 412604 186320 412616
rect 139360 412576 186320 412604
rect 139360 412564 139366 412576
rect 186314 412564 186320 412576
rect 186372 412564 186378 412616
rect 413554 411952 413560 412004
rect 413612 411992 413618 412004
rect 470134 411992 470140 412004
rect 413612 411964 470140 411992
rect 413612 411952 413618 411964
rect 470134 411952 470140 411964
rect 470192 411952 470198 412004
rect 414842 411884 414848 411936
rect 414900 411924 414906 411936
rect 543734 411924 543740 411936
rect 414900 411896 543740 411924
rect 414900 411884 414906 411896
rect 543734 411884 543740 411896
rect 543792 411884 543798 411936
rect 439498 411340 439504 411392
rect 439556 411380 439562 411392
rect 445754 411380 445760 411392
rect 439556 411352 445760 411380
rect 439556 411340 439562 411352
rect 445754 411340 445760 411352
rect 445812 411340 445818 411392
rect 418890 411272 418896 411324
rect 418948 411312 418954 411324
rect 458266 411312 458272 411324
rect 418948 411284 458272 411312
rect 418948 411272 418954 411284
rect 458266 411272 458272 411284
rect 458324 411272 458330 411324
rect 136542 411204 136548 411256
rect 136600 411244 136606 411256
rect 186406 411244 186412 411256
rect 136600 411216 186412 411244
rect 136600 411204 136606 411216
rect 186406 411204 186412 411216
rect 186464 411204 186470 411256
rect 171042 409844 171048 409896
rect 171100 409884 171106 409896
rect 186314 409884 186320 409896
rect 171100 409856 186320 409884
rect 171100 409844 171106 409856
rect 186314 409844 186320 409856
rect 186372 409844 186378 409896
rect 417510 409844 417516 409896
rect 417568 409884 417574 409896
rect 519078 409884 519084 409896
rect 417568 409856 519084 409884
rect 417568 409844 417574 409856
rect 519078 409844 519084 409856
rect 519136 409844 519142 409896
rect 413646 409776 413652 409828
rect 413704 409816 413710 409828
rect 437474 409816 437480 409828
rect 413704 409788 437480 409816
rect 413704 409776 413710 409788
rect 437474 409776 437480 409788
rect 437532 409776 437538 409828
rect 95142 409096 95148 409148
rect 95200 409136 95206 409148
rect 188430 409136 188436 409148
rect 95200 409108 188436 409136
rect 95200 409096 95206 409108
rect 188430 409096 188436 409108
rect 188488 409096 188494 409148
rect 414750 408416 414756 408468
rect 414808 408456 414814 408468
rect 437474 408456 437480 408468
rect 414808 408428 437480 408456
rect 414808 408416 414814 408428
rect 437474 408416 437480 408428
rect 437532 408416 437538 408468
rect 91002 407736 91008 407788
rect 91060 407776 91066 407788
rect 188522 407776 188528 407788
rect 91060 407748 188528 407776
rect 91060 407736 91066 407748
rect 188522 407736 188528 407748
rect 188580 407736 188586 407788
rect 129642 407056 129648 407108
rect 129700 407096 129706 407108
rect 186314 407096 186320 407108
rect 129700 407068 186320 407096
rect 129700 407056 129706 407068
rect 186314 407056 186320 407068
rect 186372 407056 186378 407108
rect 413462 407056 413468 407108
rect 413520 407096 413526 407108
rect 437474 407096 437480 407108
rect 413520 407068 437480 407096
rect 413520 407056 413526 407068
rect 437474 407056 437480 407068
rect 437532 407056 437538 407108
rect 66162 406376 66168 406428
rect 66220 406416 66226 406428
rect 164878 406416 164884 406428
rect 66220 406388 164884 406416
rect 66220 406376 66226 406388
rect 164878 406376 164884 406388
rect 164936 406376 164942 406428
rect 84102 404948 84108 405000
rect 84160 404988 84166 405000
rect 189902 404988 189908 405000
rect 84160 404960 189908 404988
rect 84160 404948 84166 404960
rect 189902 404948 189908 404960
rect 189960 404948 189966 405000
rect 124122 404268 124128 404320
rect 124180 404308 124186 404320
rect 186314 404308 186320 404320
rect 124180 404280 186320 404308
rect 124180 404268 124186 404280
rect 186314 404268 186320 404280
rect 186372 404268 186378 404320
rect 413370 404268 413376 404320
rect 413428 404308 413434 404320
rect 437474 404308 437480 404320
rect 413428 404280 437480 404308
rect 413428 404268 413434 404280
rect 437474 404268 437480 404280
rect 437532 404268 437538 404320
rect 1302 401616 1308 401668
rect 1360 401656 1366 401668
rect 53834 401656 53840 401668
rect 1360 401628 53840 401656
rect 1360 401616 1366 401628
rect 53834 401616 53840 401628
rect 53892 401656 53898 401668
rect 54938 401656 54944 401668
rect 53892 401628 54944 401656
rect 53892 401616 53898 401628
rect 54938 401616 54944 401628
rect 54996 401616 55002 401668
rect 104894 401616 104900 401668
rect 104952 401656 104958 401668
rect 189994 401656 190000 401668
rect 104952 401628 190000 401656
rect 104952 401616 104958 401628
rect 189994 401616 190000 401628
rect 190052 401616 190058 401668
rect 432598 401616 432604 401668
rect 432656 401656 432662 401668
rect 437474 401656 437480 401668
rect 432656 401628 437480 401656
rect 432656 401616 432662 401628
rect 437474 401616 437480 401628
rect 437532 401616 437538 401668
rect 121362 401548 121368 401600
rect 121420 401588 121426 401600
rect 186314 401588 186320 401600
rect 121420 401560 186320 401588
rect 121420 401548 121426 401560
rect 186314 401548 186320 401560
rect 186372 401548 186378 401600
rect 48222 400868 48228 400920
rect 48280 400908 48286 400920
rect 184290 400908 184296 400920
rect 48280 400880 184296 400908
rect 48280 400868 48286 400880
rect 184290 400868 184296 400880
rect 184348 400868 184354 400920
rect 413462 400188 413468 400240
rect 413520 400228 413526 400240
rect 437474 400228 437480 400240
rect 413520 400200 437480 400228
rect 413520 400188 413526 400200
rect 437474 400188 437480 400200
rect 437532 400188 437538 400240
rect 131206 398828 131212 398880
rect 131264 398868 131270 398880
rect 144178 398868 144184 398880
rect 131264 398840 144184 398868
rect 131264 398828 131270 398840
rect 144178 398828 144184 398840
rect 144236 398828 144242 398880
rect 425698 398828 425704 398880
rect 425756 398868 425762 398880
rect 437474 398868 437480 398880
rect 425756 398840 437480 398868
rect 425756 398828 425762 398840
rect 437474 398828 437480 398840
rect 437532 398828 437538 398880
rect 414658 398760 414664 398812
rect 414716 398800 414722 398812
rect 437566 398800 437572 398812
rect 414716 398772 437572 398800
rect 414716 398760 414722 398772
rect 437566 398760 437572 398772
rect 437624 398760 437630 398812
rect 131206 397468 131212 397520
rect 131264 397508 131270 397520
rect 142798 397508 142804 397520
rect 131264 397480 142804 397508
rect 131264 397468 131270 397480
rect 142798 397468 142804 397480
rect 142856 397468 142862 397520
rect 131206 396176 131212 396228
rect 131264 396216 131270 396228
rect 140222 396216 140228 396228
rect 131264 396188 140228 396216
rect 131264 396176 131270 396188
rect 140222 396176 140228 396188
rect 140280 396176 140286 396228
rect 131482 396108 131488 396160
rect 131540 396148 131546 396160
rect 141510 396148 141516 396160
rect 131540 396120 141516 396148
rect 131540 396108 131546 396120
rect 141510 396108 141516 396120
rect 141568 396108 141574 396160
rect 131298 396040 131304 396092
rect 131356 396080 131362 396092
rect 183002 396080 183008 396092
rect 131356 396052 183008 396080
rect 131356 396040 131362 396052
rect 183002 396040 183008 396052
rect 183060 396040 183066 396092
rect 162118 395972 162124 396024
rect 162176 396012 162182 396024
rect 186314 396012 186320 396024
rect 162176 395984 186320 396012
rect 162176 395972 162182 395984
rect 186314 395972 186320 395984
rect 186372 395972 186378 396024
rect 131206 394748 131212 394800
rect 131264 394788 131270 394800
rect 162210 394788 162216 394800
rect 131264 394760 162216 394788
rect 131264 394748 131270 394760
rect 162210 394748 162216 394760
rect 162268 394748 162274 394800
rect 131298 394680 131304 394732
rect 131356 394720 131362 394732
rect 174538 394720 174544 394732
rect 131356 394692 174544 394720
rect 131356 394680 131362 394692
rect 174538 394680 174544 394692
rect 174596 394680 174602 394732
rect 131206 393388 131212 393440
rect 131264 393428 131270 393440
rect 160738 393428 160744 393440
rect 131264 393400 160744 393428
rect 131264 393388 131270 393400
rect 160738 393388 160744 393400
rect 160796 393388 160802 393440
rect 132034 393320 132040 393372
rect 132092 393360 132098 393372
rect 181530 393360 181536 393372
rect 132092 393332 181536 393360
rect 132092 393320 132098 393332
rect 181530 393320 181536 393332
rect 181588 393320 181594 393372
rect 177390 393252 177396 393304
rect 177448 393292 177454 393304
rect 186314 393292 186320 393304
rect 177448 393264 186320 393292
rect 177448 393252 177454 393264
rect 186314 393252 186320 393264
rect 186372 393252 186378 393304
rect 413278 393252 413284 393304
rect 413336 393292 413342 393304
rect 437474 393292 437480 393304
rect 413336 393264 437480 393292
rect 413336 393252 413342 393264
rect 437474 393252 437480 393264
rect 437532 393252 437538 393304
rect 132034 392028 132040 392080
rect 132092 392068 132098 392080
rect 137462 392068 137468 392080
rect 132092 392040 137468 392068
rect 132092 392028 132098 392040
rect 137462 392028 137468 392040
rect 137520 392028 137526 392080
rect 131206 391960 131212 392012
rect 131264 392000 131270 392012
rect 159358 392000 159364 392012
rect 131264 391972 159364 392000
rect 131264 391960 131270 391972
rect 159358 391960 159364 391972
rect 159416 391960 159422 392012
rect 176010 391892 176016 391944
rect 176068 391932 176074 391944
rect 186314 391932 186320 391944
rect 176068 391904 186320 391932
rect 176068 391892 176074 391904
rect 186314 391892 186320 391904
rect 186372 391892 186378 391944
rect 413370 391212 413376 391264
rect 413428 391252 413434 391264
rect 437566 391252 437572 391264
rect 413428 391224 437572 391252
rect 413428 391212 413434 391224
rect 437566 391212 437572 391224
rect 437624 391212 437630 391264
rect 131206 390600 131212 390652
rect 131264 390640 131270 390652
rect 134702 390640 134708 390652
rect 131264 390612 134708 390640
rect 131264 390600 131270 390612
rect 134702 390600 134708 390612
rect 134760 390600 134766 390652
rect 131482 390532 131488 390584
rect 131540 390572 131546 390584
rect 152550 390572 152556 390584
rect 131540 390544 152556 390572
rect 131540 390532 131546 390544
rect 152550 390532 152556 390544
rect 152608 390532 152614 390584
rect 411990 390260 411996 390312
rect 412048 390300 412054 390312
rect 413462 390300 413468 390312
rect 412048 390272 413468 390300
rect 412048 390260 412054 390272
rect 413462 390260 413468 390272
rect 413520 390260 413526 390312
rect 131298 389784 131304 389836
rect 131356 389824 131362 389836
rect 165062 389824 165068 389836
rect 131356 389796 165068 389824
rect 131356 389784 131362 389796
rect 165062 389784 165068 389796
rect 165120 389784 165126 389836
rect 131114 389308 131120 389360
rect 131172 389348 131178 389360
rect 134518 389348 134524 389360
rect 131172 389320 134524 389348
rect 131172 389308 131178 389320
rect 134518 389308 134524 389320
rect 134576 389308 134582 389360
rect 131206 389240 131212 389292
rect 131264 389280 131270 389292
rect 134610 389280 134616 389292
rect 131264 389252 134616 389280
rect 131264 389240 131270 389252
rect 134610 389240 134616 389252
rect 134668 389240 134674 389292
rect 131482 389172 131488 389224
rect 131540 389212 131546 389224
rect 177482 389212 177488 389224
rect 131540 389184 177488 389212
rect 131540 389172 131546 389184
rect 177482 389172 177488 389184
rect 177540 389172 177546 389224
rect 435450 389172 435456 389224
rect 435508 389212 435514 389224
rect 437750 389212 437756 389224
rect 435508 389184 437756 389212
rect 435508 389172 435514 389184
rect 437750 389172 437756 389184
rect 437808 389172 437814 389224
rect 166258 389104 166264 389156
rect 166316 389144 166322 389156
rect 186406 389144 186412 389156
rect 166316 389116 186412 389144
rect 166316 389104 166322 389116
rect 186406 389104 186412 389116
rect 186464 389104 186470 389156
rect 170398 389036 170404 389088
rect 170456 389076 170462 389088
rect 186314 389076 186320 389088
rect 170456 389048 186320 389076
rect 170456 389036 170462 389048
rect 186314 389036 186320 389048
rect 186372 389036 186378 389088
rect 131206 387880 131212 387932
rect 131264 387920 131270 387932
rect 133506 387920 133512 387932
rect 131264 387892 133512 387920
rect 131264 387880 131270 387892
rect 133506 387880 133512 387892
rect 133564 387880 133570 387932
rect 131298 387812 131304 387864
rect 131356 387852 131362 387864
rect 157978 387852 157984 387864
rect 131356 387824 157984 387852
rect 131356 387812 131362 387824
rect 157978 387812 157984 387824
rect 158036 387812 158042 387864
rect 131206 386588 131212 386640
rect 131264 386628 131270 386640
rect 133414 386628 133420 386640
rect 131264 386600 133420 386628
rect 131264 386588 131270 386600
rect 133414 386588 133420 386600
rect 133472 386588 133478 386640
rect 131114 386384 131120 386436
rect 131172 386424 131178 386436
rect 184474 386424 184480 386436
rect 131172 386396 184480 386424
rect 131172 386384 131178 386396
rect 184474 386384 184480 386396
rect 184532 386384 184538 386436
rect 155218 386316 155224 386368
rect 155276 386356 155282 386368
rect 186314 386356 186320 386368
rect 155276 386328 186320 386356
rect 155276 386316 155282 386328
rect 186314 386316 186320 386328
rect 186372 386316 186378 386368
rect 417694 385636 417700 385688
rect 417752 385676 417758 385688
rect 437474 385676 437480 385688
rect 417752 385648 437480 385676
rect 417752 385636 417758 385648
rect 437474 385636 437480 385648
rect 437532 385636 437538 385688
rect 131114 385160 131120 385212
rect 131172 385200 131178 385212
rect 141418 385200 141424 385212
rect 131172 385172 141424 385200
rect 131172 385160 131178 385172
rect 141418 385160 141424 385172
rect 141476 385160 141482 385212
rect 131206 385092 131212 385144
rect 131264 385132 131270 385144
rect 155310 385132 155316 385144
rect 131264 385104 155316 385132
rect 131264 385092 131270 385104
rect 155310 385092 155316 385104
rect 155368 385092 155374 385144
rect 131298 385024 131304 385076
rect 131356 385064 131362 385076
rect 156690 385064 156696 385076
rect 131356 385036 156696 385064
rect 131356 385024 131362 385036
rect 156690 385024 156696 385036
rect 156748 385024 156754 385076
rect 131206 383732 131212 383784
rect 131264 383772 131270 383784
rect 147030 383772 147036 383784
rect 131264 383744 147036 383772
rect 131264 383732 131270 383744
rect 147030 383732 147036 383744
rect 147088 383732 147094 383784
rect 430114 383732 430120 383784
rect 430172 383772 430178 383784
rect 437474 383772 437480 383784
rect 430172 383744 437480 383772
rect 430172 383732 430178 383744
rect 437474 383732 437480 383744
rect 437532 383732 437538 383784
rect 131114 383664 131120 383716
rect 131172 383704 131178 383716
rect 182910 383704 182916 383716
rect 131172 383676 182916 383704
rect 131172 383664 131178 383676
rect 182910 383664 182916 383676
rect 182968 383664 182974 383716
rect 411806 383664 411812 383716
rect 411864 383704 411870 383716
rect 438210 383704 438216 383716
rect 411864 383676 438216 383704
rect 411864 383664 411870 383676
rect 438210 383664 438216 383676
rect 438268 383664 438274 383716
rect 131114 382304 131120 382356
rect 131172 382344 131178 382356
rect 133322 382344 133328 382356
rect 131172 382316 133328 382344
rect 131172 382304 131178 382316
rect 133322 382304 133328 382316
rect 133380 382304 133386 382356
rect 131206 382236 131212 382288
rect 131264 382276 131270 382288
rect 176194 382276 176200 382288
rect 131264 382248 176200 382276
rect 131264 382236 131270 382248
rect 176194 382236 176200 382248
rect 176252 382236 176258 382288
rect 435818 382236 435824 382288
rect 435876 382276 435882 382288
rect 437934 382276 437940 382288
rect 435876 382248 437940 382276
rect 435876 382236 435882 382248
rect 437934 382236 437940 382248
rect 437992 382236 437998 382288
rect 132218 381012 132224 381064
rect 132276 381052 132282 381064
rect 138658 381052 138664 381064
rect 132276 381024 138664 381052
rect 132276 381012 132282 381024
rect 138658 381012 138664 381024
rect 138716 381012 138722 381064
rect 131206 380944 131212 380996
rect 131264 380984 131270 380996
rect 180150 380984 180156 380996
rect 131264 380956 180156 380984
rect 131264 380944 131270 380956
rect 180150 380944 180156 380956
rect 180208 380944 180214 380996
rect 131482 380876 131488 380928
rect 131540 380916 131546 380928
rect 184382 380916 184388 380928
rect 131540 380888 184388 380916
rect 131540 380876 131546 380888
rect 184382 380876 184388 380888
rect 184440 380876 184446 380928
rect 411714 380876 411720 380928
rect 411772 380916 411778 380928
rect 416774 380916 416780 380928
rect 411772 380888 416780 380916
rect 411772 380876 411778 380888
rect 416774 380876 416780 380888
rect 416832 380876 416838 380928
rect 428826 380876 428832 380928
rect 428884 380916 428890 380928
rect 437474 380916 437480 380928
rect 428884 380888 437480 380916
rect 428884 380876 428890 380888
rect 437474 380876 437480 380888
rect 437532 380876 437538 380928
rect 144178 380808 144184 380860
rect 144236 380848 144242 380860
rect 186406 380848 186412 380860
rect 144236 380820 186412 380848
rect 144236 380808 144242 380820
rect 186406 380808 186412 380820
rect 186464 380808 186470 380860
rect 131206 379584 131212 379636
rect 131264 379624 131270 379636
rect 151170 379624 151176 379636
rect 131264 379596 151176 379624
rect 131264 379584 131270 379596
rect 151170 379584 151176 379596
rect 151228 379584 151234 379636
rect 131482 379516 131488 379568
rect 131540 379556 131546 379568
rect 173342 379556 173348 379568
rect 131540 379528 173348 379556
rect 131540 379516 131546 379528
rect 173342 379516 173348 379528
rect 173400 379516 173406 379568
rect 413278 379516 413284 379568
rect 413336 379556 413342 379568
rect 437474 379556 437480 379568
rect 413336 379528 437480 379556
rect 413336 379516 413342 379528
rect 437474 379516 437480 379528
rect 437532 379516 437538 379568
rect 142798 379448 142804 379500
rect 142856 379488 142862 379500
rect 186314 379488 186320 379500
rect 142856 379460 186320 379488
rect 142856 379448 142862 379460
rect 186314 379448 186320 379460
rect 186372 379448 186378 379500
rect 131114 378292 131120 378344
rect 131172 378332 131178 378344
rect 142890 378332 142896 378344
rect 131172 378304 142896 378332
rect 131172 378292 131178 378304
rect 142890 378292 142896 378304
rect 142948 378292 142954 378344
rect 131206 378224 131212 378276
rect 131264 378264 131270 378276
rect 146938 378264 146944 378276
rect 131264 378236 146944 378264
rect 131264 378224 131270 378236
rect 146938 378224 146944 378236
rect 146996 378224 147002 378276
rect 131298 378156 131304 378208
rect 131356 378196 131362 378208
rect 178862 378196 178868 378208
rect 131356 378168 178868 378196
rect 131356 378156 131362 378168
rect 178862 378156 178868 378168
rect 178920 378156 178926 378208
rect 554038 378156 554044 378208
rect 554096 378196 554102 378208
rect 580166 378196 580172 378208
rect 554096 378168 580172 378196
rect 554096 378156 554102 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 131942 378088 131948 378140
rect 132000 378128 132006 378140
rect 186314 378128 186320 378140
rect 132000 378100 186320 378128
rect 132000 378088 132006 378100
rect 186314 378088 186320 378100
rect 186372 378088 186378 378140
rect 131206 376796 131212 376848
rect 131264 376836 131270 376848
rect 137370 376836 137376 376848
rect 131264 376808 137376 376836
rect 131264 376796 131270 376808
rect 137370 376796 137376 376808
rect 137428 376796 137434 376848
rect 131114 376728 131120 376780
rect 131172 376768 131178 376780
rect 166258 376768 166264 376780
rect 131172 376740 166264 376768
rect 131172 376728 131178 376740
rect 166258 376728 166264 376740
rect 166316 376728 166322 376780
rect 422938 376728 422944 376780
rect 422996 376768 423002 376780
rect 437474 376768 437480 376780
rect 422996 376740 437480 376768
rect 422996 376728 423002 376740
rect 437474 376728 437480 376740
rect 437532 376728 437538 376780
rect 141510 376660 141516 376712
rect 141568 376700 141574 376712
rect 186314 376700 186320 376712
rect 141568 376672 186320 376700
rect 141568 376660 141574 376672
rect 186314 376660 186320 376672
rect 186372 376660 186378 376712
rect 131482 375436 131488 375488
rect 131540 375476 131546 375488
rect 144178 375476 144184 375488
rect 131540 375448 144184 375476
rect 131540 375436 131546 375448
rect 144178 375436 144184 375448
rect 144236 375436 144242 375488
rect 131206 375368 131212 375420
rect 131264 375408 131270 375420
rect 181622 375408 181628 375420
rect 131264 375380 181628 375408
rect 131264 375368 131270 375380
rect 181622 375368 181628 375380
rect 181680 375368 181686 375420
rect 421926 375368 421932 375420
rect 421984 375408 421990 375420
rect 437474 375408 437480 375420
rect 421984 375380 437480 375408
rect 421984 375368 421990 375380
rect 437474 375368 437480 375380
rect 437532 375368 437538 375420
rect 140222 375300 140228 375352
rect 140280 375340 140286 375352
rect 186314 375340 186320 375352
rect 140280 375312 186320 375340
rect 140280 375300 140286 375312
rect 186314 375300 186320 375312
rect 186372 375300 186378 375352
rect 183002 375232 183008 375284
rect 183060 375272 183066 375284
rect 186406 375272 186412 375284
rect 183060 375244 186412 375272
rect 183060 375232 183066 375244
rect 186406 375232 186412 375244
rect 186464 375232 186470 375284
rect 432966 374280 432972 374332
rect 433024 374320 433030 374332
rect 437474 374320 437480 374332
rect 433024 374292 437480 374320
rect 433024 374280 433030 374292
rect 437474 374280 437480 374292
rect 437532 374280 437538 374332
rect 131206 374144 131212 374196
rect 131264 374184 131270 374196
rect 140130 374184 140136 374196
rect 131264 374156 140136 374184
rect 131264 374144 131270 374156
rect 140130 374144 140136 374156
rect 140188 374144 140194 374196
rect 131114 374076 131120 374128
rect 131172 374116 131178 374128
rect 140038 374116 140044 374128
rect 131172 374088 140044 374116
rect 131172 374076 131178 374088
rect 140038 374076 140044 374088
rect 140096 374076 140102 374128
rect 131206 374008 131212 374060
rect 131264 374048 131270 374060
rect 156598 374048 156604 374060
rect 131264 374020 156604 374048
rect 131264 374008 131270 374020
rect 156598 374008 156604 374020
rect 156656 374008 156662 374060
rect 162210 373940 162216 373992
rect 162268 373980 162274 373992
rect 186314 373980 186320 373992
rect 162268 373952 186320 373980
rect 162268 373940 162274 373952
rect 186314 373940 186320 373952
rect 186372 373940 186378 373992
rect 131206 372648 131212 372700
rect 131264 372688 131270 372700
rect 142798 372688 142804 372700
rect 131264 372660 142804 372688
rect 131264 372648 131270 372660
rect 142798 372648 142804 372660
rect 142856 372648 142862 372700
rect 131482 372580 131488 372632
rect 131540 372620 131546 372632
rect 170398 372620 170404 372632
rect 131540 372592 170404 372620
rect 131540 372580 131546 372592
rect 170398 372580 170404 372592
rect 170456 372580 170462 372632
rect 174538 372512 174544 372564
rect 174596 372552 174602 372564
rect 186314 372552 186320 372564
rect 174596 372524 186320 372552
rect 174596 372512 174602 372524
rect 186314 372512 186320 372524
rect 186372 372512 186378 372564
rect 131206 371288 131212 371340
rect 131264 371328 131270 371340
rect 137278 371328 137284 371340
rect 131264 371300 137284 371328
rect 131264 371288 131270 371300
rect 137278 371288 137284 371300
rect 137336 371288 137342 371340
rect 426066 371288 426072 371340
rect 426124 371328 426130 371340
rect 437474 371328 437480 371340
rect 426124 371300 437480 371328
rect 426124 371288 426130 371300
rect 437474 371288 437480 371300
rect 437532 371288 437538 371340
rect 131114 371220 131120 371272
rect 131172 371260 131178 371272
rect 164970 371260 164976 371272
rect 131172 371232 164976 371260
rect 131172 371220 131178 371232
rect 164970 371220 164976 371232
rect 165028 371220 165034 371272
rect 411254 371220 411260 371272
rect 411312 371260 411318 371272
rect 439682 371260 439688 371272
rect 411312 371232 439688 371260
rect 411312 371220 411318 371232
rect 439682 371220 439688 371232
rect 439740 371220 439746 371272
rect 160738 371152 160744 371204
rect 160796 371192 160802 371204
rect 186314 371192 186320 371204
rect 160796 371164 186320 371192
rect 160796 371152 160802 371164
rect 186314 371152 186320 371164
rect 186372 371152 186378 371204
rect 181530 371084 181536 371136
rect 181588 371124 181594 371136
rect 186406 371124 186412 371136
rect 181588 371096 186412 371124
rect 181588 371084 181594 371096
rect 186406 371084 186412 371096
rect 186464 371084 186470 371136
rect 131206 369928 131212 369980
rect 131264 369968 131270 369980
rect 162118 369968 162124 369980
rect 131264 369940 162124 369968
rect 131264 369928 131270 369940
rect 162118 369928 162124 369940
rect 162176 369928 162182 369980
rect 131114 369860 131120 369912
rect 131172 369900 131178 369912
rect 177390 369900 177396 369912
rect 131172 369872 177396 369900
rect 131172 369860 131178 369872
rect 177390 369860 177396 369872
rect 177448 369860 177454 369912
rect 424594 369860 424600 369912
rect 424652 369900 424658 369912
rect 437474 369900 437480 369912
rect 424652 369872 437480 369900
rect 424652 369860 424658 369872
rect 437474 369860 437480 369872
rect 437532 369860 437538 369912
rect 159358 369792 159364 369844
rect 159416 369832 159422 369844
rect 186314 369832 186320 369844
rect 159416 369804 186320 369832
rect 159416 369792 159422 369804
rect 186314 369792 186320 369804
rect 186372 369792 186378 369844
rect 131482 368568 131488 368620
rect 131540 368608 131546 368620
rect 152458 368608 152464 368620
rect 131540 368580 152464 368608
rect 131540 368568 131546 368580
rect 152458 368568 152464 368580
rect 152516 368568 152522 368620
rect 131206 368500 131212 368552
rect 131264 368540 131270 368552
rect 174538 368540 174544 368552
rect 131264 368512 174544 368540
rect 131264 368500 131270 368512
rect 174538 368500 174544 368512
rect 174596 368500 174602 368552
rect 137462 368432 137468 368484
rect 137520 368472 137526 368484
rect 186314 368472 186320 368484
rect 137520 368444 186320 368472
rect 137520 368432 137526 368444
rect 186314 368432 186320 368444
rect 186372 368432 186378 368484
rect 131206 367208 131212 367260
rect 131264 367248 131270 367260
rect 135898 367248 135904 367260
rect 131264 367220 135904 367248
rect 131264 367208 131270 367220
rect 135898 367208 135904 367220
rect 135956 367208 135962 367260
rect 131114 367140 131120 367192
rect 131172 367180 131178 367192
rect 160738 367180 160744 367192
rect 131172 367152 160744 367180
rect 131172 367140 131178 367152
rect 160738 367140 160744 367152
rect 160796 367140 160802 367192
rect 131206 367072 131212 367124
rect 131264 367112 131270 367124
rect 176010 367112 176016 367124
rect 131264 367084 176016 367112
rect 131264 367072 131270 367084
rect 176010 367072 176016 367084
rect 176068 367072 176074 367124
rect 431586 367072 431592 367124
rect 431644 367112 431650 367124
rect 437474 367112 437480 367124
rect 431644 367084 437480 367112
rect 431644 367072 431650 367084
rect 437474 367072 437480 367084
rect 437532 367072 437538 367124
rect 134702 367004 134708 367056
rect 134760 367044 134766 367056
rect 186406 367044 186412 367056
rect 134760 367016 186412 367044
rect 134760 367004 134766 367016
rect 186406 367004 186412 367016
rect 186464 367004 186470 367056
rect 165062 366936 165068 366988
rect 165120 366976 165126 366988
rect 186314 366976 186320 366988
rect 165120 366948 186320 366976
rect 165120 366936 165126 366948
rect 186314 366936 186320 366948
rect 186372 366936 186378 366988
rect 131206 365712 131212 365764
rect 131264 365752 131270 365764
rect 163682 365752 163688 365764
rect 131264 365724 163688 365752
rect 131264 365712 131270 365724
rect 163682 365712 163688 365724
rect 163740 365712 163746 365764
rect 432874 365712 432880 365764
rect 432932 365752 432938 365764
rect 437474 365752 437480 365764
rect 432932 365724 437480 365752
rect 432932 365712 432938 365724
rect 437474 365712 437480 365724
rect 437532 365712 437538 365764
rect 152550 365644 152556 365696
rect 152608 365684 152614 365696
rect 186314 365684 186320 365696
rect 152608 365656 186320 365684
rect 152608 365644 152614 365656
rect 186314 365644 186320 365656
rect 186372 365644 186378 365696
rect 433978 364556 433984 364608
rect 434036 364596 434042 364608
rect 437474 364596 437480 364608
rect 434036 364568 437480 364596
rect 434036 364556 434042 364568
rect 437474 364556 437480 364568
rect 437532 364556 437538 364608
rect 131114 364420 131120 364472
rect 131172 364460 131178 364472
rect 169110 364460 169116 364472
rect 131172 364432 169116 364460
rect 131172 364420 131178 364432
rect 169110 364420 169116 364432
rect 169168 364420 169174 364472
rect 131206 364352 131212 364404
rect 131264 364392 131270 364404
rect 181530 364392 181536 364404
rect 131264 364364 181536 364392
rect 131264 364352 131270 364364
rect 181530 364352 181536 364364
rect 181588 364352 181594 364404
rect 558178 364352 558184 364404
rect 558236 364392 558242 364404
rect 580166 364392 580172 364404
rect 558236 364364 580172 364392
rect 558236 364352 558242 364364
rect 580166 364352 580172 364364
rect 580224 364352 580230 364404
rect 134518 364284 134524 364336
rect 134576 364324 134582 364336
rect 186314 364324 186320 364336
rect 134576 364296 186320 364324
rect 134576 364284 134582 364296
rect 186314 364284 186320 364296
rect 186372 364284 186378 364336
rect 131114 363060 131120 363112
rect 131172 363100 131178 363112
rect 133230 363100 133236 363112
rect 131172 363072 133236 363100
rect 131172 363060 131178 363072
rect 133230 363060 133236 363072
rect 133288 363060 133294 363112
rect 131206 362992 131212 363044
rect 131264 363032 131270 363044
rect 152734 363032 152740 363044
rect 131264 363004 152740 363032
rect 131264 362992 131270 363004
rect 152734 362992 152740 363004
rect 152792 362992 152798 363044
rect 131482 362924 131488 362976
rect 131540 362964 131546 362976
rect 159358 362964 159364 362976
rect 131540 362936 159364 362964
rect 131540 362924 131546 362936
rect 159358 362924 159364 362936
rect 159416 362924 159422 362976
rect 415302 362924 415308 362976
rect 415360 362964 415366 362976
rect 437474 362964 437480 362976
rect 415360 362936 437480 362964
rect 415360 362924 415366 362936
rect 437474 362924 437480 362936
rect 437532 362924 437538 362976
rect 177482 362856 177488 362908
rect 177540 362896 177546 362908
rect 186314 362896 186320 362908
rect 177540 362868 186320 362896
rect 177540 362856 177546 362868
rect 186314 362856 186320 362868
rect 186372 362856 186378 362908
rect 132218 362176 132224 362228
rect 132276 362216 132282 362228
rect 173250 362216 173256 362228
rect 132276 362188 173256 362216
rect 132276 362176 132282 362188
rect 173250 362176 173256 362188
rect 173308 362176 173314 362228
rect 131206 361632 131212 361684
rect 131264 361672 131270 361684
rect 148502 361672 148508 361684
rect 131264 361644 148508 361672
rect 131264 361632 131270 361644
rect 148502 361632 148508 361644
rect 148560 361632 148566 361684
rect 131114 361564 131120 361616
rect 131172 361604 131178 361616
rect 178770 361604 178776 361616
rect 131172 361576 178776 361604
rect 131172 361564 131178 361576
rect 178770 361564 178776 361576
rect 178828 361564 178834 361616
rect 134610 361496 134616 361548
rect 134668 361536 134674 361548
rect 186314 361536 186320 361548
rect 134668 361508 186320 361536
rect 134668 361496 134674 361508
rect 186314 361496 186320 361508
rect 186372 361496 186378 361548
rect 157978 361428 157984 361480
rect 158036 361468 158042 361480
rect 186406 361468 186412 361480
rect 158036 361440 186412 361468
rect 158036 361428 158042 361440
rect 186406 361428 186412 361440
rect 186464 361428 186470 361480
rect 131114 360272 131120 360324
rect 131172 360312 131178 360324
rect 134518 360312 134524 360324
rect 131172 360284 134524 360312
rect 131172 360272 131178 360284
rect 134518 360272 134524 360284
rect 134576 360272 134582 360324
rect 131206 360204 131212 360256
rect 131264 360244 131270 360256
rect 158254 360244 158260 360256
rect 131264 360216 158260 360244
rect 131264 360204 131270 360216
rect 158254 360204 158260 360216
rect 158312 360204 158318 360256
rect 414842 360204 414848 360256
rect 414900 360244 414906 360256
rect 437474 360244 437480 360256
rect 414900 360216 437480 360244
rect 414900 360204 414906 360216
rect 437474 360204 437480 360216
rect 437532 360204 437538 360256
rect 133506 360136 133512 360188
rect 133564 360176 133570 360188
rect 186314 360176 186320 360188
rect 133564 360148 186320 360176
rect 133564 360136 133570 360148
rect 186314 360136 186320 360148
rect 186372 360136 186378 360188
rect 411254 359320 411260 359372
rect 411312 359360 411318 359372
rect 412910 359360 412916 359372
rect 411312 359332 412916 359360
rect 411312 359320 411318 359332
rect 412910 359320 412916 359332
rect 412968 359320 412974 359372
rect 132034 358844 132040 358896
rect 132092 358884 132098 358896
rect 165154 358884 165160 358896
rect 132092 358856 165160 358884
rect 132092 358844 132098 358856
rect 165154 358844 165160 358856
rect 165212 358844 165218 358896
rect 131206 358776 131212 358828
rect 131264 358816 131270 358828
rect 177574 358816 177580 358828
rect 131264 358788 177580 358816
rect 131264 358776 131270 358788
rect 177574 358776 177580 358788
rect 177632 358776 177638 358828
rect 184474 358708 184480 358760
rect 184532 358748 184538 358760
rect 187418 358748 187424 358760
rect 184532 358720 187424 358748
rect 184532 358708 184538 358720
rect 187418 358708 187424 358720
rect 187476 358708 187482 358760
rect 131114 357484 131120 357536
rect 131172 357524 131178 357536
rect 166442 357524 166448 357536
rect 131172 357496 166448 357524
rect 131172 357484 131178 357496
rect 166442 357484 166448 357496
rect 166500 357484 166506 357536
rect 131206 357416 131212 357468
rect 131264 357456 131270 357468
rect 183094 357456 183100 357468
rect 131264 357428 183100 357456
rect 131264 357416 131270 357428
rect 183094 357416 183100 357428
rect 183152 357416 183158 357468
rect 414750 357416 414756 357468
rect 414808 357456 414814 357468
rect 437474 357456 437480 357468
rect 414808 357428 437480 357456
rect 414808 357416 414814 357428
rect 437474 357416 437480 357428
rect 437532 357416 437538 357468
rect 133414 357348 133420 357400
rect 133472 357388 133478 357400
rect 186314 357388 186320 357400
rect 133472 357360 186320 357388
rect 133472 357348 133478 357360
rect 186314 357348 186320 357360
rect 186372 357348 186378 357400
rect 156690 357280 156696 357332
rect 156748 357320 156754 357332
rect 186406 357320 186412 357332
rect 156748 357292 186412 357320
rect 156748 357280 156754 357292
rect 186406 357280 186412 357292
rect 186464 357280 186470 357332
rect 131206 356192 131212 356244
rect 131264 356232 131270 356244
rect 138842 356232 138848 356244
rect 131264 356204 138848 356232
rect 131264 356192 131270 356204
rect 138842 356192 138848 356204
rect 138900 356192 138906 356244
rect 131114 356124 131120 356176
rect 131172 356164 131178 356176
rect 145742 356164 145748 356176
rect 131172 356136 145748 356164
rect 131172 356124 131178 356136
rect 145742 356124 145748 356136
rect 145800 356124 145806 356176
rect 131298 356056 131304 356108
rect 131356 356096 131362 356108
rect 158162 356096 158168 356108
rect 131356 356068 158168 356096
rect 131356 356056 131362 356068
rect 158162 356056 158168 356068
rect 158220 356056 158226 356108
rect 428734 356056 428740 356108
rect 428792 356096 428798 356108
rect 437474 356096 437480 356108
rect 428792 356068 437480 356096
rect 428792 356056 428798 356068
rect 437474 356056 437480 356068
rect 437532 356056 437538 356108
rect 141418 355988 141424 356040
rect 141476 356028 141482 356040
rect 186314 356028 186320 356040
rect 141476 356000 186320 356028
rect 141476 355988 141482 356000
rect 186314 355988 186320 356000
rect 186372 355988 186378 356040
rect 131206 354764 131212 354816
rect 131264 354804 131270 354816
rect 141510 354804 141516 354816
rect 131264 354776 141516 354804
rect 131264 354764 131270 354776
rect 141510 354764 141516 354776
rect 141568 354764 141574 354816
rect 131298 354696 131304 354748
rect 131356 354736 131362 354748
rect 156782 354736 156788 354748
rect 131356 354708 156788 354736
rect 131356 354696 131362 354708
rect 156782 354696 156788 354708
rect 156840 354696 156846 354748
rect 427078 354696 427084 354748
rect 427136 354736 427142 354748
rect 437474 354736 437480 354748
rect 427136 354708 437480 354736
rect 427136 354696 427142 354708
rect 437474 354696 437480 354708
rect 437532 354696 437538 354748
rect 155310 354628 155316 354680
rect 155368 354668 155374 354680
rect 186314 354668 186320 354680
rect 155368 354640 186320 354668
rect 155368 354628 155374 354640
rect 186314 354628 186320 354640
rect 186372 354628 186378 354680
rect 131206 353336 131212 353388
rect 131264 353376 131270 353388
rect 155494 353376 155500 353388
rect 131264 353348 155500 353376
rect 131264 353336 131270 353348
rect 155494 353336 155500 353348
rect 155552 353336 155558 353388
rect 131114 353268 131120 353320
rect 131172 353308 131178 353320
rect 184566 353308 184572 353320
rect 131172 353280 184572 353308
rect 131172 353268 131178 353280
rect 184566 353268 184572 353280
rect 184624 353268 184630 353320
rect 424502 353268 424508 353320
rect 424560 353308 424566 353320
rect 437474 353308 437480 353320
rect 424560 353280 437480 353308
rect 424560 353268 424566 353280
rect 437474 353268 437480 353280
rect 437532 353268 437538 353320
rect 147030 353200 147036 353252
rect 147088 353240 147094 353252
rect 186314 353240 186320 353252
rect 147088 353212 186320 353240
rect 147088 353200 147094 353212
rect 186314 353200 186320 353212
rect 186372 353200 186378 353252
rect 182910 353132 182916 353184
rect 182968 353172 182974 353184
rect 186406 353172 186412 353184
rect 182968 353144 186412 353172
rect 182968 353132 182974 353144
rect 186406 353132 186412 353144
rect 186464 353132 186470 353184
rect 411254 353132 411260 353184
rect 411312 353172 411318 353184
rect 413370 353172 413376 353184
rect 411312 353144 413376 353172
rect 411312 353132 411318 353144
rect 413370 353132 413376 353144
rect 413428 353132 413434 353184
rect 131206 352044 131212 352096
rect 131264 352084 131270 352096
rect 141694 352084 141700 352096
rect 131264 352056 141700 352084
rect 131264 352044 131270 352056
rect 141694 352044 141700 352056
rect 141752 352044 141758 352096
rect 131114 351976 131120 352028
rect 131172 352016 131178 352028
rect 144454 352016 144460 352028
rect 131172 351988 144460 352016
rect 131172 351976 131178 351988
rect 144454 351976 144460 351988
rect 144512 351976 144518 352028
rect 131482 351908 131488 351960
rect 131540 351948 131546 351960
rect 148410 351948 148416 351960
rect 131540 351920 148416 351948
rect 131540 351908 131546 351920
rect 148410 351908 148416 351920
rect 148468 351908 148474 351960
rect 133322 351840 133328 351892
rect 133380 351880 133386 351892
rect 186314 351880 186320 351892
rect 133380 351852 186320 351880
rect 133380 351840 133386 351852
rect 186314 351840 186320 351852
rect 186372 351840 186378 351892
rect 131114 350616 131120 350668
rect 131172 350656 131178 350668
rect 141602 350656 141608 350668
rect 131172 350628 141608 350656
rect 131172 350616 131178 350628
rect 141602 350616 141608 350628
rect 141660 350616 141666 350668
rect 131206 350548 131212 350600
rect 131264 350588 131270 350600
rect 176102 350588 176108 350600
rect 131264 350560 176108 350588
rect 131264 350548 131270 350560
rect 176102 350548 176108 350560
rect 176160 350548 176166 350600
rect 420362 350548 420368 350600
rect 420420 350588 420426 350600
rect 437474 350588 437480 350600
rect 420420 350560 437480 350588
rect 420420 350548 420426 350560
rect 437474 350548 437480 350560
rect 437532 350548 437538 350600
rect 176194 350480 176200 350532
rect 176252 350520 176258 350532
rect 186314 350520 186320 350532
rect 176252 350492 186320 350520
rect 176252 350480 176258 350492
rect 186314 350480 186320 350492
rect 186372 350480 186378 350532
rect 131206 349188 131212 349240
rect 131264 349228 131270 349240
rect 147214 349228 147220 349240
rect 131264 349200 147220 349228
rect 131264 349188 131270 349200
rect 147214 349188 147220 349200
rect 147272 349188 147278 349240
rect 131114 349120 131120 349172
rect 131172 349160 131178 349172
rect 174722 349160 174728 349172
rect 131172 349132 174728 349160
rect 131172 349120 131178 349132
rect 174722 349120 174728 349132
rect 174780 349120 174786 349172
rect 435634 349120 435640 349172
rect 435692 349160 435698 349172
rect 437474 349160 437480 349172
rect 435692 349132 437480 349160
rect 435692 349120 435698 349132
rect 437474 349120 437480 349132
rect 437532 349120 437538 349172
rect 138658 349052 138664 349104
rect 138716 349092 138722 349104
rect 186314 349092 186320 349104
rect 138716 349064 186320 349092
rect 138716 349052 138722 349064
rect 186314 349052 186320 349064
rect 186372 349052 186378 349104
rect 184382 348984 184388 349036
rect 184440 349024 184446 349036
rect 186406 349024 186412 349036
rect 184440 348996 186412 349024
rect 184440 348984 184446 348996
rect 186406 348984 186412 348996
rect 186464 348984 186470 349036
rect 131206 348304 131212 348356
rect 131264 348344 131270 348356
rect 134886 348344 134892 348356
rect 131264 348316 134892 348344
rect 131264 348304 131270 348316
rect 134886 348304 134892 348316
rect 134944 348304 134950 348356
rect 131482 347828 131488 347880
rect 131540 347868 131546 347880
rect 134794 347868 134800 347880
rect 131540 347840 134800 347868
rect 131540 347828 131546 347840
rect 134794 347828 134800 347840
rect 134852 347828 134858 347880
rect 131298 347760 131304 347812
rect 131356 347800 131362 347812
rect 145650 347800 145656 347812
rect 131356 347772 145656 347800
rect 131356 347760 131362 347772
rect 145650 347760 145656 347772
rect 145708 347760 145714 347812
rect 423122 347760 423128 347812
rect 423180 347800 423186 347812
rect 437474 347800 437480 347812
rect 423180 347772 437480 347800
rect 423180 347760 423186 347772
rect 437474 347760 437480 347772
rect 437532 347760 437538 347812
rect 180150 347692 180156 347744
rect 180208 347732 180214 347744
rect 186314 347732 186320 347744
rect 180208 347704 186320 347732
rect 180208 347692 180214 347704
rect 186314 347692 186320 347704
rect 186372 347692 186378 347744
rect 131206 346468 131212 346520
rect 131264 346508 131270 346520
rect 162302 346508 162308 346520
rect 131264 346480 162308 346508
rect 131264 346468 131270 346480
rect 162302 346468 162308 346480
rect 162360 346468 162366 346520
rect 131114 346400 131120 346452
rect 131172 346440 131178 346452
rect 180242 346440 180248 346452
rect 131172 346412 180248 346440
rect 131172 346400 131178 346412
rect 180242 346400 180248 346412
rect 180300 346400 180306 346452
rect 430022 346400 430028 346452
rect 430080 346440 430086 346452
rect 437474 346440 437480 346452
rect 430080 346412 437480 346440
rect 430080 346400 430086 346412
rect 437474 346400 437480 346412
rect 437532 346400 437538 346452
rect 151170 346332 151176 346384
rect 151228 346372 151234 346384
rect 186314 346372 186320 346384
rect 151228 346344 186320 346372
rect 151228 346332 151234 346344
rect 186314 346332 186320 346344
rect 186372 346332 186378 346384
rect 131206 345176 131212 345228
rect 131264 345216 131270 345228
rect 143074 345216 143080 345228
rect 131264 345188 143080 345216
rect 131264 345176 131270 345188
rect 143074 345176 143080 345188
rect 143132 345176 143138 345228
rect 131114 345108 131120 345160
rect 131172 345148 131178 345160
rect 155402 345148 155408 345160
rect 131172 345120 155408 345148
rect 131172 345108 131178 345120
rect 155402 345108 155408 345120
rect 155460 345108 155466 345160
rect 131206 345040 131212 345092
rect 131264 345080 131270 345092
rect 170582 345080 170588 345092
rect 131264 345052 170588 345080
rect 131264 345040 131270 345052
rect 170582 345040 170588 345052
rect 170640 345040 170646 345092
rect 429930 345040 429936 345092
rect 429988 345080 429994 345092
rect 437474 345080 437480 345092
rect 429988 345052 437480 345080
rect 429988 345040 429994 345052
rect 437474 345040 437480 345052
rect 437532 345040 437538 345092
rect 173342 344972 173348 345024
rect 173400 345012 173406 345024
rect 186314 345012 186320 345024
rect 173400 344984 186320 345012
rect 173400 344972 173406 344984
rect 186314 344972 186320 344984
rect 186372 344972 186378 345024
rect 131298 343680 131304 343732
rect 131356 343720 131362 343732
rect 153838 343720 153844 343732
rect 131356 343692 153844 343720
rect 131356 343680 131362 343692
rect 153838 343680 153844 343692
rect 153896 343680 153902 343732
rect 411254 343680 411260 343732
rect 411312 343720 411318 343732
rect 413002 343720 413008 343732
rect 411312 343692 413008 343720
rect 411312 343680 411318 343692
rect 413002 343680 413008 343692
rect 413060 343680 413066 343732
rect 131206 343612 131212 343664
rect 131264 343652 131270 343664
rect 173434 343652 173440 343664
rect 131264 343624 173440 343652
rect 131264 343612 131270 343624
rect 173434 343612 173440 343624
rect 173492 343612 173498 343664
rect 142890 343544 142896 343596
rect 142948 343584 142954 343596
rect 186314 343584 186320 343596
rect 142948 343556 186320 343584
rect 142948 343544 142954 343556
rect 186314 343544 186320 343556
rect 186372 343544 186378 343596
rect 178862 343476 178868 343528
rect 178920 343516 178926 343528
rect 186406 343516 186412 343528
rect 178920 343488 186412 343516
rect 178920 343476 178926 343488
rect 186406 343476 186412 343488
rect 186464 343476 186470 343528
rect 131206 342320 131212 342372
rect 131264 342360 131270 342372
rect 144362 342360 144368 342372
rect 131264 342332 144368 342360
rect 131264 342320 131270 342332
rect 144362 342320 144368 342332
rect 144420 342320 144426 342372
rect 423030 342320 423036 342372
rect 423088 342360 423094 342372
rect 437474 342360 437480 342372
rect 423088 342332 437480 342360
rect 423088 342320 423094 342332
rect 437474 342320 437480 342332
rect 437532 342320 437538 342372
rect 131482 342252 131488 342304
rect 131540 342292 131546 342304
rect 159542 342292 159548 342304
rect 131540 342264 159548 342292
rect 131540 342252 131546 342264
rect 159542 342252 159548 342264
rect 159600 342252 159606 342304
rect 411254 342252 411260 342304
rect 411312 342292 411318 342304
rect 439774 342292 439780 342304
rect 411312 342264 439780 342292
rect 411312 342252 411318 342264
rect 439774 342252 439780 342264
rect 439832 342252 439838 342304
rect 146938 342184 146944 342236
rect 146996 342224 147002 342236
rect 186314 342224 186320 342236
rect 146996 342196 186320 342224
rect 146996 342184 147002 342196
rect 186314 342184 186320 342196
rect 186372 342184 186378 342236
rect 131206 341028 131212 341080
rect 131264 341068 131270 341080
rect 149698 341068 149704 341080
rect 131264 341040 149704 341068
rect 131264 341028 131270 341040
rect 149698 341028 149704 341040
rect 149756 341028 149762 341080
rect 131298 340960 131304 341012
rect 131356 341000 131362 341012
rect 160922 341000 160928 341012
rect 131356 340972 160928 341000
rect 131356 340960 131362 340972
rect 160922 340960 160928 340972
rect 160980 340960 160986 341012
rect 131114 340892 131120 340944
rect 131172 340932 131178 340944
rect 178862 340932 178868 340944
rect 131172 340904 178868 340932
rect 131172 340892 131178 340904
rect 178862 340892 178868 340904
rect 178920 340892 178926 340944
rect 166258 340824 166264 340876
rect 166316 340864 166322 340876
rect 186314 340864 186320 340876
rect 166316 340836 186320 340864
rect 166316 340824 166322 340836
rect 186314 340824 186320 340836
rect 186372 340824 186378 340876
rect 132034 340144 132040 340196
rect 132092 340184 132098 340196
rect 180334 340184 180340 340196
rect 132092 340156 180340 340184
rect 132092 340144 132098 340156
rect 180334 340144 180340 340156
rect 180392 340144 180398 340196
rect 131298 339532 131304 339584
rect 131356 339572 131362 339584
rect 137554 339572 137560 339584
rect 131356 339544 137560 339572
rect 131356 339532 131362 339544
rect 137554 339532 137560 339544
rect 137612 339532 137618 339584
rect 131206 339464 131212 339516
rect 131264 339504 131270 339516
rect 166350 339504 166356 339516
rect 131264 339476 166356 339504
rect 131264 339464 131270 339476
rect 166350 339464 166356 339476
rect 166408 339464 166414 339516
rect 435542 339464 435548 339516
rect 435600 339504 435606 339516
rect 437842 339504 437848 339516
rect 435600 339476 437848 339504
rect 435600 339464 435606 339476
rect 437842 339464 437848 339476
rect 437900 339464 437906 339516
rect 137370 339396 137376 339448
rect 137428 339436 137434 339448
rect 186314 339436 186320 339448
rect 137428 339408 186320 339436
rect 137428 339396 137434 339408
rect 186314 339396 186320 339408
rect 186372 339396 186378 339448
rect 181622 339328 181628 339380
rect 181680 339368 181686 339380
rect 186406 339368 186412 339380
rect 181680 339340 186412 339368
rect 181680 339328 181686 339340
rect 186406 339328 186412 339340
rect 186464 339328 186470 339380
rect 131206 338172 131212 338224
rect 131264 338212 131270 338224
rect 137462 338212 137468 338224
rect 131264 338184 137468 338212
rect 131264 338172 131270 338184
rect 137462 338172 137468 338184
rect 137520 338172 137526 338224
rect 131114 338104 131120 338156
rect 131172 338144 131178 338156
rect 152642 338144 152648 338156
rect 131172 338116 152648 338144
rect 131172 338104 131178 338116
rect 152642 338104 152648 338116
rect 152700 338104 152706 338156
rect 417602 338104 417608 338156
rect 417660 338144 417666 338156
rect 437474 338144 437480 338156
rect 417660 338116 437480 338144
rect 417660 338104 417666 338116
rect 437474 338104 437480 338116
rect 437532 338104 437538 338156
rect 144178 338036 144184 338088
rect 144236 338076 144242 338088
rect 186314 338076 186320 338088
rect 144236 338048 186320 338076
rect 144236 338036 144242 338048
rect 186314 338036 186320 338048
rect 186372 338036 186378 338088
rect 411254 338036 411260 338088
rect 411312 338076 411318 338088
rect 417694 338076 417700 338088
rect 411312 338048 417700 338076
rect 411312 338036 411318 338048
rect 417694 338036 417700 338048
rect 417752 338036 417758 338088
rect 131206 336880 131212 336932
rect 131264 336920 131270 336932
rect 147030 336920 147036 336932
rect 131264 336892 147036 336920
rect 131264 336880 131270 336892
rect 147030 336880 147036 336892
rect 147088 336880 147094 336932
rect 132034 336812 132040 336864
rect 132092 336852 132098 336864
rect 151262 336852 151268 336864
rect 132092 336824 151268 336852
rect 132092 336812 132098 336824
rect 151262 336812 151268 336824
rect 151320 336812 151326 336864
rect 131482 336744 131488 336796
rect 131540 336784 131546 336796
rect 181622 336784 181628 336796
rect 131540 336756 181628 336784
rect 131540 336744 131546 336756
rect 181622 336744 181628 336756
rect 181680 336744 181686 336796
rect 425974 336744 425980 336796
rect 426032 336784 426038 336796
rect 437474 336784 437480 336796
rect 426032 336756 437480 336784
rect 426032 336744 426038 336756
rect 437474 336744 437480 336756
rect 437532 336744 437538 336796
rect 140130 336676 140136 336728
rect 140188 336716 140194 336728
rect 186314 336716 186320 336728
rect 140188 336688 186320 336716
rect 140188 336676 140194 336688
rect 186314 336676 186320 336688
rect 186372 336676 186378 336728
rect 131206 335384 131212 335436
rect 131264 335424 131270 335436
rect 140222 335424 140228 335436
rect 131264 335396 140228 335424
rect 131264 335384 131270 335396
rect 140222 335384 140228 335396
rect 140280 335384 140286 335436
rect 131114 335316 131120 335368
rect 131172 335356 131178 335368
rect 147122 335356 147128 335368
rect 131172 335328 147128 335356
rect 131172 335316 131178 335328
rect 147122 335316 147128 335328
rect 147180 335316 147186 335368
rect 140038 335248 140044 335300
rect 140096 335288 140102 335300
rect 186314 335288 186320 335300
rect 140096 335260 186320 335288
rect 140096 335248 140102 335260
rect 186314 335248 186320 335260
rect 186372 335248 186378 335300
rect 156598 335180 156604 335232
rect 156656 335220 156662 335232
rect 186406 335220 186412 335232
rect 156656 335192 186412 335220
rect 156656 335180 156662 335192
rect 186406 335180 186412 335192
rect 186464 335180 186470 335232
rect 132218 334024 132224 334076
rect 132276 334064 132282 334076
rect 142982 334064 142988 334076
rect 132276 334036 142988 334064
rect 132276 334024 132282 334036
rect 142982 334024 142988 334036
rect 143040 334024 143046 334076
rect 131206 333956 131212 334008
rect 131264 333996 131270 334008
rect 163590 333996 163596 334008
rect 131264 333968 163596 333996
rect 131264 333956 131270 333968
rect 163590 333956 163596 333968
rect 163648 333956 163654 334008
rect 142798 333888 142804 333940
rect 142856 333928 142862 333940
rect 186314 333928 186320 333940
rect 142856 333900 186320 333928
rect 142856 333888 142862 333900
rect 186314 333888 186320 333900
rect 186372 333888 186378 333940
rect 131114 332732 131120 332784
rect 131172 332772 131178 332784
rect 140130 332772 140136 332784
rect 131172 332744 140136 332772
rect 131172 332732 131178 332744
rect 140130 332732 140136 332744
rect 140188 332732 140194 332784
rect 131298 332664 131304 332716
rect 131356 332704 131362 332716
rect 142890 332704 142896 332716
rect 131356 332676 142896 332704
rect 131356 332664 131362 332676
rect 142890 332664 142896 332676
rect 142948 332664 142954 332716
rect 131206 332596 131212 332648
rect 131264 332636 131270 332648
rect 183002 332636 183008 332648
rect 131264 332608 183008 332636
rect 131264 332596 131270 332608
rect 183002 332596 183008 332608
rect 183060 332596 183066 332648
rect 419166 332596 419172 332648
rect 419224 332636 419230 332648
rect 437474 332636 437480 332648
rect 419224 332608 437480 332636
rect 419224 332596 419230 332608
rect 437474 332596 437480 332608
rect 437532 332596 437538 332648
rect 170398 332528 170404 332580
rect 170456 332568 170462 332580
rect 186314 332568 186320 332580
rect 170456 332540 186320 332568
rect 170456 332528 170462 332540
rect 186314 332528 186320 332540
rect 186372 332528 186378 332580
rect 132218 331304 132224 331356
rect 132276 331344 132282 331356
rect 140038 331344 140044 331356
rect 132276 331316 140044 331344
rect 132276 331304 132282 331316
rect 140038 331304 140044 331316
rect 140096 331304 140102 331356
rect 131482 331236 131488 331288
rect 131540 331276 131546 331288
rect 170490 331276 170496 331288
rect 131540 331248 170496 331276
rect 131540 331236 131546 331248
rect 170490 331236 170496 331248
rect 170548 331236 170554 331288
rect 416222 331236 416228 331288
rect 416280 331276 416286 331288
rect 437474 331276 437480 331288
rect 416280 331248 437480 331276
rect 416280 331236 416286 331248
rect 437474 331236 437480 331248
rect 437532 331236 437538 331288
rect 137278 331168 137284 331220
rect 137336 331208 137342 331220
rect 186406 331208 186412 331220
rect 137336 331180 186412 331208
rect 137336 331168 137342 331180
rect 186406 331168 186412 331180
rect 186464 331168 186470 331220
rect 164970 331100 164976 331152
rect 165028 331140 165034 331152
rect 186314 331140 186320 331152
rect 165028 331112 186320 331140
rect 165028 331100 165034 331112
rect 186314 331100 186320 331112
rect 186372 331100 186378 331152
rect 417694 330488 417700 330540
rect 417752 330528 417758 330540
rect 437566 330528 437572 330540
rect 417752 330500 437572 330528
rect 417752 330488 417758 330500
rect 437566 330488 437572 330500
rect 437624 330488 437630 330540
rect 132218 329944 132224 329996
rect 132276 329984 132282 329996
rect 133506 329984 133512 329996
rect 132276 329956 133512 329984
rect 132276 329944 132282 329956
rect 133506 329944 133512 329956
rect 133564 329944 133570 329996
rect 131114 329876 131120 329928
rect 131172 329916 131178 329928
rect 159450 329916 159456 329928
rect 131172 329888 159456 329916
rect 131172 329876 131178 329888
rect 159450 329876 159456 329888
rect 159508 329876 159514 329928
rect 431494 329876 431500 329928
rect 431552 329916 431558 329928
rect 437474 329916 437480 329928
rect 431552 329888 437480 329916
rect 431552 329876 431558 329888
rect 437474 329876 437480 329888
rect 437532 329876 437538 329928
rect 131206 329808 131212 329860
rect 131264 329848 131270 329860
rect 165062 329848 165068 329860
rect 131264 329820 165068 329848
rect 131264 329808 131270 329820
rect 165062 329808 165068 329820
rect 165120 329808 165126 329860
rect 411254 329808 411260 329860
rect 411312 329848 411318 329860
rect 439590 329848 439596 329860
rect 411312 329820 439596 329848
rect 411312 329808 411318 329820
rect 439590 329808 439596 329820
rect 439648 329808 439654 329860
rect 131942 329740 131948 329792
rect 132000 329780 132006 329792
rect 186314 329780 186320 329792
rect 132000 329752 186320 329780
rect 132000 329740 132006 329752
rect 186314 329740 186320 329752
rect 186372 329740 186378 329792
rect 131206 328516 131212 328568
rect 131264 328556 131270 328568
rect 152550 328556 152556 328568
rect 131264 328528 152556 328556
rect 131264 328516 131270 328528
rect 152550 328516 152556 328528
rect 152608 328516 152614 328568
rect 131298 328448 131304 328500
rect 131356 328488 131362 328500
rect 174630 328488 174636 328500
rect 131356 328460 174636 328488
rect 131356 328448 131362 328460
rect 174630 328448 174636 328460
rect 174688 328448 174694 328500
rect 421834 328448 421840 328500
rect 421892 328488 421898 328500
rect 437474 328488 437480 328500
rect 421892 328460 437480 328488
rect 421892 328448 421898 328460
rect 437474 328448 437480 328460
rect 437532 328448 437538 328500
rect 177390 328380 177396 328432
rect 177448 328420 177454 328432
rect 186314 328420 186320 328432
rect 177448 328392 186320 328420
rect 177448 328380 177454 328392
rect 186314 328380 186320 328392
rect 186372 328380 186378 328432
rect 131114 327156 131120 327208
rect 131172 327196 131178 327208
rect 166258 327196 166264 327208
rect 131172 327168 166264 327196
rect 131172 327156 131178 327168
rect 166258 327156 166264 327168
rect 166316 327156 166322 327208
rect 131206 327088 131212 327140
rect 131264 327128 131270 327140
rect 184474 327128 184480 327140
rect 131264 327100 184480 327128
rect 131264 327088 131270 327100
rect 184474 327088 184480 327100
rect 184532 327088 184538 327140
rect 162118 327020 162124 327072
rect 162176 327060 162182 327072
rect 186314 327060 186320 327072
rect 162176 327032 186320 327060
rect 162176 327020 162182 327032
rect 186314 327020 186320 327032
rect 186372 327020 186378 327072
rect 174538 326952 174544 327004
rect 174596 326992 174602 327004
rect 186406 326992 186412 327004
rect 174596 326964 186412 326992
rect 174596 326952 174602 326964
rect 186406 326952 186412 326964
rect 186464 326952 186470 327004
rect 427170 326340 427176 326392
rect 427228 326380 427234 326392
rect 438486 326380 438492 326392
rect 427228 326352 438492 326380
rect 427228 326340 427234 326352
rect 438486 326340 438492 326352
rect 438544 326340 438550 326392
rect 132218 325796 132224 325848
rect 132276 325836 132282 325848
rect 160830 325836 160836 325848
rect 132276 325808 160836 325836
rect 132276 325796 132282 325808
rect 160830 325796 160836 325808
rect 160888 325796 160894 325848
rect 131206 325728 131212 325780
rect 131264 325768 131270 325780
rect 158070 325768 158076 325780
rect 131264 325740 158076 325768
rect 131264 325728 131270 325740
rect 158070 325728 158076 325740
rect 158128 325728 158134 325780
rect 131298 325660 131304 325712
rect 131356 325700 131362 325712
rect 133414 325700 133420 325712
rect 131356 325672 133420 325700
rect 131356 325660 131362 325672
rect 133414 325660 133420 325672
rect 133472 325660 133478 325712
rect 411254 325660 411260 325712
rect 411312 325700 411318 325712
rect 431218 325700 431224 325712
rect 411312 325672 431224 325700
rect 411312 325660 411318 325672
rect 431218 325660 431224 325672
rect 431276 325660 431282 325712
rect 152458 325592 152464 325644
rect 152516 325632 152522 325644
rect 186314 325632 186320 325644
rect 152516 325604 186320 325632
rect 152516 325592 152522 325604
rect 186314 325592 186320 325604
rect 186372 325592 186378 325644
rect 131482 324368 131488 324420
rect 131540 324408 131546 324420
rect 151170 324408 151176 324420
rect 131540 324380 151176 324408
rect 131540 324368 131546 324380
rect 151170 324368 151176 324380
rect 151228 324368 151234 324420
rect 131206 324300 131212 324352
rect 131264 324340 131270 324352
rect 169018 324340 169024 324352
rect 131264 324312 169024 324340
rect 131264 324300 131270 324312
rect 169018 324300 169024 324312
rect 169076 324300 169082 324352
rect 411254 324300 411260 324352
rect 411312 324340 411318 324352
rect 439866 324340 439872 324352
rect 411312 324312 439872 324340
rect 411312 324300 411318 324312
rect 439866 324300 439872 324312
rect 439924 324300 439930 324352
rect 551370 324300 551376 324352
rect 551428 324340 551434 324352
rect 580166 324340 580172 324352
rect 551428 324312 580172 324340
rect 551428 324300 551434 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 135898 324232 135904 324284
rect 135956 324272 135962 324284
rect 186314 324272 186320 324284
rect 135956 324244 186320 324272
rect 135956 324232 135962 324244
rect 186314 324232 186320 324244
rect 186372 324232 186378 324284
rect 131482 323076 131488 323128
rect 131540 323116 131546 323128
rect 137370 323116 137376 323128
rect 131540 323088 137376 323116
rect 131540 323076 131546 323088
rect 137370 323076 137376 323088
rect 137428 323076 137434 323128
rect 131114 323008 131120 323060
rect 131172 323048 131178 323060
rect 156690 323048 156696 323060
rect 131172 323020 156696 323048
rect 131172 323008 131178 323020
rect 156690 323008 156696 323020
rect 156748 323008 156754 323060
rect 131206 322940 131212 322992
rect 131264 322980 131270 322992
rect 177482 322980 177488 322992
rect 131264 322952 177488 322980
rect 131264 322940 131270 322952
rect 177482 322940 177488 322952
rect 177540 322940 177546 322992
rect 160738 322872 160744 322924
rect 160796 322912 160802 322924
rect 186314 322912 186320 322924
rect 160796 322884 186320 322912
rect 160796 322872 160802 322884
rect 186314 322872 186320 322884
rect 186372 322872 186378 322924
rect 176010 322804 176016 322856
rect 176068 322844 176074 322856
rect 186406 322844 186412 322856
rect 176068 322816 186412 322844
rect 176068 322804 176074 322816
rect 186406 322804 186412 322816
rect 186464 322804 186470 322856
rect 417786 322192 417792 322244
rect 417844 322232 417850 322244
rect 438394 322232 438400 322244
rect 417844 322204 438400 322232
rect 417844 322192 417850 322204
rect 438394 322192 438400 322204
rect 438452 322192 438458 322244
rect 131206 321648 131212 321700
rect 131264 321688 131270 321700
rect 144270 321688 144276 321700
rect 131264 321660 144276 321688
rect 131264 321648 131270 321660
rect 144270 321648 144276 321660
rect 144328 321648 144334 321700
rect 131114 321580 131120 321632
rect 131172 321620 131178 321632
rect 155310 321620 155316 321632
rect 131172 321592 155316 321620
rect 131172 321580 131178 321592
rect 155310 321580 155316 321592
rect 155368 321580 155374 321632
rect 173250 321512 173256 321564
rect 173308 321552 173314 321564
rect 186314 321552 186320 321564
rect 173308 321524 186320 321552
rect 173308 321512 173314 321524
rect 186314 321512 186320 321524
rect 186372 321512 186378 321564
rect 420270 320832 420276 320884
rect 420328 320872 420334 320884
rect 437474 320872 437480 320884
rect 420328 320844 437480 320872
rect 420328 320832 420334 320844
rect 437474 320832 437480 320844
rect 437532 320832 437538 320884
rect 131114 320220 131120 320272
rect 131172 320260 131178 320272
rect 162210 320260 162216 320272
rect 131172 320232 162216 320260
rect 131172 320220 131178 320232
rect 162210 320220 162216 320232
rect 162268 320220 162274 320272
rect 131206 320152 131212 320204
rect 131264 320192 131270 320204
rect 176010 320192 176016 320204
rect 131264 320164 176016 320192
rect 131264 320152 131270 320164
rect 176010 320152 176016 320164
rect 176068 320152 176074 320204
rect 163682 320084 163688 320136
rect 163740 320124 163746 320136
rect 186314 320124 186320 320136
rect 163740 320096 186320 320124
rect 163740 320084 163746 320096
rect 186314 320084 186320 320096
rect 186372 320084 186378 320136
rect 132218 318860 132224 318912
rect 132276 318900 132282 318912
rect 156598 318900 156604 318912
rect 132276 318872 156604 318900
rect 132276 318860 132282 318872
rect 156598 318860 156604 318872
rect 156656 318860 156662 318912
rect 131206 318792 131212 318844
rect 131264 318832 131270 318844
rect 173250 318832 173256 318844
rect 131264 318804 173256 318832
rect 131264 318792 131270 318804
rect 173250 318792 173256 318804
rect 173308 318792 173314 318844
rect 429838 318792 429844 318844
rect 429896 318832 429902 318844
rect 437474 318832 437480 318844
rect 429896 318804 437480 318832
rect 429896 318792 429902 318804
rect 437474 318792 437480 318804
rect 437532 318792 437538 318844
rect 169110 318724 169116 318776
rect 169168 318764 169174 318776
rect 186314 318764 186320 318776
rect 169168 318736 186320 318764
rect 169168 318724 169174 318736
rect 186314 318724 186320 318736
rect 186372 318724 186378 318776
rect 131482 317432 131488 317484
rect 131540 317472 131546 317484
rect 174538 317472 174544 317484
rect 131540 317444 174544 317472
rect 131540 317432 131546 317444
rect 174538 317432 174544 317444
rect 174596 317432 174602 317484
rect 411254 317432 411260 317484
rect 411312 317472 411318 317484
rect 425790 317472 425796 317484
rect 411312 317444 425796 317472
rect 411312 317432 411318 317444
rect 425790 317432 425796 317444
rect 425848 317432 425854 317484
rect 159358 317364 159364 317416
rect 159416 317404 159422 317416
rect 186314 317404 186320 317416
rect 159416 317376 186320 317404
rect 159416 317364 159422 317376
rect 186314 317364 186320 317376
rect 186372 317364 186378 317416
rect 431954 317364 431960 317416
rect 432012 317404 432018 317416
rect 438302 317404 438308 317416
rect 432012 317376 438308 317404
rect 432012 317364 432018 317376
rect 438302 317364 438308 317376
rect 438360 317364 438366 317416
rect 181530 317296 181536 317348
rect 181588 317336 181594 317348
rect 186406 317336 186412 317348
rect 181588 317308 186412 317336
rect 181588 317296 181594 317308
rect 186406 317296 186412 317308
rect 186464 317296 186470 317348
rect 132218 316072 132224 316124
rect 132276 316112 132282 316124
rect 133322 316112 133328 316124
rect 132276 316084 133328 316112
rect 132276 316072 132282 316084
rect 133322 316072 133328 316084
rect 133380 316072 133386 316124
rect 131206 316004 131212 316056
rect 131264 316044 131270 316056
rect 155218 316044 155224 316056
rect 131264 316016 155224 316044
rect 131264 316004 131270 316016
rect 155218 316004 155224 316016
rect 155276 316004 155282 316056
rect 411254 316004 411260 316056
rect 411312 316044 411318 316056
rect 428458 316044 428464 316056
rect 411312 316016 428464 316044
rect 411312 316004 411318 316016
rect 428458 316004 428464 316016
rect 428516 316004 428522 316056
rect 133230 315936 133236 315988
rect 133288 315976 133294 315988
rect 186314 315976 186320 315988
rect 133288 315948 186320 315976
rect 133288 315936 133294 315948
rect 186314 315936 186320 315948
rect 186372 315936 186378 315988
rect 131482 314712 131488 314764
rect 131540 314752 131546 314764
rect 138750 314752 138756 314764
rect 131540 314724 138756 314752
rect 131540 314712 131546 314724
rect 138750 314712 138756 314724
rect 138808 314712 138814 314764
rect 131206 314644 131212 314696
rect 131264 314684 131270 314696
rect 180150 314684 180156 314696
rect 131264 314656 180156 314684
rect 131264 314644 131270 314656
rect 180150 314644 180156 314656
rect 180208 314644 180214 314696
rect 419074 314644 419080 314696
rect 419132 314684 419138 314696
rect 437474 314684 437480 314696
rect 419132 314656 437480 314684
rect 419132 314644 419138 314656
rect 437474 314644 437480 314656
rect 437532 314644 437538 314696
rect 152734 314576 152740 314628
rect 152792 314616 152798 314628
rect 186314 314616 186320 314628
rect 152792 314588 186320 314616
rect 152792 314576 152798 314588
rect 186314 314576 186320 314588
rect 186372 314576 186378 314628
rect 131298 313896 131304 313948
rect 131356 313936 131362 313948
rect 170398 313936 170404 313948
rect 131356 313908 170404 313936
rect 131356 313896 131362 313908
rect 170398 313896 170404 313908
rect 170456 313896 170462 313948
rect 131206 313352 131212 313404
rect 131264 313392 131270 313404
rect 152458 313392 152464 313404
rect 131264 313364 152464 313392
rect 131264 313352 131270 313364
rect 152458 313352 152464 313364
rect 152516 313352 152522 313404
rect 131114 313284 131120 313336
rect 131172 313324 131178 313336
rect 157978 313324 157984 313336
rect 131172 313296 157984 313324
rect 131172 313284 131178 313296
rect 157978 313284 157984 313296
rect 158036 313284 158042 313336
rect 411254 313284 411260 313336
rect 411312 313324 411318 313336
rect 421558 313324 421564 313336
rect 411312 313296 421564 313324
rect 411312 313284 411318 313296
rect 421558 313284 421564 313296
rect 421616 313284 421622 313336
rect 421742 313284 421748 313336
rect 421800 313324 421806 313336
rect 437474 313324 437480 313336
rect 421800 313296 437480 313324
rect 421800 313284 421806 313296
rect 437474 313284 437480 313296
rect 437532 313284 437538 313336
rect 148502 313216 148508 313268
rect 148560 313256 148566 313268
rect 186406 313256 186412 313268
rect 148560 313228 186412 313256
rect 148560 313216 148566 313228
rect 186406 313216 186412 313228
rect 186464 313216 186470 313268
rect 178770 313148 178776 313200
rect 178828 313188 178834 313200
rect 186314 313188 186320 313200
rect 178828 313160 186320 313188
rect 178828 313148 178834 313160
rect 186314 313148 186320 313160
rect 186372 313148 186378 313200
rect 131114 311924 131120 311976
rect 131172 311964 131178 311976
rect 148318 311964 148324 311976
rect 131172 311936 148324 311964
rect 131172 311924 131178 311936
rect 148318 311924 148324 311936
rect 148376 311924 148382 311976
rect 131206 311856 131212 311908
rect 131264 311896 131270 311908
rect 164970 311896 164976 311908
rect 131264 311868 164976 311896
rect 131264 311856 131270 311868
rect 164970 311856 164976 311868
rect 165028 311856 165034 311908
rect 411254 311856 411260 311908
rect 411312 311896 411318 311908
rect 424318 311896 424324 311908
rect 411312 311868 424324 311896
rect 411312 311856 411318 311868
rect 424318 311856 424324 311868
rect 424376 311856 424382 311908
rect 434070 311856 434076 311908
rect 434128 311896 434134 311908
rect 438762 311896 438768 311908
rect 434128 311868 438768 311896
rect 434128 311856 434134 311868
rect 438762 311856 438768 311868
rect 438820 311856 438826 311908
rect 556798 311856 556804 311908
rect 556856 311896 556862 311908
rect 580166 311896 580172 311908
rect 556856 311868 580172 311896
rect 556856 311856 556862 311868
rect 580166 311856 580172 311868
rect 580224 311856 580230 311908
rect 134518 311788 134524 311840
rect 134576 311828 134582 311840
rect 186314 311828 186320 311840
rect 134576 311800 186320 311828
rect 134576 311788 134582 311800
rect 186314 311788 186320 311800
rect 186372 311788 186378 311840
rect 131482 310564 131488 310616
rect 131540 310604 131546 310616
rect 159358 310604 159364 310616
rect 131540 310576 159364 310604
rect 131540 310564 131546 310576
rect 159358 310564 159364 310576
rect 159416 310564 159422 310616
rect 131206 310496 131212 310548
rect 131264 310536 131270 310548
rect 182910 310536 182916 310548
rect 131264 310508 182916 310536
rect 131264 310496 131270 310508
rect 182910 310496 182916 310508
rect 182968 310496 182974 310548
rect 414658 310496 414664 310548
rect 414716 310536 414722 310548
rect 437474 310536 437480 310548
rect 414716 310508 437480 310536
rect 414716 310496 414722 310508
rect 437474 310496 437480 310508
rect 437532 310496 437538 310548
rect 180334 310428 180340 310480
rect 180392 310468 180398 310480
rect 186314 310468 186320 310480
rect 180392 310440 186320 310468
rect 180392 310428 180398 310440
rect 186314 310428 186320 310440
rect 186372 310428 186378 310480
rect 131298 309748 131304 309800
rect 131356 309788 131362 309800
rect 184382 309788 184388 309800
rect 131356 309760 184388 309788
rect 131356 309748 131362 309760
rect 184382 309748 184388 309760
rect 184440 309748 184446 309800
rect 420914 309748 420920 309800
rect 420972 309788 420978 309800
rect 431954 309788 431960 309800
rect 420972 309760 431960 309788
rect 420972 309748 420978 309760
rect 431954 309748 431960 309760
rect 432012 309748 432018 309800
rect 131114 309612 131120 309664
rect 131172 309652 131178 309664
rect 134702 309652 134708 309664
rect 131172 309624 134708 309652
rect 131172 309612 131178 309624
rect 134702 309612 134708 309624
rect 134760 309612 134766 309664
rect 131206 309136 131212 309188
rect 131264 309176 131270 309188
rect 141418 309176 141424 309188
rect 131264 309148 141424 309176
rect 131264 309136 131270 309148
rect 141418 309136 141424 309148
rect 141476 309136 141482 309188
rect 411254 309136 411260 309188
rect 411312 309176 411318 309188
rect 420914 309176 420920 309188
rect 411312 309148 420920 309176
rect 411312 309136 411318 309148
rect 420914 309136 420920 309148
rect 420972 309136 420978 309188
rect 158254 309068 158260 309120
rect 158312 309108 158318 309120
rect 186314 309108 186320 309120
rect 158312 309080 186320 309108
rect 158312 309068 158318 309080
rect 186314 309068 186320 309080
rect 186372 309068 186378 309120
rect 410518 309068 410524 309120
rect 410576 309108 410582 309120
rect 417786 309108 417792 309120
rect 410576 309080 417792 309108
rect 410576 309068 410582 309080
rect 417786 309068 417792 309080
rect 417844 309068 417850 309120
rect 165154 309000 165160 309052
rect 165212 309040 165218 309052
rect 186406 309040 186412 309052
rect 165212 309012 186412 309040
rect 165212 309000 165218 309012
rect 186406 309000 186412 309012
rect 186464 309000 186470 309052
rect 131206 307912 131212 307964
rect 131264 307952 131270 307964
rect 134610 307952 134616 307964
rect 131264 307924 134616 307952
rect 131264 307912 131270 307924
rect 134610 307912 134616 307924
rect 134668 307912 134674 307964
rect 131114 307844 131120 307896
rect 131172 307884 131178 307896
rect 145558 307884 145564 307896
rect 131172 307856 145564 307884
rect 131172 307844 131178 307856
rect 145558 307844 145564 307856
rect 145616 307844 145622 307896
rect 131482 307776 131488 307828
rect 131540 307816 131546 307828
rect 160738 307816 160744 307828
rect 131540 307788 160744 307816
rect 131540 307776 131546 307788
rect 160738 307776 160744 307788
rect 160796 307776 160802 307828
rect 432690 307776 432696 307828
rect 432748 307816 432754 307828
rect 437474 307816 437480 307828
rect 432748 307788 437480 307816
rect 432748 307776 432754 307788
rect 437474 307776 437480 307788
rect 437532 307776 437538 307828
rect 177574 307708 177580 307760
rect 177632 307748 177638 307760
rect 186314 307748 186320 307760
rect 177632 307720 186320 307748
rect 177632 307708 177638 307720
rect 186314 307708 186320 307720
rect 186372 307708 186378 307760
rect 424686 307028 424692 307080
rect 424744 307068 424750 307080
rect 438394 307068 438400 307080
rect 424744 307040 438400 307068
rect 424744 307028 424750 307040
rect 438394 307028 438400 307040
rect 438452 307028 438458 307080
rect 131114 306416 131120 306468
rect 131172 306456 131178 306468
rect 142798 306456 142804 306468
rect 131172 306428 142804 306456
rect 131172 306416 131178 306428
rect 142798 306416 142804 306428
rect 142856 306416 142862 306468
rect 131206 306348 131212 306400
rect 131264 306388 131270 306400
rect 177390 306388 177396 306400
rect 131264 306360 177396 306388
rect 131264 306348 131270 306360
rect 177390 306348 177396 306360
rect 177448 306348 177454 306400
rect 166442 306280 166448 306332
rect 166500 306320 166506 306332
rect 186314 306320 186320 306332
rect 166500 306292 186320 306320
rect 166500 306280 166506 306292
rect 186314 306280 186320 306292
rect 186372 306280 186378 306332
rect 409966 306280 409972 306332
rect 410024 306320 410030 306332
rect 430114 306320 430120 306332
rect 410024 306292 430120 306320
rect 410024 306280 410030 306292
rect 430114 306280 430120 306292
rect 430172 306280 430178 306332
rect 131482 305124 131488 305176
rect 131540 305164 131546 305176
rect 178770 305164 178776 305176
rect 131540 305136 178776 305164
rect 131540 305124 131546 305136
rect 178770 305124 178776 305136
rect 178828 305124 178834 305176
rect 131114 305056 131120 305108
rect 131172 305096 131178 305108
rect 137278 305096 137284 305108
rect 131172 305068 137284 305096
rect 131172 305056 131178 305068
rect 137278 305056 137284 305068
rect 137336 305056 137342 305108
rect 131206 304988 131212 305040
rect 131264 305028 131270 305040
rect 133230 305028 133236 305040
rect 131264 305000 133236 305028
rect 131264 304988 131270 305000
rect 133230 304988 133236 305000
rect 133288 304988 133294 305040
rect 428642 304988 428648 305040
rect 428700 305028 428706 305040
rect 437474 305028 437480 305040
rect 428700 305000 437480 305028
rect 428700 304988 428706 305000
rect 437474 304988 437480 305000
rect 437532 304988 437538 305040
rect 158162 304920 158168 304972
rect 158220 304960 158226 304972
rect 186406 304960 186412 304972
rect 158220 304932 186412 304960
rect 158220 304920 158226 304932
rect 186406 304920 186412 304932
rect 186464 304920 186470 304972
rect 183094 304852 183100 304904
rect 183152 304892 183158 304904
rect 186682 304892 186688 304904
rect 183152 304864 186688 304892
rect 183152 304852 183158 304864
rect 186682 304852 186688 304864
rect 186740 304852 186746 304904
rect 421006 304240 421012 304292
rect 421064 304280 421070 304292
rect 435818 304280 435824 304292
rect 421064 304252 435824 304280
rect 421064 304240 421070 304252
rect 435818 304240 435824 304252
rect 435876 304240 435882 304292
rect 131298 303696 131304 303748
rect 131356 303736 131362 303748
rect 144178 303736 144184 303748
rect 131356 303708 144184 303736
rect 131356 303696 131362 303708
rect 144178 303696 144184 303708
rect 144236 303696 144242 303748
rect 131206 303628 131212 303680
rect 131264 303668 131270 303680
rect 181530 303668 181536 303680
rect 131264 303640 181536 303668
rect 131264 303628 131270 303640
rect 181530 303628 181536 303640
rect 181588 303628 181594 303680
rect 411254 303628 411260 303680
rect 411312 303668 411318 303680
rect 421006 303668 421012 303680
rect 411312 303640 421012 303668
rect 411312 303628 411318 303640
rect 421006 303628 421012 303640
rect 421064 303628 421070 303680
rect 435726 303628 435732 303680
rect 435784 303668 435790 303680
rect 438670 303668 438676 303680
rect 435784 303640 438676 303668
rect 435784 303628 435790 303640
rect 438670 303628 438676 303640
rect 438728 303628 438734 303680
rect 145742 303560 145748 303612
rect 145800 303600 145806 303612
rect 186314 303600 186320 303612
rect 145800 303572 186320 303600
rect 145800 303560 145806 303572
rect 186314 303560 186320 303572
rect 186372 303560 186378 303612
rect 131114 302268 131120 302320
rect 131172 302308 131178 302320
rect 135898 302308 135904 302320
rect 131172 302280 135904 302308
rect 131172 302268 131178 302280
rect 135898 302268 135904 302280
rect 135956 302268 135962 302320
rect 131206 302200 131212 302252
rect 131264 302240 131270 302252
rect 162118 302240 162124 302252
rect 131264 302212 162124 302240
rect 131264 302200 131270 302212
rect 162118 302200 162124 302212
rect 162176 302200 162182 302252
rect 432782 302200 432788 302252
rect 432840 302240 432846 302252
rect 438026 302240 438032 302252
rect 432840 302212 438032 302240
rect 432840 302200 432846 302212
rect 438026 302200 438032 302212
rect 438084 302200 438090 302252
rect 138842 302132 138848 302184
rect 138900 302172 138906 302184
rect 186314 302172 186320 302184
rect 138900 302144 186320 302172
rect 138900 302132 138906 302144
rect 186314 302132 186320 302144
rect 186372 302132 186378 302184
rect 411530 302132 411536 302184
rect 411588 302172 411594 302184
rect 428826 302172 428832 302184
rect 411588 302144 428832 302172
rect 411588 302132 411594 302144
rect 428826 302132 428832 302144
rect 428884 302132 428890 302184
rect 431402 301452 431408 301504
rect 431460 301492 431466 301504
rect 437566 301492 437572 301504
rect 431460 301464 437572 301492
rect 431460 301452 431466 301464
rect 437566 301452 437572 301464
rect 437624 301452 437630 301504
rect 131206 300908 131212 300960
rect 131264 300948 131270 300960
rect 138658 300948 138664 300960
rect 131264 300920 138664 300948
rect 131264 300908 131270 300920
rect 138658 300908 138664 300920
rect 138716 300908 138722 300960
rect 131482 300840 131488 300892
rect 131540 300880 131546 300892
rect 146938 300880 146944 300892
rect 131540 300852 146944 300880
rect 131540 300840 131546 300852
rect 146938 300840 146944 300852
rect 146996 300840 147002 300892
rect 156782 300772 156788 300824
rect 156840 300812 156846 300824
rect 186314 300812 186320 300824
rect 156840 300784 186320 300812
rect 156840 300772 156846 300784
rect 186314 300772 186320 300784
rect 186372 300772 186378 300824
rect 410518 300772 410524 300824
rect 410576 300812 410582 300824
rect 413278 300812 413284 300824
rect 410576 300784 413284 300812
rect 410576 300772 410582 300784
rect 413278 300772 413284 300784
rect 413336 300772 413342 300824
rect 439774 300772 439780 300824
rect 439832 300812 439838 300824
rect 552198 300812 552204 300824
rect 439832 300784 552204 300812
rect 439832 300772 439838 300784
rect 552198 300772 552204 300784
rect 552256 300772 552262 300824
rect 439866 300704 439872 300756
rect 439924 300744 439930 300756
rect 550542 300744 550548 300756
rect 439924 300716 550548 300744
rect 439924 300704 439930 300716
rect 550542 300704 550548 300716
rect 550600 300704 550606 300756
rect 428826 300092 428832 300144
rect 428884 300132 428890 300144
rect 438578 300132 438584 300144
rect 428884 300104 438584 300132
rect 428884 300092 428890 300104
rect 438578 300092 438584 300104
rect 438636 300092 438642 300144
rect 131114 299888 131120 299940
rect 131172 299928 131178 299940
rect 134518 299928 134524 299940
rect 131172 299900 134524 299928
rect 131172 299888 131178 299900
rect 134518 299888 134524 299900
rect 134576 299888 134582 299940
rect 141510 299412 141516 299464
rect 141568 299452 141574 299464
rect 186314 299452 186320 299464
rect 141568 299424 186320 299452
rect 141568 299412 141574 299424
rect 186314 299412 186320 299424
rect 186372 299412 186378 299464
rect 184566 299344 184572 299396
rect 184624 299384 184630 299396
rect 186406 299384 186412 299396
rect 184624 299356 186412 299384
rect 184624 299344 184630 299356
rect 186406 299344 186412 299356
rect 186464 299344 186470 299396
rect 522298 298120 522304 298172
rect 522356 298160 522362 298172
rect 580166 298160 580172 298172
rect 522356 298132 580172 298160
rect 522356 298120 522362 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 155494 298052 155500 298104
rect 155552 298092 155558 298104
rect 186314 298092 186320 298104
rect 155552 298064 186320 298092
rect 155552 298052 155558 298064
rect 186314 298052 186320 298064
rect 186372 298052 186378 298104
rect 418982 298052 418988 298104
rect 419040 298092 419046 298104
rect 545482 298092 545488 298104
rect 419040 298064 545488 298092
rect 419040 298052 419046 298064
rect 545482 298052 545488 298064
rect 545540 298052 545546 298104
rect 421650 297984 421656 298036
rect 421708 298024 421714 298036
rect 528738 298024 528744 298036
rect 421708 297996 528744 298024
rect 421708 297984 421714 297996
rect 528738 297984 528744 297996
rect 528796 297984 528802 298036
rect 411254 297916 411260 297968
rect 411312 297956 411318 297968
rect 422938 297956 422944 297968
rect 411312 297928 422944 297956
rect 411312 297916 411318 297928
rect 422938 297916 422944 297928
rect 422996 297916 423002 297968
rect 431310 297916 431316 297968
rect 431368 297956 431374 297968
rect 520274 297956 520280 297968
rect 431368 297928 520280 297956
rect 431368 297916 431374 297928
rect 520274 297916 520280 297928
rect 520332 297916 520338 297968
rect 428550 297848 428556 297900
rect 428608 297888 428614 297900
rect 511994 297888 512000 297900
rect 428608 297860 512000 297888
rect 428608 297848 428614 297860
rect 511994 297848 512000 297860
rect 512052 297848 512058 297900
rect 424410 297780 424416 297832
rect 424468 297820 424474 297832
rect 503162 297820 503168 297832
rect 424468 297792 503168 297820
rect 424468 297780 424474 297792
rect 503162 297780 503168 297792
rect 503220 297780 503226 297832
rect 425882 297712 425888 297764
rect 425940 297752 425946 297764
rect 494698 297752 494704 297764
rect 425940 297724 494704 297752
rect 425940 297712 425946 297724
rect 494698 297712 494704 297724
rect 494756 297712 494762 297764
rect 132126 297372 132132 297424
rect 132184 297412 132190 297424
rect 141510 297412 141516 297424
rect 132184 297384 141516 297412
rect 132184 297372 132190 297384
rect 141510 297372 141516 297384
rect 141568 297372 141574 297424
rect 141694 296624 141700 296676
rect 141752 296664 141758 296676
rect 186314 296664 186320 296676
rect 141752 296636 186320 296664
rect 141752 296624 141758 296636
rect 186314 296624 186320 296636
rect 186372 296624 186378 296676
rect 410150 296624 410156 296676
rect 410208 296664 410214 296676
rect 421926 296664 421932 296676
rect 410208 296636 421932 296664
rect 410208 296624 410214 296636
rect 421926 296624 421932 296636
rect 421984 296624 421990 296676
rect 422938 295944 422944 295996
rect 422996 295984 423002 295996
rect 438394 295984 438400 295996
rect 422996 295956 438400 295984
rect 422996 295944 423002 295956
rect 438394 295944 438400 295956
rect 438452 295944 438458 295996
rect 477494 295944 477500 295996
rect 477552 295984 477558 295996
rect 544378 295984 544384 295996
rect 477552 295956 544384 295984
rect 477552 295944 477558 295956
rect 544378 295944 544384 295956
rect 544436 295944 544442 295996
rect 144454 295264 144460 295316
rect 144512 295304 144518 295316
rect 186314 295304 186320 295316
rect 144512 295276 186320 295304
rect 144512 295264 144518 295276
rect 186314 295264 186320 295276
rect 186372 295264 186378 295316
rect 148410 295196 148416 295248
rect 148468 295236 148474 295248
rect 186406 295236 186412 295248
rect 148468 295208 186412 295236
rect 148468 295196 148474 295208
rect 186406 295196 186412 295208
rect 186464 295196 186470 295248
rect 420178 294652 420184 294704
rect 420236 294692 420242 294704
rect 511994 294692 512000 294704
rect 420236 294664 512000 294692
rect 420236 294652 420242 294664
rect 511994 294652 512000 294664
rect 512052 294652 512058 294704
rect 416130 294584 416136 294636
rect 416188 294624 416194 294636
rect 512178 294624 512184 294636
rect 416188 294596 512184 294624
rect 416188 294584 416194 294596
rect 512178 294584 512184 294596
rect 512236 294584 512242 294636
rect 141602 293904 141608 293956
rect 141660 293944 141666 293956
rect 186314 293944 186320 293956
rect 141660 293916 186320 293944
rect 141660 293904 141666 293916
rect 186314 293904 186320 293916
rect 186372 293904 186378 293956
rect 439682 293904 439688 293956
rect 439740 293944 439746 293956
rect 441614 293944 441620 293956
rect 439740 293916 441620 293944
rect 439740 293904 439746 293916
rect 441614 293904 441620 293916
rect 441672 293904 441678 293956
rect 419626 293224 419632 293276
rect 419684 293264 419690 293276
rect 432966 293264 432972 293276
rect 419684 293236 432972 293264
rect 419684 293224 419690 293236
rect 432966 293224 432972 293236
rect 433024 293224 433030 293276
rect 411254 292544 411260 292596
rect 411312 292584 411318 292596
rect 419626 292584 419632 292596
rect 411312 292556 419632 292584
rect 411312 292544 411318 292556
rect 419626 292544 419632 292556
rect 419684 292544 419690 292596
rect 176102 292476 176108 292528
rect 176160 292516 176166 292528
rect 186314 292516 186320 292528
rect 176160 292488 186320 292516
rect 176160 292476 176166 292488
rect 186314 292476 186320 292488
rect 186372 292476 186378 292528
rect 419626 291864 419632 291916
rect 419684 291904 419690 291916
rect 437014 291904 437020 291916
rect 419684 291876 437020 291904
rect 419684 291864 419690 291876
rect 437014 291864 437020 291876
rect 437072 291864 437078 291916
rect 131942 291796 131948 291848
rect 132000 291836 132006 291848
rect 176194 291836 176200 291848
rect 132000 291808 176200 291836
rect 132000 291796 132006 291808
rect 176194 291796 176200 291808
rect 176252 291796 176258 291848
rect 416038 291796 416044 291848
rect 416096 291836 416102 291848
rect 512086 291836 512092 291848
rect 416096 291808 512092 291836
rect 416096 291796 416102 291808
rect 512086 291796 512092 291808
rect 512144 291796 512150 291848
rect 411254 291184 411260 291236
rect 411312 291224 411318 291236
rect 419626 291224 419632 291236
rect 411312 291196 419632 291224
rect 411312 291184 411318 291196
rect 419626 291184 419632 291196
rect 419684 291184 419690 291236
rect 147214 291116 147220 291168
rect 147272 291156 147278 291168
rect 186406 291156 186412 291168
rect 147272 291128 186412 291156
rect 147272 291116 147278 291128
rect 186406 291116 186412 291128
rect 186464 291116 186470 291168
rect 174722 291048 174728 291100
rect 174780 291088 174786 291100
rect 186314 291088 186320 291100
rect 174780 291060 186320 291088
rect 174780 291048 174786 291060
rect 186314 291048 186320 291060
rect 186372 291048 186378 291100
rect 134886 289756 134892 289808
rect 134944 289796 134950 289808
rect 186314 289796 186320 289808
rect 134944 289768 186320 289796
rect 134944 289756 134950 289768
rect 186314 289756 186320 289768
rect 186372 289756 186378 289808
rect 415394 289076 415400 289128
rect 415452 289116 415458 289128
rect 426066 289116 426072 289128
rect 415452 289088 426072 289116
rect 415452 289076 415458 289088
rect 426066 289076 426072 289088
rect 426124 289076 426130 289128
rect 411254 288396 411260 288448
rect 411312 288436 411318 288448
rect 415394 288436 415400 288448
rect 411312 288408 415400 288436
rect 411312 288396 411318 288408
rect 415394 288396 415400 288408
rect 415452 288396 415458 288448
rect 145650 288328 145656 288380
rect 145708 288368 145714 288380
rect 186314 288368 186320 288380
rect 145708 288340 186320 288368
rect 145708 288328 145714 288340
rect 186314 288328 186320 288340
rect 186372 288328 186378 288380
rect 411254 287036 411260 287088
rect 411312 287076 411318 287088
rect 418154 287076 418160 287088
rect 411312 287048 418160 287076
rect 411312 287036 411318 287048
rect 418154 287036 418160 287048
rect 418212 287076 418218 287088
rect 424594 287076 424600 287088
rect 418212 287048 424600 287076
rect 418212 287036 418218 287048
rect 424594 287036 424600 287048
rect 424652 287036 424658 287088
rect 134794 286968 134800 287020
rect 134852 287008 134858 287020
rect 186314 287008 186320 287020
rect 134852 286980 186320 287008
rect 134852 286968 134858 286980
rect 186314 286968 186320 286980
rect 186372 286968 186378 287020
rect 180242 286900 180248 286952
rect 180300 286940 180306 286952
rect 186406 286940 186412 286952
rect 180300 286912 186412 286940
rect 180300 286900 180306 286912
rect 186406 286900 186412 286912
rect 186464 286900 186470 286952
rect 162302 285608 162308 285660
rect 162360 285648 162366 285660
rect 186314 285648 186320 285660
rect 162360 285620 186320 285648
rect 162360 285608 162366 285620
rect 186314 285608 186320 285620
rect 186372 285608 186378 285660
rect 419810 284928 419816 284980
rect 419868 284968 419874 284980
rect 431586 284968 431592 284980
rect 419868 284940 431592 284968
rect 419868 284928 419874 284940
rect 431586 284928 431592 284940
rect 431644 284928 431650 284980
rect 411254 284316 411260 284368
rect 411312 284356 411318 284368
rect 419810 284356 419816 284368
rect 411312 284328 419816 284356
rect 411312 284316 411318 284328
rect 419810 284316 419816 284328
rect 419868 284316 419874 284368
rect 143074 284248 143080 284300
rect 143132 284288 143138 284300
rect 186314 284288 186320 284300
rect 143132 284260 186320 284288
rect 143132 284248 143138 284260
rect 186314 284248 186320 284260
rect 186372 284248 186378 284300
rect 418246 283636 418252 283688
rect 418304 283676 418310 283688
rect 432874 283676 432880 283688
rect 418304 283648 432880 283676
rect 418304 283636 418310 283648
rect 432874 283636 432880 283648
rect 432932 283636 432938 283688
rect 414934 283568 414940 283620
rect 414992 283608 414998 283620
rect 438486 283608 438492 283620
rect 414992 283580 438492 283608
rect 414992 283568 414998 283580
rect 438486 283568 438492 283580
rect 438544 283568 438550 283620
rect 411254 282888 411260 282940
rect 411312 282928 411318 282940
rect 418246 282928 418252 282940
rect 411312 282900 418252 282928
rect 411312 282888 411318 282900
rect 418246 282888 418252 282900
rect 418304 282888 418310 282940
rect 155402 282820 155408 282872
rect 155460 282860 155466 282872
rect 186314 282860 186320 282872
rect 155460 282832 186320 282860
rect 155460 282820 155466 282832
rect 186314 282820 186320 282832
rect 186372 282820 186378 282872
rect 170582 282752 170588 282804
rect 170640 282792 170646 282804
rect 186406 282792 186412 282804
rect 170640 282764 186412 282792
rect 170640 282752 170646 282764
rect 186406 282752 186412 282764
rect 186464 282752 186470 282804
rect 153838 281460 153844 281512
rect 153896 281500 153902 281512
rect 186314 281500 186320 281512
rect 153896 281472 186320 281500
rect 153896 281460 153902 281472
rect 186314 281460 186320 281472
rect 186372 281460 186378 281512
rect 418338 280780 418344 280832
rect 418396 280820 418402 280832
rect 433978 280820 433984 280832
rect 418396 280792 433984 280820
rect 418396 280780 418402 280792
rect 433978 280780 433984 280792
rect 434036 280780 434042 280832
rect 411254 280168 411260 280220
rect 411312 280208 411318 280220
rect 418338 280208 418344 280220
rect 411312 280180 418344 280208
rect 411312 280168 411318 280180
rect 418338 280168 418344 280180
rect 418396 280168 418402 280220
rect 173434 280100 173440 280152
rect 173492 280140 173498 280152
rect 186314 280140 186320 280152
rect 173492 280112 186320 280140
rect 173492 280100 173498 280112
rect 186314 280100 186320 280112
rect 186372 280100 186378 280152
rect 132034 279420 132040 279472
rect 132092 279460 132098 279472
rect 173342 279460 173348 279472
rect 132092 279432 173348 279460
rect 132092 279420 132098 279432
rect 173342 279420 173348 279432
rect 173400 279420 173406 279472
rect 411254 279420 411260 279472
rect 411312 279460 411318 279472
rect 415302 279460 415308 279472
rect 411312 279432 415308 279460
rect 411312 279420 411318 279432
rect 415302 279420 415308 279432
rect 415360 279460 415366 279472
rect 416866 279460 416872 279472
rect 415360 279432 416872 279460
rect 415360 279420 415366 279432
rect 416866 279420 416872 279432
rect 416924 279420 416930 279472
rect 144362 278672 144368 278724
rect 144420 278712 144426 278724
rect 186314 278712 186320 278724
rect 144420 278684 186320 278712
rect 144420 278672 144426 278684
rect 186314 278672 186320 278684
rect 186372 278672 186378 278724
rect 159542 277312 159548 277364
rect 159600 277352 159606 277364
rect 186314 277352 186320 277364
rect 159600 277324 186320 277352
rect 159600 277312 159606 277324
rect 186314 277312 186320 277324
rect 186372 277312 186378 277364
rect 178862 277244 178868 277296
rect 178920 277284 178926 277296
rect 186406 277284 186412 277296
rect 178920 277256 186412 277284
rect 178920 277244 178926 277256
rect 186406 277244 186412 277256
rect 186464 277244 186470 277296
rect 411254 276836 411260 276888
rect 411312 276876 411318 276888
rect 414014 276876 414020 276888
rect 411312 276848 414020 276876
rect 411312 276836 411318 276848
rect 414014 276836 414020 276848
rect 414072 276876 414078 276888
rect 414842 276876 414848 276888
rect 414072 276848 414848 276876
rect 414072 276836 414078 276848
rect 414842 276836 414848 276848
rect 414900 276836 414906 276888
rect 160922 275952 160928 276004
rect 160980 275992 160986 276004
rect 186314 275992 186320 276004
rect 160980 275964 186320 275992
rect 160980 275952 160986 275964
rect 186314 275952 186320 275964
rect 186372 275952 186378 276004
rect 416682 275272 416688 275324
rect 416740 275312 416746 275324
rect 436922 275312 436928 275324
rect 416740 275284 436928 275312
rect 416740 275272 416746 275284
rect 436922 275272 436928 275284
rect 436980 275272 436986 275324
rect 411254 274660 411260 274712
rect 411312 274700 411318 274712
rect 415486 274700 415492 274712
rect 411312 274672 415492 274700
rect 411312 274660 411318 274672
rect 415486 274660 415492 274672
rect 415544 274700 415550 274712
rect 416682 274700 416688 274712
rect 415544 274672 416688 274700
rect 415544 274660 415550 274672
rect 416682 274660 416688 274672
rect 416740 274660 416746 274712
rect 149698 274592 149704 274644
rect 149756 274632 149762 274644
rect 186314 274632 186320 274644
rect 149756 274604 186320 274632
rect 149756 274592 149762 274604
rect 186314 274592 186320 274604
rect 186372 274592 186378 274644
rect 137554 273164 137560 273216
rect 137612 273204 137618 273216
rect 186314 273204 186320 273216
rect 137612 273176 186320 273204
rect 137612 273164 137618 273176
rect 186314 273164 186320 273176
rect 186372 273164 186378 273216
rect 411254 273164 411260 273216
rect 411312 273204 411318 273216
rect 413094 273204 413100 273216
rect 411312 273176 413100 273204
rect 411312 273164 411318 273176
rect 413094 273164 413100 273176
rect 413152 273204 413158 273216
rect 414750 273204 414756 273216
rect 413152 273176 414756 273204
rect 413152 273164 413158 273176
rect 414750 273164 414756 273176
rect 414808 273164 414814 273216
rect 166350 273096 166356 273148
rect 166408 273136 166414 273148
rect 186406 273136 186412 273148
rect 166408 273108 186412 273136
rect 166408 273096 166414 273108
rect 186406 273096 186412 273108
rect 186464 273096 186470 273148
rect 515398 271872 515404 271924
rect 515456 271912 515462 271924
rect 579798 271912 579804 271924
rect 515456 271884 579804 271912
rect 515456 271872 515462 271884
rect 579798 271872 579804 271884
rect 579856 271872 579862 271924
rect 152642 271804 152648 271856
rect 152700 271844 152706 271856
rect 186314 271844 186320 271856
rect 152700 271816 186320 271844
rect 152700 271804 152706 271816
rect 186314 271804 186320 271816
rect 186372 271804 186378 271856
rect 416682 271124 416688 271176
rect 416740 271164 416746 271176
rect 428734 271164 428740 271176
rect 416740 271136 428740 271164
rect 416740 271124 416746 271136
rect 428734 271124 428740 271136
rect 428792 271124 428798 271176
rect 411254 270512 411260 270564
rect 411312 270552 411318 270564
rect 415578 270552 415584 270564
rect 411312 270524 415584 270552
rect 411312 270512 411318 270524
rect 415578 270512 415584 270524
rect 415636 270552 415642 270564
rect 416682 270552 416688 270564
rect 415636 270524 416688 270552
rect 415636 270512 415642 270524
rect 416682 270512 416688 270524
rect 416740 270512 416746 270564
rect 137462 270444 137468 270496
rect 137520 270484 137526 270496
rect 186314 270484 186320 270496
rect 137520 270456 186320 270484
rect 137520 270444 137526 270456
rect 186314 270444 186320 270456
rect 186372 270444 186378 270496
rect 151262 269016 151268 269068
rect 151320 269056 151326 269068
rect 186314 269056 186320 269068
rect 151320 269028 186320 269056
rect 151320 269016 151326 269028
rect 186314 269016 186320 269028
rect 186372 269016 186378 269068
rect 181622 268948 181628 269000
rect 181680 268988 181686 269000
rect 186406 268988 186412 269000
rect 181680 268960 186412 268988
rect 181680 268948 181686 268960
rect 186406 268948 186412 268960
rect 186464 268948 186470 269000
rect 416958 268336 416964 268388
rect 417016 268376 417022 268388
rect 427078 268376 427084 268388
rect 417016 268348 427084 268376
rect 417016 268336 417022 268348
rect 427078 268336 427084 268348
rect 427136 268336 427142 268388
rect 411254 267724 411260 267776
rect 411312 267764 411318 267776
rect 416958 267764 416964 267776
rect 411312 267736 416964 267764
rect 411312 267724 411318 267736
rect 416958 267724 416964 267736
rect 417016 267724 417022 267776
rect 147030 267656 147036 267708
rect 147088 267696 147094 267708
rect 186314 267696 186320 267708
rect 147088 267668 186320 267696
rect 147088 267656 147094 267668
rect 186314 267656 186320 267668
rect 186372 267656 186378 267708
rect 411254 266976 411260 267028
rect 411312 267016 411318 267028
rect 414106 267016 414112 267028
rect 411312 266988 414112 267016
rect 411312 266976 411318 266988
rect 414106 266976 414112 266988
rect 414164 267016 414170 267028
rect 424502 267016 424508 267028
rect 414164 266988 424508 267016
rect 414164 266976 414170 266988
rect 424502 266976 424508 266988
rect 424560 266976 424566 267028
rect 147122 266296 147128 266348
rect 147180 266336 147186 266348
rect 186314 266336 186320 266348
rect 147180 266308 186320 266336
rect 147180 266296 147186 266308
rect 186314 266296 186320 266308
rect 186372 266296 186378 266348
rect 140222 264868 140228 264920
rect 140280 264908 140286 264920
rect 186314 264908 186320 264920
rect 140280 264880 186320 264908
rect 140280 264868 140286 264880
rect 186314 264868 186320 264880
rect 186372 264868 186378 264920
rect 163590 264800 163596 264852
rect 163648 264840 163654 264852
rect 186406 264840 186412 264852
rect 163648 264812 186412 264840
rect 163648 264800 163654 264812
rect 186406 264800 186412 264812
rect 186464 264800 186470 264852
rect 411254 263576 411260 263628
rect 411312 263616 411318 263628
rect 415670 263616 415676 263628
rect 411312 263588 415676 263616
rect 411312 263576 411318 263588
rect 415670 263576 415676 263588
rect 415728 263616 415734 263628
rect 420362 263616 420368 263628
rect 415728 263588 420368 263616
rect 415728 263576 415734 263588
rect 420362 263576 420368 263588
rect 420420 263576 420426 263628
rect 142982 263508 142988 263560
rect 143040 263548 143046 263560
rect 186314 263548 186320 263560
rect 143040 263520 186320 263548
rect 143040 263508 143046 263520
rect 186314 263508 186320 263520
rect 186372 263508 186378 263560
rect 411254 262828 411260 262880
rect 411312 262868 411318 262880
rect 414198 262868 414204 262880
rect 411312 262840 414204 262868
rect 411312 262828 411318 262840
rect 414198 262828 414204 262840
rect 414256 262868 414262 262880
rect 435634 262868 435640 262880
rect 414256 262840 435640 262868
rect 414256 262828 414262 262840
rect 435634 262828 435640 262840
rect 435692 262828 435698 262880
rect 140130 262148 140136 262200
rect 140188 262188 140194 262200
rect 186314 262188 186320 262200
rect 140188 262160 186320 262188
rect 140188 262148 140194 262160
rect 186314 262148 186320 262160
rect 186372 262148 186378 262200
rect 142890 260788 142896 260840
rect 142948 260828 142954 260840
rect 186314 260828 186320 260840
rect 142948 260800 186320 260828
rect 142948 260788 142954 260800
rect 186314 260788 186320 260800
rect 186372 260788 186378 260840
rect 411254 259428 411260 259480
rect 411312 259468 411318 259480
rect 417050 259468 417056 259480
rect 411312 259440 417056 259468
rect 411312 259428 411318 259440
rect 417050 259428 417056 259440
rect 417108 259468 417114 259480
rect 423122 259468 423128 259480
rect 417108 259440 423128 259468
rect 417108 259428 417114 259440
rect 423122 259428 423128 259440
rect 423180 259428 423186 259480
rect 140038 259360 140044 259412
rect 140096 259400 140102 259412
rect 186314 259400 186320 259412
rect 140096 259372 186320 259400
rect 140096 259360 140102 259372
rect 186314 259360 186320 259372
rect 186372 259360 186378 259412
rect 183002 259292 183008 259344
rect 183060 259332 183066 259344
rect 186406 259332 186412 259344
rect 183060 259304 186412 259332
rect 183060 259292 183066 259304
rect 186406 259292 186412 259304
rect 186464 259292 186470 259344
rect 411254 258680 411260 258732
rect 411312 258720 411318 258732
rect 414290 258720 414296 258732
rect 411312 258692 414296 258720
rect 411312 258680 411318 258692
rect 414290 258680 414296 258692
rect 414348 258720 414354 258732
rect 430022 258720 430028 258732
rect 414348 258692 430028 258720
rect 414348 258680 414354 258692
rect 430022 258680 430028 258692
rect 430080 258680 430086 258732
rect 555418 258068 555424 258120
rect 555476 258108 555482 258120
rect 580166 258108 580172 258120
rect 555476 258080 580172 258108
rect 555476 258068 555482 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 170490 258000 170496 258052
rect 170548 258040 170554 258052
rect 186314 258040 186320 258052
rect 170548 258012 186320 258040
rect 170548 258000 170554 258012
rect 186314 258000 186320 258012
rect 186372 258000 186378 258052
rect 159450 256640 159456 256692
rect 159508 256680 159514 256692
rect 186314 256680 186320 256692
rect 159508 256652 186320 256680
rect 159508 256640 159514 256652
rect 186314 256640 186320 256652
rect 186372 256640 186378 256692
rect 417326 255960 417332 256012
rect 417384 256000 417390 256012
rect 429930 256000 429936 256012
rect 417384 255972 429936 256000
rect 417384 255960 417390 255972
rect 429930 255960 429936 255972
rect 429988 255960 429994 256012
rect 430022 255960 430028 256012
rect 430080 256000 430086 256012
rect 438302 256000 438308 256012
rect 430080 255972 438308 256000
rect 430080 255960 430086 255972
rect 438302 255960 438308 255972
rect 438360 255960 438366 256012
rect 411254 255280 411260 255332
rect 411312 255320 411318 255332
rect 417142 255320 417148 255332
rect 411312 255292 417148 255320
rect 411312 255280 411318 255292
rect 417142 255280 417148 255292
rect 417200 255320 417206 255332
rect 417326 255320 417332 255332
rect 417200 255292 417332 255320
rect 417200 255280 417206 255292
rect 417326 255280 417332 255292
rect 417384 255280 417390 255332
rect 133506 255212 133512 255264
rect 133564 255252 133570 255264
rect 186314 255252 186320 255264
rect 133564 255224 186320 255252
rect 133564 255212 133570 255224
rect 186314 255212 186320 255224
rect 186372 255212 186378 255264
rect 165062 255144 165068 255196
rect 165120 255184 165126 255196
rect 186406 255184 186412 255196
rect 165120 255156 186412 255184
rect 165120 255144 165126 255156
rect 186406 255144 186412 255156
rect 186464 255144 186470 255196
rect 411254 254532 411260 254584
rect 411312 254572 411318 254584
rect 414382 254572 414388 254584
rect 411312 254544 414388 254572
rect 411312 254532 411318 254544
rect 414382 254532 414388 254544
rect 414440 254572 414446 254584
rect 423030 254572 423036 254584
rect 414440 254544 423036 254572
rect 414440 254532 414446 254544
rect 423030 254532 423036 254544
rect 423088 254532 423094 254584
rect 152550 253852 152556 253904
rect 152608 253892 152614 253904
rect 186314 253892 186320 253904
rect 152608 253864 186320 253892
rect 152608 253852 152614 253864
rect 186314 253852 186320 253864
rect 186372 253852 186378 253904
rect 174630 252492 174636 252544
rect 174688 252532 174694 252544
rect 186314 252532 186320 252544
rect 174688 252504 186320 252532
rect 174688 252492 174694 252504
rect 186314 252492 186320 252504
rect 186372 252492 186378 252544
rect 410794 252492 410800 252544
rect 410852 252532 410858 252544
rect 427170 252532 427176 252544
rect 410852 252504 427176 252532
rect 410852 252492 410858 252504
rect 427170 252492 427176 252504
rect 427228 252492 427234 252544
rect 166258 251132 166264 251184
rect 166316 251172 166322 251184
rect 186314 251172 186320 251184
rect 166316 251144 186320 251172
rect 166316 251132 166322 251144
rect 186314 251132 186320 251144
rect 186372 251132 186378 251184
rect 184474 251064 184480 251116
rect 184532 251104 184538 251116
rect 186406 251104 186412 251116
rect 184532 251076 186412 251104
rect 184532 251064 184538 251076
rect 186406 251064 186412 251076
rect 186464 251064 186470 251116
rect 411254 250452 411260 250504
rect 411312 250492 411318 250504
rect 411622 250492 411628 250504
rect 411312 250464 411628 250492
rect 411312 250452 411318 250464
rect 411622 250452 411628 250464
rect 411680 250492 411686 250504
rect 435542 250492 435548 250504
rect 411680 250464 435548 250492
rect 411680 250452 411686 250464
rect 435542 250452 435548 250464
rect 435600 250452 435606 250504
rect 160830 249704 160836 249756
rect 160888 249744 160894 249756
rect 186314 249744 186320 249756
rect 160888 249716 186320 249744
rect 160888 249704 160894 249716
rect 186314 249704 186320 249716
rect 186372 249704 186378 249756
rect 133414 248344 133420 248396
rect 133472 248384 133478 248396
rect 186314 248384 186320 248396
rect 133472 248356 186320 248384
rect 133472 248344 133478 248356
rect 186314 248344 186320 248356
rect 186372 248344 186378 248396
rect 411806 247664 411812 247716
rect 411864 247704 411870 247716
rect 417602 247704 417608 247716
rect 411864 247676 417608 247704
rect 411864 247664 411870 247676
rect 417602 247664 417608 247676
rect 417660 247664 417666 247716
rect 158070 246984 158076 247036
rect 158128 247024 158134 247036
rect 186314 247024 186320 247036
rect 158128 246996 186320 247024
rect 158128 246984 158134 246996
rect 186314 246984 186320 246996
rect 186372 246984 186378 247036
rect 169018 246916 169024 246968
rect 169076 246956 169082 246968
rect 186406 246956 186412 246968
rect 169076 246928 186412 246956
rect 169076 246916 169082 246928
rect 186406 246916 186412 246928
rect 186464 246916 186470 246968
rect 417326 246304 417332 246356
rect 417384 246344 417390 246356
rect 425974 246344 425980 246356
rect 417384 246316 425980 246344
rect 417384 246304 417390 246316
rect 425974 246304 425980 246316
rect 426032 246304 426038 246356
rect 411254 245624 411260 245676
rect 411312 245664 411318 245676
rect 417326 245664 417332 245676
rect 411312 245636 417332 245664
rect 411312 245624 411318 245636
rect 417326 245624 417332 245636
rect 417384 245624 417390 245676
rect 151170 245556 151176 245608
rect 151228 245596 151234 245608
rect 186314 245596 186320 245608
rect 151228 245568 186320 245596
rect 151228 245556 151234 245568
rect 186314 245556 186320 245568
rect 186372 245556 186378 245608
rect 520918 244264 520924 244316
rect 520976 244304 520982 244316
rect 579798 244304 579804 244316
rect 520976 244276 579804 244304
rect 520976 244264 520982 244276
rect 579798 244264 579804 244276
rect 579856 244264 579862 244316
rect 156690 244196 156696 244248
rect 156748 244236 156754 244248
rect 186314 244236 186320 244248
rect 156748 244208 186320 244236
rect 156748 244196 156754 244208
rect 186314 244196 186320 244208
rect 186372 244196 186378 244248
rect 410794 244196 410800 244248
rect 410852 244236 410858 244248
rect 417694 244236 417700 244248
rect 410852 244208 417700 244236
rect 410852 244196 410858 244208
rect 417694 244196 417700 244208
rect 417752 244196 417758 244248
rect 137370 242836 137376 242888
rect 137428 242876 137434 242888
rect 186314 242876 186320 242888
rect 137428 242848 186320 242876
rect 137428 242836 137434 242848
rect 186314 242836 186320 242848
rect 186372 242836 186378 242888
rect 411254 241816 411260 241868
rect 411312 241856 411318 241868
rect 414474 241856 414480 241868
rect 411312 241828 414480 241856
rect 411312 241816 411318 241828
rect 414474 241816 414480 241828
rect 414532 241856 414538 241868
rect 419166 241856 419172 241868
rect 414532 241828 419172 241856
rect 414532 241816 414538 241828
rect 419166 241816 419172 241828
rect 419224 241816 419230 241868
rect 155310 241408 155316 241460
rect 155368 241448 155374 241460
rect 186406 241448 186412 241460
rect 155368 241420 186412 241448
rect 155368 241408 155374 241420
rect 186406 241408 186412 241420
rect 186464 241408 186470 241460
rect 177482 241340 177488 241392
rect 177540 241380 177546 241392
rect 186314 241380 186320 241392
rect 177540 241352 186320 241380
rect 177540 241340 177546 241352
rect 186314 241340 186320 241352
rect 186372 241340 186378 241392
rect 144270 240048 144276 240100
rect 144328 240088 144334 240100
rect 186314 240088 186320 240100
rect 144328 240060 186320 240088
rect 144328 240048 144334 240060
rect 186314 240048 186320 240060
rect 186372 240048 186378 240100
rect 411254 240048 411260 240100
rect 411312 240088 411318 240100
rect 416222 240088 416228 240100
rect 411312 240060 416228 240088
rect 411312 240048 411318 240060
rect 416222 240048 416228 240060
rect 416280 240048 416286 240100
rect 162210 238688 162216 238740
rect 162268 238728 162274 238740
rect 186314 238728 186320 238740
rect 162268 238700 186320 238728
rect 162268 238688 162274 238700
rect 186314 238688 186320 238700
rect 186372 238688 186378 238740
rect 416682 238008 416688 238060
rect 416740 238048 416746 238060
rect 431494 238048 431500 238060
rect 416740 238020 431500 238048
rect 416740 238008 416746 238020
rect 431494 238008 431500 238020
rect 431552 238008 431558 238060
rect 411254 237396 411260 237448
rect 411312 237436 411318 237448
rect 415762 237436 415768 237448
rect 411312 237408 415768 237436
rect 411312 237396 411318 237408
rect 415762 237396 415768 237408
rect 415820 237436 415826 237448
rect 416682 237436 416688 237448
rect 415820 237408 416688 237436
rect 415820 237396 415826 237408
rect 416682 237396 416688 237408
rect 416740 237396 416746 237448
rect 176010 237328 176016 237380
rect 176068 237368 176074 237380
rect 186314 237368 186320 237380
rect 176068 237340 186320 237368
rect 176068 237328 176074 237340
rect 186314 237328 186320 237340
rect 186372 237328 186378 237380
rect 409414 237328 409420 237380
rect 409472 237368 409478 237380
rect 421834 237368 421840 237380
rect 409472 237340 421840 237368
rect 409472 237328 409478 237340
rect 421834 237328 421840 237340
rect 421892 237328 421898 237380
rect 176194 237260 176200 237312
rect 176252 237300 176258 237312
rect 186406 237300 186412 237312
rect 176252 237272 186412 237300
rect 176252 237260 176258 237272
rect 186406 237260 186412 237272
rect 186464 237260 186470 237312
rect 156598 235900 156604 235952
rect 156656 235940 156662 235952
rect 186314 235940 186320 235952
rect 156656 235912 186320 235940
rect 156656 235900 156662 235912
rect 186314 235900 186320 235912
rect 186372 235900 186378 235952
rect 173250 234540 173256 234592
rect 173308 234580 173314 234592
rect 186314 234580 186320 234592
rect 173308 234552 186320 234580
rect 173308 234540 173314 234552
rect 186314 234540 186320 234552
rect 186372 234540 186378 234592
rect 411254 233248 411260 233300
rect 411312 233288 411318 233300
rect 415854 233288 415860 233300
rect 411312 233260 415860 233288
rect 411312 233248 411318 233260
rect 415854 233248 415860 233260
rect 415912 233288 415918 233300
rect 420270 233288 420276 233300
rect 415912 233260 420276 233288
rect 415912 233248 415918 233260
rect 420270 233248 420276 233260
rect 420328 233248 420334 233300
rect 141510 233180 141516 233232
rect 141568 233220 141574 233232
rect 186314 233220 186320 233232
rect 141568 233192 186320 233220
rect 141568 233180 141574 233192
rect 186314 233180 186320 233192
rect 186372 233180 186378 233232
rect 469214 233180 469220 233232
rect 469272 233220 469278 233232
rect 579982 233220 579988 233232
rect 469272 233192 579988 233220
rect 469272 233180 469278 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 174538 233112 174544 233164
rect 174596 233152 174602 233164
rect 186406 233152 186412 233164
rect 174596 233124 186412 233152
rect 174596 233112 174602 233124
rect 186406 233112 186412 233124
rect 186464 233112 186470 233164
rect 133322 231752 133328 231804
rect 133380 231792 133386 231804
rect 186314 231792 186320 231804
rect 133380 231764 186320 231792
rect 133380 231752 133386 231764
rect 186314 231752 186320 231764
rect 186372 231752 186378 231804
rect 411346 231072 411352 231124
rect 411404 231112 411410 231124
rect 412082 231112 412088 231124
rect 411404 231084 412088 231112
rect 411404 231072 411410 231084
rect 412082 231072 412088 231084
rect 412140 231112 412146 231124
rect 434070 231112 434076 231124
rect 412140 231084 434076 231112
rect 412140 231072 412146 231084
rect 434070 231072 434076 231084
rect 434128 231072 434134 231124
rect 155218 230392 155224 230444
rect 155276 230432 155282 230444
rect 186314 230432 186320 230444
rect 155276 230404 186320 230432
rect 155276 230392 155282 230404
rect 186314 230392 186320 230404
rect 186372 230392 186378 230444
rect 415946 229712 415952 229764
rect 416004 229752 416010 229764
rect 428826 229752 428832 229764
rect 416004 229724 428832 229752
rect 416004 229712 416010 229724
rect 428826 229712 428832 229724
rect 428884 229712 428890 229764
rect 411254 229100 411260 229152
rect 411312 229140 411318 229152
rect 415946 229140 415952 229152
rect 411312 229112 415952 229140
rect 411312 229100 411318 229112
rect 415946 229100 415952 229112
rect 416004 229100 416010 229152
rect 138750 229032 138756 229084
rect 138808 229072 138814 229084
rect 186314 229072 186320 229084
rect 138808 229044 186320 229072
rect 138808 229032 138814 229044
rect 186314 229032 186320 229044
rect 186372 229032 186378 229084
rect 180150 228964 180156 229016
rect 180208 229004 180214 229016
rect 186406 229004 186412 229016
rect 180208 228976 186412 229004
rect 180208 228964 180214 228976
rect 186406 228964 186412 228976
rect 186464 228964 186470 229016
rect 409506 227740 409512 227792
rect 409564 227780 409570 227792
rect 414934 227780 414940 227792
rect 409564 227752 414940 227780
rect 409564 227740 409570 227752
rect 414934 227740 414940 227752
rect 414992 227740 414998 227792
rect 170398 227672 170404 227724
rect 170456 227712 170462 227724
rect 186314 227712 186320 227724
rect 170456 227684 186320 227712
rect 170456 227672 170462 227684
rect 186314 227672 186320 227684
rect 186372 227672 186378 227724
rect 157978 226244 157984 226296
rect 158036 226284 158042 226296
rect 186314 226284 186320 226296
rect 158036 226256 186320 226284
rect 158036 226244 158042 226256
rect 186314 226244 186320 226256
rect 186372 226244 186378 226296
rect 411530 225564 411536 225616
rect 411588 225604 411594 225616
rect 424686 225604 424692 225616
rect 411588 225576 424692 225604
rect 411588 225564 411594 225576
rect 424686 225564 424692 225576
rect 424744 225564 424750 225616
rect 152458 224884 152464 224936
rect 152516 224924 152522 224936
rect 186314 224924 186320 224936
rect 152516 224896 186320 224924
rect 152516 224884 152522 224896
rect 186314 224884 186320 224896
rect 186372 224884 186378 224936
rect 184382 224816 184388 224868
rect 184440 224856 184446 224868
rect 186406 224856 186412 224868
rect 184440 224828 186412 224856
rect 184440 224816 184446 224828
rect 186406 224816 186412 224828
rect 186464 224816 186470 224868
rect 415302 224204 415308 224256
rect 415360 224244 415366 224256
rect 429838 224244 429844 224256
rect 415360 224216 429844 224244
rect 415360 224204 415366 224216
rect 429838 224204 429844 224216
rect 429896 224204 429902 224256
rect 411254 223592 411260 223644
rect 411312 223632 411318 223644
rect 414566 223632 414572 223644
rect 411312 223604 414572 223632
rect 411312 223592 411318 223604
rect 414566 223592 414572 223604
rect 414624 223632 414630 223644
rect 415302 223632 415308 223644
rect 414624 223604 415308 223632
rect 414624 223592 414630 223604
rect 415302 223592 415308 223604
rect 415360 223592 415366 223644
rect 148318 223524 148324 223576
rect 148376 223564 148382 223576
rect 186314 223564 186320 223576
rect 148376 223536 186320 223564
rect 148376 223524 148382 223536
rect 186314 223524 186320 223536
rect 186372 223524 186378 223576
rect 164970 222096 164976 222148
rect 165028 222136 165034 222148
rect 186314 222136 186320 222148
rect 165028 222108 186320 222136
rect 165028 222096 165034 222108
rect 186314 222096 186320 222108
rect 186372 222096 186378 222148
rect 410794 222096 410800 222148
rect 410852 222136 410858 222148
rect 435726 222136 435732 222148
rect 410852 222108 435732 222136
rect 410852 222096 410858 222108
rect 435726 222096 435732 222108
rect 435784 222096 435790 222148
rect 159358 220736 159364 220788
rect 159416 220776 159422 220788
rect 186406 220776 186412 220788
rect 159416 220748 186412 220776
rect 159416 220736 159422 220748
rect 186406 220736 186412 220748
rect 186464 220736 186470 220788
rect 182910 220668 182916 220720
rect 182968 220708 182974 220720
rect 186498 220708 186504 220720
rect 182968 220680 186504 220708
rect 182968 220668 182974 220680
rect 186498 220668 186504 220680
rect 186556 220668 186562 220720
rect 411990 220056 411996 220108
rect 412048 220096 412054 220108
rect 419074 220096 419080 220108
rect 412048 220068 419080 220096
rect 412048 220056 412054 220068
rect 419074 220056 419080 220068
rect 419132 220056 419138 220108
rect 134702 219376 134708 219428
rect 134760 219416 134766 219428
rect 186314 219416 186320 219428
rect 134760 219388 186320 219416
rect 134760 219376 134766 219388
rect 186314 219376 186320 219388
rect 186372 219376 186378 219428
rect 460934 219376 460940 219428
rect 460992 219416 460998 219428
rect 580166 219416 580172 219428
rect 460992 219388 580172 219416
rect 460992 219376 460998 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 141418 217948 141424 218000
rect 141476 217988 141482 218000
rect 186314 217988 186320 218000
rect 141476 217960 186320 217988
rect 141476 217948 141482 217960
rect 186314 217948 186320 217960
rect 186372 217948 186378 218000
rect 411254 217268 411260 217320
rect 411312 217308 411318 217320
rect 414750 217308 414756 217320
rect 411312 217280 414756 217308
rect 411312 217268 411318 217280
rect 414750 217268 414756 217280
rect 414808 217308 414814 217320
rect 421742 217308 421748 217320
rect 414808 217280 421748 217308
rect 414808 217268 414814 217280
rect 421742 217268 421748 217280
rect 421800 217268 421806 217320
rect 145558 216588 145564 216640
rect 145616 216628 145622 216640
rect 186314 216628 186320 216640
rect 145616 216600 186320 216628
rect 145616 216588 145622 216600
rect 186314 216588 186320 216600
rect 186372 216588 186378 216640
rect 412082 216588 412088 216640
rect 412140 216628 412146 216640
rect 432782 216628 432788 216640
rect 412140 216600 432788 216628
rect 412140 216588 412146 216600
rect 432782 216588 432788 216600
rect 432840 216588 432846 216640
rect 134610 215228 134616 215280
rect 134668 215268 134674 215280
rect 186406 215268 186412 215280
rect 134668 215240 186412 215268
rect 134668 215228 134674 215240
rect 186406 215228 186412 215240
rect 186464 215228 186470 215280
rect 160738 215160 160744 215212
rect 160796 215200 160802 215212
rect 186314 215200 186320 215212
rect 160796 215172 186320 215200
rect 160796 215160 160802 215172
rect 186314 215160 186320 215172
rect 186372 215160 186378 215212
rect 142798 213868 142804 213920
rect 142856 213908 142862 213920
rect 186314 213908 186320 213920
rect 142856 213880 186320 213908
rect 142856 213868 142862 213880
rect 186314 213868 186320 213880
rect 186372 213868 186378 213920
rect 411254 213324 411260 213376
rect 411312 213364 411318 213376
rect 414658 213364 414664 213376
rect 411312 213336 414664 213364
rect 411312 213324 411318 213336
rect 414658 213324 414664 213336
rect 414716 213324 414722 213376
rect 177390 212440 177396 212492
rect 177448 212480 177454 212492
rect 186314 212480 186320 212492
rect 177448 212452 186320 212480
rect 177448 212440 177454 212452
rect 186314 212440 186320 212452
rect 186372 212440 186378 212492
rect 411254 211760 411260 211812
rect 411312 211800 411318 211812
rect 413186 211800 413192 211812
rect 411312 211772 413192 211800
rect 411312 211760 411318 211772
rect 413186 211760 413192 211772
rect 413244 211800 413250 211812
rect 432690 211800 432696 211812
rect 413244 211772 432696 211800
rect 413244 211760 413250 211772
rect 432690 211760 432696 211772
rect 432748 211760 432754 211812
rect 137278 211080 137284 211132
rect 137336 211120 137342 211132
rect 186314 211120 186320 211132
rect 137336 211092 186320 211120
rect 137336 211080 137342 211092
rect 186314 211080 186320 211092
rect 186372 211080 186378 211132
rect 178770 211012 178776 211064
rect 178828 211052 178834 211064
rect 186406 211052 186412 211064
rect 178828 211024 186412 211052
rect 178828 211012 178834 211024
rect 186406 211012 186412 211024
rect 186464 211012 186470 211064
rect 133230 209720 133236 209772
rect 133288 209760 133294 209772
rect 186314 209760 186320 209772
rect 133288 209732 186320 209760
rect 133288 209720 133294 209732
rect 186314 209720 186320 209732
rect 186372 209720 186378 209772
rect 411622 209040 411628 209092
rect 411680 209080 411686 209092
rect 431402 209080 431408 209092
rect 411680 209052 431408 209080
rect 411680 209040 411686 209052
rect 431402 209040 431408 209052
rect 431460 209040 431466 209092
rect 144178 208292 144184 208344
rect 144236 208332 144242 208344
rect 186314 208332 186320 208344
rect 144236 208304 186320 208332
rect 144236 208292 144242 208304
rect 186314 208292 186320 208304
rect 186372 208292 186378 208344
rect 411346 207612 411352 207664
rect 411404 207652 411410 207664
rect 428642 207652 428648 207664
rect 411404 207624 428648 207652
rect 411404 207612 411410 207624
rect 428642 207612 428648 207624
rect 428700 207612 428706 207664
rect 135898 206932 135904 206984
rect 135956 206972 135962 206984
rect 186314 206972 186320 206984
rect 135956 206944 186320 206972
rect 135956 206932 135962 206944
rect 186314 206932 186320 206944
rect 186372 206932 186378 206984
rect 181530 206864 181536 206916
rect 181588 206904 181594 206916
rect 186406 206904 186412 206916
rect 181588 206876 186412 206904
rect 181588 206864 181594 206876
rect 186406 206864 186412 206876
rect 186464 206864 186470 206916
rect 519538 205640 519544 205692
rect 519596 205680 519602 205692
rect 580166 205680 580172 205692
rect 519596 205652 580172 205680
rect 519596 205640 519602 205652
rect 580166 205640 580172 205652
rect 580224 205640 580230 205692
rect 162118 205572 162124 205624
rect 162176 205612 162182 205624
rect 186314 205612 186320 205624
rect 162176 205584 186320 205612
rect 162176 205572 162182 205584
rect 186314 205572 186320 205584
rect 186372 205572 186378 205624
rect 413922 204892 413928 204944
rect 413980 204932 413986 204944
rect 436830 204932 436836 204944
rect 413980 204904 436836 204932
rect 413980 204892 413986 204904
rect 436830 204892 436836 204904
rect 436888 204892 436894 204944
rect 411254 204280 411260 204332
rect 411312 204320 411318 204332
rect 413370 204320 413376 204332
rect 411312 204292 413376 204320
rect 411312 204280 411318 204292
rect 413370 204280 413376 204292
rect 413428 204320 413434 204332
rect 413922 204320 413928 204332
rect 413428 204292 413928 204320
rect 413428 204280 413434 204292
rect 413922 204280 413928 204292
rect 413980 204280 413986 204332
rect 146938 204212 146944 204264
rect 146996 204252 147002 204264
rect 186314 204252 186320 204264
rect 146996 204224 186320 204252
rect 146996 204212 147002 204224
rect 186314 204212 186320 204224
rect 186372 204212 186378 204264
rect 415302 203532 415308 203584
rect 415360 203572 415366 203584
rect 430022 203572 430028 203584
rect 415360 203544 430028 203572
rect 415360 203532 415366 203544
rect 430022 203532 430028 203544
rect 430080 203532 430086 203584
rect 411254 203056 411260 203108
rect 411312 203096 411318 203108
rect 414842 203096 414848 203108
rect 411312 203068 414848 203096
rect 411312 203056 411318 203068
rect 414842 203056 414848 203068
rect 414900 203096 414906 203108
rect 415302 203096 415308 203108
rect 414900 203068 415308 203096
rect 414900 203056 414906 203068
rect 415302 203056 415308 203068
rect 415360 203056 415366 203108
rect 138658 202784 138664 202836
rect 138716 202824 138722 202836
rect 186406 202824 186412 202836
rect 138716 202796 186412 202824
rect 138716 202784 138722 202796
rect 186406 202784 186412 202796
rect 186464 202784 186470 202836
rect 173342 202716 173348 202768
rect 173400 202756 173406 202768
rect 186314 202756 186320 202768
rect 173400 202728 186320 202756
rect 173400 202716 173406 202728
rect 186314 202716 186320 202728
rect 186372 202716 186378 202768
rect 412634 202104 412640 202156
rect 412692 202144 412698 202156
rect 536834 202144 536840 202156
rect 412692 202116 536840 202144
rect 412692 202104 412698 202116
rect 536834 202104 536840 202116
rect 536892 202104 536898 202156
rect 134518 201424 134524 201476
rect 134576 201464 134582 201476
rect 186314 201464 186320 201476
rect 134576 201436 186320 201464
rect 134576 201424 134582 201436
rect 186314 201424 186320 201436
rect 186372 201424 186378 201476
rect 411254 200744 411260 200796
rect 411312 200784 411318 200796
rect 422938 200784 422944 200796
rect 411312 200756 422944 200784
rect 411312 200744 411318 200756
rect 422938 200744 422944 200756
rect 422996 200744 423002 200796
rect 401042 199996 401048 200048
rect 401100 200036 401106 200048
rect 412266 200036 412272 200048
rect 401100 200008 412272 200036
rect 401100 199996 401106 200008
rect 412266 199996 412272 200008
rect 412324 199996 412330 200048
rect 404998 199928 405004 199980
rect 405056 199968 405062 199980
rect 415394 199968 415400 199980
rect 405056 199940 415400 199968
rect 405056 199928 405062 199940
rect 415394 199928 415400 199940
rect 415452 199928 415458 199980
rect 400950 199860 400956 199912
rect 401008 199900 401014 199912
rect 411438 199900 411444 199912
rect 401008 199872 411444 199900
rect 401008 199860 401014 199872
rect 411438 199860 411444 199872
rect 411496 199860 411502 199912
rect 399570 199792 399576 199844
rect 399628 199832 399634 199844
rect 412174 199832 412180 199844
rect 399628 199804 412180 199832
rect 399628 199792 399634 199804
rect 412174 199792 412180 199804
rect 412232 199792 412238 199844
rect 407758 199724 407764 199776
rect 407816 199764 407822 199776
rect 419810 199764 419816 199776
rect 407816 199736 419816 199764
rect 407816 199724 407822 199736
rect 419810 199724 419816 199736
rect 419868 199724 419874 199776
rect 398374 199656 398380 199708
rect 398432 199696 398438 199708
rect 410426 199696 410432 199708
rect 398432 199668 410432 199696
rect 398432 199656 398438 199668
rect 410426 199656 410432 199668
rect 410484 199656 410490 199708
rect 194594 199588 194600 199640
rect 194652 199628 194658 199640
rect 195606 199628 195612 199640
rect 194652 199600 195612 199628
rect 194652 199588 194658 199600
rect 195606 199588 195612 199600
rect 195664 199588 195670 199640
rect 399202 199588 399208 199640
rect 399260 199628 399266 199640
rect 411806 199628 411812 199640
rect 399260 199600 411812 199628
rect 399260 199588 399266 199600
rect 411806 199588 411812 199600
rect 411864 199588 411870 199640
rect 406378 199520 406384 199572
rect 406436 199560 406442 199572
rect 419718 199560 419724 199572
rect 406436 199532 419724 199560
rect 406436 199520 406442 199532
rect 419718 199520 419724 199532
rect 419776 199520 419782 199572
rect 393222 199452 393228 199504
rect 393280 199492 393286 199504
rect 411254 199492 411260 199504
rect 393280 199464 411260 199492
rect 393280 199452 393286 199464
rect 411254 199452 411260 199464
rect 411312 199452 411318 199504
rect 261846 199384 261852 199436
rect 261904 199424 261910 199436
rect 552014 199424 552020 199436
rect 261904 199396 552020 199424
rect 261904 199384 261910 199396
rect 552014 199384 552020 199396
rect 552072 199384 552078 199436
rect 189718 199112 189724 199164
rect 189776 199152 189782 199164
rect 239582 199152 239588 199164
rect 189776 199124 239588 199152
rect 189776 199112 189782 199124
rect 239582 199112 239588 199124
rect 239640 199112 239646 199164
rect 188338 199044 188344 199096
rect 188396 199084 188402 199096
rect 259638 199084 259644 199096
rect 188396 199056 259644 199084
rect 188396 199044 188402 199056
rect 259638 199044 259644 199056
rect 259696 199044 259702 199096
rect 189810 198976 189816 199028
rect 189868 199016 189874 199028
rect 327534 199016 327540 199028
rect 189868 198988 327540 199016
rect 189868 198976 189874 198988
rect 327534 198976 327540 198988
rect 327592 198976 327598 199028
rect 185578 198908 185584 198960
rect 185636 198948 185642 198960
rect 271966 198948 271972 198960
rect 185636 198920 271972 198948
rect 185636 198908 185642 198920
rect 271966 198908 271972 198920
rect 272024 198908 272030 198960
rect 296162 198908 296168 198960
rect 296220 198948 296226 198960
rect 436738 198948 436744 198960
rect 296220 198920 436744 198948
rect 296220 198908 296226 198920
rect 436738 198908 436744 198920
rect 436796 198908 436802 198960
rect 131850 198840 131856 198892
rect 131908 198880 131914 198892
rect 311986 198880 311992 198892
rect 131908 198852 311992 198880
rect 131908 198840 131914 198852
rect 311986 198840 311992 198852
rect 312044 198840 312050 198892
rect 133138 198772 133144 198824
rect 133196 198812 133202 198824
rect 319622 198812 319628 198824
rect 133196 198784 319628 198812
rect 133196 198772 133202 198784
rect 319622 198772 319628 198784
rect 319680 198772 319686 198824
rect 344186 198772 344192 198824
rect 344244 198812 344250 198824
rect 425698 198812 425704 198824
rect 344244 198784 425704 198812
rect 344244 198772 344250 198784
rect 425698 198772 425704 198784
rect 425756 198772 425762 198824
rect 189994 198704 190000 198756
rect 190052 198744 190058 198756
rect 194594 198744 194600 198756
rect 190052 198716 194600 198744
rect 190052 198704 190058 198716
rect 194594 198704 194600 198716
rect 194652 198704 194658 198756
rect 208210 198704 208216 198756
rect 208268 198744 208274 198756
rect 435450 198744 435456 198756
rect 208268 198716 435456 198744
rect 208268 198704 208274 198716
rect 435450 198704 435456 198716
rect 435508 198704 435514 198756
rect 182818 198636 182824 198688
rect 182876 198676 182882 198688
rect 379606 198676 379612 198688
rect 182876 198648 379612 198676
rect 182876 198636 182882 198648
rect 379606 198636 379612 198648
rect 379664 198636 379670 198688
rect 397362 198636 397368 198688
rect 397420 198676 397426 198688
rect 413370 198676 413376 198688
rect 397420 198648 413376 198676
rect 397420 198636 397426 198648
rect 413370 198636 413376 198648
rect 413428 198636 413434 198688
rect 184198 198568 184204 198620
rect 184256 198608 184262 198620
rect 351454 198608 351460 198620
rect 184256 198580 351460 198608
rect 184256 198568 184262 198580
rect 351454 198568 351460 198580
rect 351512 198568 351518 198620
rect 368106 198568 368112 198620
rect 368164 198608 368170 198620
rect 432598 198608 432604 198620
rect 368164 198580 432604 198608
rect 368164 198568 368170 198580
rect 432598 198568 432604 198580
rect 432656 198568 432662 198620
rect 188430 198500 188436 198552
rect 188488 198540 188494 198552
rect 339494 198540 339500 198552
rect 188488 198512 339500 198540
rect 188488 198500 188494 198512
rect 339494 198500 339500 198512
rect 339552 198500 339558 198552
rect 364242 198500 364248 198552
rect 364300 198540 364306 198552
rect 412634 198540 412640 198552
rect 364300 198512 412640 198540
rect 364300 198500 364306 198512
rect 412634 198500 412640 198512
rect 412692 198500 412698 198552
rect 188522 198432 188528 198484
rect 188580 198472 188586 198484
rect 323486 198472 323492 198484
rect 188580 198444 323492 198472
rect 188580 198432 188586 198444
rect 323486 198432 323492 198444
rect 323544 198432 323550 198484
rect 397270 198432 397276 198484
rect 397328 198472 397334 198484
rect 413186 198472 413192 198484
rect 397328 198444 413192 198472
rect 397328 198432 397334 198444
rect 413186 198432 413192 198444
rect 413244 198432 413250 198484
rect 163498 198364 163504 198416
rect 163556 198404 163562 198416
rect 267734 198404 267740 198416
rect 163556 198376 267740 198404
rect 163556 198364 163562 198376
rect 267734 198364 267740 198376
rect 267792 198364 267798 198416
rect 397178 198364 397184 198416
rect 397236 198404 397242 198416
rect 414750 198404 414756 198416
rect 397236 198376 414756 198404
rect 397236 198364 397242 198376
rect 414750 198364 414756 198376
rect 414808 198364 414814 198416
rect 184290 198296 184296 198348
rect 184348 198336 184354 198348
rect 279510 198336 279516 198348
rect 184348 198308 279516 198336
rect 184348 198296 184354 198308
rect 279510 198296 279516 198308
rect 279568 198296 279574 198348
rect 395798 198296 395804 198348
rect 395856 198336 395862 198348
rect 414106 198336 414112 198348
rect 395856 198308 414112 198336
rect 395856 198296 395862 198308
rect 414106 198296 414112 198308
rect 414164 198296 414170 198348
rect 177298 198228 177304 198280
rect 177356 198268 177362 198280
rect 255590 198268 255596 198280
rect 177356 198240 255596 198268
rect 177356 198228 177362 198240
rect 255590 198228 255596 198240
rect 255648 198228 255654 198280
rect 395890 198228 395896 198280
rect 395948 198268 395954 198280
rect 414382 198268 414388 198280
rect 395948 198240 414388 198268
rect 395948 198228 395954 198240
rect 414382 198228 414388 198240
rect 414440 198228 414446 198280
rect 175918 198160 175924 198212
rect 175976 198200 175982 198212
rect 243630 198200 243636 198212
rect 175976 198172 243636 198200
rect 175976 198160 175982 198172
rect 243630 198160 243636 198172
rect 243688 198160 243694 198212
rect 395706 198160 395712 198212
rect 395764 198200 395770 198212
rect 414290 198200 414296 198212
rect 395764 198172 414296 198200
rect 395764 198160 395770 198172
rect 414290 198160 414296 198172
rect 414348 198160 414354 198212
rect 185670 198092 185676 198144
rect 185728 198132 185734 198144
rect 247494 198132 247500 198144
rect 185728 198104 247500 198132
rect 185728 198092 185734 198104
rect 247494 198092 247500 198104
rect 247552 198092 247558 198144
rect 395430 198092 395436 198144
rect 395488 198132 395494 198144
rect 395488 198104 395752 198132
rect 395488 198092 395494 198104
rect 178678 198024 178684 198076
rect 178736 198064 178742 198076
rect 235534 198064 235540 198076
rect 178736 198036 235540 198064
rect 178736 198024 178742 198036
rect 235534 198024 235540 198036
rect 235592 198024 235598 198076
rect 323578 198024 323584 198076
rect 323636 198064 323642 198076
rect 395614 198064 395620 198076
rect 323636 198036 395620 198064
rect 323636 198024 323642 198036
rect 395614 198024 395620 198036
rect 395672 198024 395678 198076
rect 395724 198064 395752 198104
rect 396718 198092 396724 198144
rect 396776 198132 396782 198144
rect 415486 198132 415492 198144
rect 396776 198104 415492 198132
rect 396776 198092 396782 198104
rect 415486 198092 415492 198104
rect 415544 198092 415550 198144
rect 414198 198064 414204 198076
rect 395724 198036 414204 198064
rect 414198 198024 414204 198036
rect 414256 198024 414262 198076
rect 164878 197956 164884 198008
rect 164936 197996 164942 198008
rect 219526 197996 219532 198008
rect 164936 197968 219532 197996
rect 164936 197956 164942 197968
rect 219526 197956 219532 197968
rect 219584 197956 219590 198008
rect 224218 197956 224224 198008
rect 224276 197996 224282 198008
rect 261846 197996 261852 198008
rect 224276 197968 261852 197996
rect 224276 197956 224282 197968
rect 261846 197956 261852 197968
rect 261904 197956 261910 198008
rect 264146 197956 264152 198008
rect 264204 197996 264210 198008
rect 280246 197996 280252 198008
rect 264204 197968 280252 197996
rect 264204 197956 264210 197968
rect 280246 197956 280252 197968
rect 280304 197956 280310 198008
rect 319438 197956 319444 198008
rect 319496 197996 319502 198008
rect 391566 197996 391572 198008
rect 319496 197968 391572 197996
rect 319496 197956 319502 197968
rect 391566 197956 391572 197968
rect 391624 197956 391630 198008
rect 395522 197956 395528 198008
rect 395580 197996 395586 198008
rect 415578 197996 415584 198008
rect 395580 197968 415584 197996
rect 395580 197956 395586 197968
rect 415578 197956 415584 197968
rect 415636 197956 415642 198008
rect 189902 197888 189908 197940
rect 189960 197928 189966 197940
rect 227714 197928 227720 197940
rect 189960 197900 227720 197928
rect 189960 197888 189966 197900
rect 227714 197888 227720 197900
rect 227772 197888 227778 197940
rect 403618 197888 403624 197940
rect 403676 197928 403682 197940
rect 418338 197928 418344 197940
rect 403676 197900 418344 197928
rect 403676 197888 403682 197900
rect 418338 197888 418344 197900
rect 418396 197888 418402 197940
rect 188890 197820 188896 197872
rect 188948 197860 188954 197872
rect 212534 197860 212540 197872
rect 188948 197832 212540 197860
rect 188948 197820 188954 197832
rect 212534 197820 212540 197832
rect 212592 197820 212598 197872
rect 399754 197820 399760 197872
rect 399812 197860 399818 197872
rect 411346 197860 411352 197872
rect 399812 197832 411352 197860
rect 399812 197820 399818 197832
rect 411346 197820 411352 197832
rect 411404 197820 411410 197872
rect 186222 197752 186228 197804
rect 186280 197792 186286 197804
rect 200114 197792 200120 197804
rect 186280 197764 200120 197792
rect 186280 197752 186286 197764
rect 200114 197752 200120 197764
rect 200172 197752 200178 197804
rect 400858 197752 400864 197804
rect 400916 197792 400922 197804
rect 411714 197792 411720 197804
rect 400916 197764 411720 197792
rect 400916 197752 400922 197764
rect 411714 197752 411720 197764
rect 411772 197752 411778 197804
rect 395614 197344 395620 197396
rect 395672 197384 395678 197396
rect 395798 197384 395804 197396
rect 395672 197356 395804 197384
rect 395672 197344 395678 197356
rect 395798 197344 395804 197356
rect 395856 197344 395862 197396
rect 148962 197276 148968 197328
rect 149020 197316 149026 197328
rect 383654 197316 383660 197328
rect 149020 197288 383660 197316
rect 149020 197276 149026 197288
rect 383654 197276 383660 197288
rect 383712 197276 383718 197328
rect 151078 197208 151084 197260
rect 151136 197248 151142 197260
rect 375558 197248 375564 197260
rect 151136 197220 375564 197248
rect 151136 197208 151142 197220
rect 375558 197208 375564 197220
rect 375616 197208 375622 197260
rect 131022 197140 131028 197192
rect 131080 197180 131086 197192
rect 355502 197180 355508 197192
rect 131080 197152 355508 197180
rect 131080 197140 131086 197152
rect 355502 197140 355508 197152
rect 355560 197140 355566 197192
rect 131758 197072 131764 197124
rect 131816 197112 131822 197124
rect 331582 197112 331588 197124
rect 131816 197084 331588 197112
rect 131816 197072 131822 197084
rect 331582 197072 331588 197084
rect 331640 197072 331646 197124
rect 130470 197004 130476 197056
rect 130528 197044 130534 197056
rect 315574 197044 315580 197056
rect 130528 197016 315580 197044
rect 130528 197004 130534 197016
rect 315574 197004 315580 197016
rect 315632 197004 315638 197056
rect 130378 196936 130384 196988
rect 130436 196976 130442 196988
rect 303614 196976 303620 196988
rect 130436 196948 303620 196976
rect 130436 196936 130442 196948
rect 303614 196936 303620 196948
rect 303672 196936 303678 196988
rect 397822 196800 397828 196852
rect 397880 196840 397886 196852
rect 409322 196840 409328 196852
rect 397880 196812 409328 196840
rect 397880 196800 397886 196812
rect 409322 196800 409328 196812
rect 409380 196800 409386 196852
rect 398742 196732 398748 196784
rect 398800 196772 398806 196784
rect 410334 196772 410340 196784
rect 398800 196744 410340 196772
rect 398800 196732 398806 196744
rect 410334 196732 410340 196744
rect 410392 196732 410398 196784
rect 399110 196664 399116 196716
rect 399168 196704 399174 196716
rect 411898 196704 411904 196716
rect 399168 196676 411904 196704
rect 399168 196664 399174 196676
rect 411898 196664 411904 196676
rect 411956 196664 411962 196716
rect 399018 196596 399024 196648
rect 399076 196636 399082 196648
rect 411990 196636 411996 196648
rect 399076 196608 411996 196636
rect 399076 196596 399082 196608
rect 411990 196596 411996 196608
rect 412048 196596 412054 196648
rect 396994 195916 397000 195968
rect 397052 195956 397058 195968
rect 415946 195956 415952 195968
rect 397052 195928 415952 195956
rect 397052 195916 397058 195928
rect 415946 195916 415952 195928
rect 416004 195916 416010 195968
rect 395982 195848 395988 195900
rect 396040 195888 396046 195900
rect 415854 195888 415860 195900
rect 396040 195860 415860 195888
rect 396040 195848 396046 195860
rect 415854 195848 415860 195860
rect 415912 195848 415918 195900
rect 394418 195780 394424 195832
rect 394476 195820 394482 195832
rect 414474 195820 414480 195832
rect 394476 195792 414480 195820
rect 394476 195780 394482 195792
rect 414474 195780 414480 195792
rect 414532 195780 414538 195832
rect 396902 195712 396908 195764
rect 396960 195752 396966 195764
rect 417142 195752 417148 195764
rect 396960 195724 417148 195752
rect 396960 195712 396966 195724
rect 417142 195712 417148 195724
rect 417200 195712 417206 195764
rect 392670 195644 392676 195696
rect 392728 195684 392734 195696
rect 413094 195684 413100 195696
rect 392728 195656 413100 195684
rect 392728 195644 392734 195656
rect 413094 195644 413100 195656
rect 413152 195644 413158 195696
rect 392578 195576 392584 195628
rect 392636 195616 392642 195628
rect 414014 195616 414020 195628
rect 392636 195588 414020 195616
rect 392636 195576 392642 195588
rect 414014 195576 414020 195588
rect 414072 195576 414078 195628
rect 393130 195508 393136 195560
rect 393188 195548 393194 195560
rect 415762 195548 415768 195560
rect 393188 195520 415768 195548
rect 393188 195508 393194 195520
rect 415762 195508 415768 195520
rect 415820 195508 415826 195560
rect 394326 195440 394332 195492
rect 394384 195480 394390 195492
rect 417050 195480 417056 195492
rect 394384 195452 417056 195480
rect 394384 195440 394390 195452
rect 417050 195440 417056 195452
rect 417108 195440 417114 195492
rect 392946 195372 392952 195424
rect 393004 195412 393010 195424
rect 415670 195412 415676 195424
rect 393004 195384 415676 195412
rect 393004 195372 393010 195384
rect 415670 195372 415676 195384
rect 415728 195372 415734 195424
rect 393038 195304 393044 195356
rect 393096 195344 393102 195356
rect 417234 195344 417240 195356
rect 393096 195316 417240 195344
rect 393096 195304 393102 195316
rect 417234 195304 417240 195316
rect 417292 195304 417298 195356
rect 400122 195236 400128 195288
rect 400180 195276 400186 195288
rect 503714 195276 503720 195288
rect 400180 195248 503720 195276
rect 400180 195236 400186 195248
rect 503714 195236 503720 195248
rect 503772 195236 503778 195288
rect 397086 195168 397092 195220
rect 397144 195208 397150 195220
rect 414566 195208 414572 195220
rect 397144 195180 414572 195208
rect 397144 195168 397150 195180
rect 414566 195168 414572 195180
rect 414624 195168 414630 195220
rect 403802 195100 403808 195152
rect 403860 195140 403866 195152
rect 421006 195140 421012 195152
rect 403860 195112 421012 195140
rect 403860 195100 403866 195112
rect 421006 195100 421012 195112
rect 421064 195100 421070 195152
rect 403710 195032 403716 195084
rect 403768 195072 403774 195084
rect 418246 195072 418252 195084
rect 403768 195044 418252 195072
rect 403768 195032 403774 195044
rect 418246 195032 418252 195044
rect 418304 195032 418310 195084
rect 204162 193808 204168 193860
rect 204220 193848 204226 193860
rect 284938 193848 284944 193860
rect 204220 193820 284944 193848
rect 204220 193808 204226 193820
rect 284938 193808 284944 193820
rect 284996 193808 285002 193860
rect 452654 193128 452660 193180
rect 452712 193168 452718 193180
rect 580166 193168 580172 193180
rect 452712 193140 580172 193168
rect 452712 193128 452718 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 401226 192924 401232 192976
rect 401284 192964 401290 192976
rect 419626 192964 419632 192976
rect 401284 192936 419632 192964
rect 401284 192924 401290 192936
rect 419626 192924 419632 192936
rect 419684 192924 419690 192976
rect 394602 192856 394608 192908
rect 394660 192896 394666 192908
rect 414842 192896 414848 192908
rect 394660 192868 414848 192896
rect 394660 192856 394666 192868
rect 414842 192856 414848 192868
rect 414900 192856 414906 192908
rect 401134 192788 401140 192840
rect 401192 192828 401198 192840
rect 420914 192828 420920 192840
rect 401192 192800 420920 192828
rect 401192 192788 401198 192800
rect 420914 192788 420920 192800
rect 420972 192788 420978 192840
rect 394510 192720 394516 192772
rect 394568 192760 394574 192772
rect 414658 192760 414664 192772
rect 394568 192732 414664 192760
rect 394568 192720 394574 192732
rect 414658 192720 414664 192732
rect 414716 192720 414722 192772
rect 392762 192652 392768 192704
rect 392820 192692 392826 192704
rect 416866 192692 416872 192704
rect 392820 192664 416872 192692
rect 392820 192652 392826 192664
rect 416866 192652 416872 192664
rect 416924 192652 416930 192704
rect 393958 192584 393964 192636
rect 394016 192624 394022 192636
rect 418154 192624 418160 192636
rect 394016 192596 418160 192624
rect 394016 192584 394022 192596
rect 418154 192584 418160 192596
rect 418212 192584 418218 192636
rect 389818 192516 389824 192568
rect 389876 192556 389882 192568
rect 416774 192556 416780 192568
rect 389876 192528 416780 192556
rect 389876 192516 389882 192528
rect 416774 192516 416780 192528
rect 416832 192516 416838 192568
rect 189258 192448 189264 192500
rect 189316 192488 189322 192500
rect 224954 192488 224960 192500
rect 189316 192460 224960 192488
rect 189316 192448 189322 192460
rect 224954 192448 224960 192460
rect 225012 192448 225018 192500
rect 282178 192448 282184 192500
rect 282236 192488 282242 192500
rect 413002 192488 413008 192500
rect 282236 192460 413008 192488
rect 282236 192448 282242 192460
rect 413002 192448 413008 192460
rect 413060 192448 413066 192500
rect 400674 191836 400680 191888
rect 400732 191876 400738 191888
rect 404262 191876 404268 191888
rect 400732 191848 404268 191876
rect 400732 191836 400738 191848
rect 404262 191836 404268 191848
rect 404320 191836 404326 191888
rect 188706 191156 188712 191208
rect 188764 191196 188770 191208
rect 235994 191196 236000 191208
rect 188764 191168 236000 191196
rect 188764 191156 188770 191168
rect 235994 191156 236000 191168
rect 236052 191156 236058 191208
rect 187142 191088 187148 191140
rect 187200 191128 187206 191140
rect 509234 191128 509240 191140
rect 187200 191100 509240 191128
rect 187200 191088 187206 191100
rect 509234 191088 509240 191100
rect 509292 191088 509298 191140
rect 189166 189728 189172 189780
rect 189224 189768 189230 189780
rect 248414 189768 248420 189780
rect 189224 189740 248420 189768
rect 189224 189728 189230 189740
rect 248414 189728 248420 189740
rect 248472 189728 248478 189780
rect 282362 189728 282368 189780
rect 282420 189768 282426 189780
rect 412910 189768 412916 189780
rect 282420 189740 412916 189768
rect 282420 189728 282426 189740
rect 412910 189728 412916 189740
rect 412968 189728 412974 189780
rect 169846 188300 169852 188352
rect 169904 188340 169910 188352
rect 407114 188340 407120 188352
rect 169904 188312 407120 188340
rect 169904 188300 169910 188312
rect 407114 188300 407120 188312
rect 407172 188300 407178 188352
rect 397454 187688 397460 187740
rect 397512 187728 397518 187740
rect 400674 187728 400680 187740
rect 397512 187700 400680 187728
rect 397512 187688 397518 187700
rect 400674 187688 400680 187700
rect 400732 187688 400738 187740
rect 187234 186940 187240 186992
rect 187292 186980 187298 186992
rect 286318 186980 286324 186992
rect 187292 186952 286324 186980
rect 187292 186940 187298 186952
rect 286318 186940 286324 186952
rect 286376 186940 286382 186992
rect 187510 184152 187516 184204
rect 187568 184192 187574 184204
rect 395338 184192 395344 184204
rect 187568 184164 395344 184192
rect 187568 184152 187574 184164
rect 395338 184152 395344 184164
rect 395396 184152 395402 184204
rect 390554 182860 390560 182912
rect 390612 182900 390618 182912
rect 397454 182900 397460 182912
rect 390612 182872 397460 182900
rect 390612 182860 390618 182872
rect 397454 182860 397460 182872
rect 397512 182860 397518 182912
rect 188798 182792 188804 182844
rect 188856 182832 188862 182844
rect 466454 182832 466460 182844
rect 188856 182804 466460 182832
rect 188856 182792 188862 182804
rect 466454 182792 466460 182804
rect 466512 182792 466518 182844
rect 387334 181024 387340 181076
rect 387392 181064 387398 181076
rect 390554 181064 390560 181076
rect 387392 181036 390560 181064
rect 387392 181024 387398 181036
rect 390554 181024 390560 181036
rect 390612 181024 390618 181076
rect 186866 180072 186872 180124
rect 186924 180112 186930 180124
rect 309778 180112 309784 180124
rect 186924 180084 309784 180112
rect 186924 180072 186930 180084
rect 309778 180072 309784 180084
rect 309836 180072 309842 180124
rect 442994 179324 443000 179376
rect 443052 179364 443058 179376
rect 580166 179364 580172 179376
rect 443052 179336 580172 179364
rect 443052 179324 443058 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 274634 178644 274640 178696
rect 274692 178684 274698 178696
rect 349798 178684 349804 178696
rect 274692 178656 349804 178684
rect 274692 178644 274698 178656
rect 349798 178644 349804 178656
rect 349856 178644 349862 178696
rect 187602 177284 187608 177336
rect 187660 177324 187666 177336
rect 305638 177324 305644 177336
rect 187660 177296 305644 177324
rect 187660 177284 187666 177296
rect 305638 177284 305644 177296
rect 305696 177284 305702 177336
rect 384298 175176 384304 175228
rect 384356 175216 384362 175228
rect 387334 175216 387340 175228
rect 384356 175188 387340 175216
rect 384356 175176 384362 175188
rect 387334 175176 387340 175188
rect 387392 175176 387398 175228
rect 382274 168376 382280 168428
rect 382332 168416 382338 168428
rect 384298 168416 384304 168428
rect 382332 168388 384304 168416
rect 382332 168376 382338 168388
rect 384298 168376 384304 168388
rect 384356 168376 384362 168428
rect 289078 165588 289084 165640
rect 289136 165628 289142 165640
rect 580166 165628 580172 165640
rect 289136 165600 580172 165628
rect 289136 165588 289142 165600
rect 580166 165588 580172 165600
rect 580224 165588 580230 165640
rect 381538 164772 381544 164824
rect 381596 164812 381602 164824
rect 382274 164812 382280 164824
rect 381596 164784 382280 164812
rect 381596 164772 381602 164784
rect 382274 164772 382280 164784
rect 382332 164772 382338 164824
rect 187326 155184 187332 155236
rect 187384 155224 187390 155236
rect 510890 155224 510896 155236
rect 187384 155196 510896 155224
rect 187384 155184 187390 155196
rect 510890 155184 510896 155196
rect 510948 155184 510954 155236
rect 379514 154300 379520 154352
rect 379572 154340 379578 154352
rect 381538 154340 381544 154352
rect 379572 154312 381544 154340
rect 379572 154300 379578 154312
rect 381538 154300 381544 154312
rect 381596 154300 381602 154352
rect 428458 153824 428464 153876
rect 428516 153864 428522 153876
rect 580626 153864 580632 153876
rect 428516 153836 580632 153864
rect 428516 153824 428522 153836
rect 580626 153824 580632 153836
rect 580684 153824 580690 153876
rect 431218 153144 431224 153196
rect 431276 153184 431282 153196
rect 580166 153184 580172 153196
rect 431276 153156 580172 153184
rect 431276 153144 431282 153156
rect 580166 153144 580172 153156
rect 580224 153144 580230 153196
rect 170214 152464 170220 152516
rect 170272 152504 170278 152516
rect 371234 152504 371240 152516
rect 170272 152476 371240 152504
rect 170272 152464 170278 152476
rect 371234 152464 371240 152476
rect 371292 152464 371298 152516
rect 168926 151036 168932 151088
rect 168984 151076 168990 151088
rect 282914 151076 282920 151088
rect 168984 151048 282920 151076
rect 168984 151036 168990 151048
rect 282914 151036 282920 151048
rect 282972 151036 282978 151088
rect 424318 151036 424324 151088
rect 424376 151076 424382 151088
rect 580534 151076 580540 151088
rect 424376 151048 580540 151076
rect 424376 151036 424382 151048
rect 580534 151036 580540 151048
rect 580592 151036 580598 151088
rect 188982 149676 188988 149728
rect 189040 149716 189046 149728
rect 281534 149716 281540 149728
rect 189040 149688 281540 149716
rect 189040 149676 189046 149688
rect 281534 149676 281540 149688
rect 281592 149676 281598 149728
rect 282270 149676 282276 149728
rect 282328 149716 282334 149728
rect 412818 149716 412824 149728
rect 282328 149688 412824 149716
rect 282328 149676 282334 149688
rect 412818 149676 412824 149688
rect 412876 149676 412882 149728
rect 421558 149676 421564 149728
rect 421616 149716 421622 149728
rect 580350 149716 580356 149728
rect 421616 149688 580356 149716
rect 421616 149676 421622 149688
rect 580350 149676 580356 149688
rect 580408 149676 580414 149728
rect 168834 148316 168840 148368
rect 168892 148356 168898 148368
rect 299474 148356 299480 148368
rect 168892 148328 299480 148356
rect 168892 148316 168898 148328
rect 299474 148316 299480 148328
rect 299532 148316 299538 148368
rect 425790 148316 425796 148368
rect 425848 148356 425854 148368
rect 580258 148356 580264 148368
rect 425848 148328 580264 148356
rect 425848 148316 425854 148328
rect 580258 148316 580264 148328
rect 580316 148316 580322 148368
rect 406010 146956 406016 147008
rect 406068 146996 406074 147008
rect 439498 146996 439504 147008
rect 406068 146968 439504 146996
rect 406068 146956 406074 146968
rect 439498 146956 439504 146968
rect 439556 146956 439562 147008
rect 439590 146956 439596 147008
rect 439648 146996 439654 147008
rect 512270 146996 512276 147008
rect 439648 146968 512276 146996
rect 439648 146956 439654 146968
rect 512270 146956 512276 146968
rect 512328 146956 512334 147008
rect 211154 146888 211160 146940
rect 211212 146928 211218 146940
rect 280154 146928 280160 146940
rect 211212 146900 280160 146928
rect 211212 146888 211218 146900
rect 280154 146888 280160 146900
rect 280212 146888 280218 146940
rect 282454 146888 282460 146940
rect 282512 146928 282518 146940
rect 412726 146928 412732 146940
rect 282512 146900 412732 146928
rect 282512 146888 282518 146900
rect 412726 146888 412732 146900
rect 412784 146888 412790 146940
rect 485774 146888 485780 146940
rect 485832 146928 485838 146940
rect 562318 146928 562324 146940
rect 485832 146900 562324 146928
rect 485832 146888 485838 146900
rect 562318 146888 562324 146900
rect 562376 146888 562382 146940
rect 379514 146316 379520 146328
rect 378152 146288 379520 146316
rect 377306 146208 377312 146260
rect 377364 146248 377370 146260
rect 378152 146248 378180 146288
rect 379514 146276 379520 146288
rect 379572 146276 379578 146328
rect 377364 146220 378180 146248
rect 377364 146208 377370 146220
rect 169202 145528 169208 145580
rect 169260 145568 169266 145580
rect 215294 145568 215300 145580
rect 169260 145540 215300 145568
rect 169260 145528 169266 145540
rect 215294 145528 215300 145540
rect 215352 145528 215358 145580
rect 398466 144236 398472 144288
rect 398524 144276 398530 144288
rect 410518 144276 410524 144288
rect 398524 144248 410524 144276
rect 398524 144236 398530 144248
rect 410518 144236 410524 144248
rect 410576 144236 410582 144288
rect 189074 144168 189080 144220
rect 189132 144208 189138 144220
rect 580442 144208 580448 144220
rect 189132 144180 580448 144208
rect 189132 144168 189138 144180
rect 580442 144168 580448 144180
rect 580500 144168 580506 144220
rect 194594 143488 194600 143540
rect 194652 143528 194658 143540
rect 195054 143528 195060 143540
rect 194652 143500 195060 143528
rect 194652 143488 194658 143500
rect 195054 143488 195060 143500
rect 195112 143528 195118 143540
rect 418890 143528 418896 143540
rect 195112 143500 418896 143528
rect 195112 143488 195118 143500
rect 418890 143488 418896 143500
rect 418948 143488 418954 143540
rect 192570 143420 192576 143472
rect 192628 143460 192634 143472
rect 406010 143460 406016 143472
rect 192628 143432 406016 143460
rect 192628 143420 192634 143432
rect 406010 143420 406016 143432
rect 406068 143420 406074 143472
rect 188338 142876 188344 142928
rect 188396 142916 188402 142928
rect 195054 142916 195060 142928
rect 188396 142888 195060 142916
rect 188396 142876 188402 142888
rect 195054 142876 195060 142888
rect 195112 142876 195118 142928
rect 398558 142876 398564 142928
rect 398616 142916 398622 142928
rect 409414 142916 409420 142928
rect 398616 142888 409420 142916
rect 398616 142876 398622 142888
rect 409414 142876 409420 142888
rect 409472 142876 409478 142928
rect 417418 142876 417424 142928
rect 417476 142916 417482 142928
rect 454678 142916 454684 142928
rect 417476 142888 454684 142916
rect 417476 142876 417482 142888
rect 454678 142876 454684 142888
rect 454736 142876 454742 142928
rect 176194 142808 176200 142860
rect 176252 142848 176258 142860
rect 191834 142848 191840 142860
rect 176252 142820 191840 142848
rect 176252 142808 176258 142820
rect 191834 142808 191840 142820
rect 191892 142848 191898 142860
rect 192570 142848 192576 142860
rect 191892 142820 192576 142848
rect 191892 142808 191898 142820
rect 192570 142808 192576 142820
rect 192628 142808 192634 142860
rect 274266 142808 274272 142860
rect 274324 142848 274330 142860
rect 323578 142848 323584 142860
rect 274324 142820 323584 142848
rect 274324 142808 274330 142820
rect 323578 142808 323584 142820
rect 323636 142808 323642 142860
rect 376018 142808 376024 142860
rect 376076 142848 376082 142860
rect 377306 142848 377312 142860
rect 376076 142820 377312 142848
rect 376076 142808 376082 142820
rect 377306 142808 377312 142820
rect 377364 142808 377370 142860
rect 399386 142808 399392 142860
rect 399444 142848 399450 142860
rect 411530 142848 411536 142860
rect 399444 142820 411536 142848
rect 399444 142808 399450 142820
rect 411530 142808 411536 142820
rect 411588 142808 411594 142860
rect 418798 142808 418804 142860
rect 418856 142848 418862 142860
rect 479150 142848 479156 142860
rect 418856 142820 479156 142848
rect 418856 142808 418862 142820
rect 479150 142808 479156 142820
rect 479208 142808 479214 142860
rect 14 142672 20 142724
rect 72 142712 78 142724
rect 1302 142712 1308 142724
rect 72 142684 1308 142712
rect 72 142672 78 142684
rect 1302 142672 1308 142684
rect 1360 142672 1366 142724
rect 1302 142196 1308 142248
rect 1360 142236 1366 142248
rect 176194 142236 176200 142248
rect 1360 142208 176200 142236
rect 1360 142196 1366 142208
rect 176194 142196 176200 142208
rect 176252 142196 176258 142248
rect 1394 142128 1400 142180
rect 1452 142168 1458 142180
rect 188338 142168 188344 142180
rect 1452 142140 188344 142168
rect 1452 142128 1458 142140
rect 188338 142128 188344 142140
rect 188396 142128 188402 142180
rect 398650 141720 398656 141772
rect 398708 141760 398714 141772
rect 409506 141760 409512 141772
rect 398708 141732 409512 141760
rect 398708 141720 398714 141732
rect 409506 141720 409512 141732
rect 409564 141720 409570 141772
rect 394142 141652 394148 141704
rect 394200 141692 394206 141704
rect 404998 141692 405004 141704
rect 394200 141664 405004 141692
rect 394200 141652 394206 141664
rect 404998 141652 405004 141664
rect 405056 141652 405062 141704
rect 399294 141584 399300 141636
rect 399352 141624 399358 141636
rect 411622 141624 411628 141636
rect 399352 141596 411628 141624
rect 399352 141584 399358 141596
rect 411622 141584 411628 141596
rect 411680 141584 411686 141636
rect 438210 141584 438216 141636
rect 438268 141624 438274 141636
rect 509326 141624 509332 141636
rect 438268 141596 509332 141624
rect 438268 141584 438274 141596
rect 509326 141584 509332 141596
rect 509384 141584 509390 141636
rect 394234 141516 394240 141568
rect 394292 141556 394298 141568
rect 406378 141556 406384 141568
rect 394292 141528 406384 141556
rect 394292 141516 394298 141528
rect 406378 141516 406384 141528
rect 406436 141516 406442 141568
rect 438118 141516 438124 141568
rect 438176 141556 438182 141568
rect 509418 141556 509424 141568
rect 438176 141528 509424 141556
rect 438176 141516 438182 141528
rect 509418 141516 509424 141528
rect 509476 141516 509482 141568
rect 395798 141448 395804 141500
rect 395856 141488 395862 141500
rect 419534 141488 419540 141500
rect 395856 141460 419540 141488
rect 395856 141448 395862 141460
rect 419534 141448 419540 141460
rect 419592 141448 419598 141500
rect 435358 141448 435364 141500
rect 435416 141488 435422 141500
rect 510706 141488 510712 141500
rect 435416 141460 510712 141488
rect 435416 141448 435422 141460
rect 510706 141448 510712 141460
rect 510764 141448 510770 141500
rect 198734 141380 198740 141432
rect 198792 141420 198798 141432
rect 518158 141420 518164 141432
rect 198792 141392 518164 141420
rect 198792 141380 198798 141392
rect 518158 141380 518164 141392
rect 518216 141380 518222 141432
rect 168190 141040 168196 141092
rect 168248 141080 168254 141092
rect 173158 141080 173164 141092
rect 168248 141052 173164 141080
rect 168248 141040 168254 141052
rect 173158 141040 173164 141052
rect 173216 141040 173222 141092
rect 170122 140972 170128 141024
rect 170180 141012 170186 141024
rect 393774 141012 393780 141024
rect 170180 140984 393780 141012
rect 170180 140972 170186 140984
rect 393774 140972 393780 140984
rect 393832 141012 393838 141024
rect 394234 141012 394240 141024
rect 393832 140984 394240 141012
rect 393832 140972 393838 140984
rect 394234 140972 394240 140984
rect 394292 140972 394298 141024
rect 169662 140904 169668 140956
rect 169720 140944 169726 140956
rect 393866 140944 393872 140956
rect 169720 140916 393872 140944
rect 169720 140904 169726 140916
rect 393866 140904 393872 140916
rect 393924 140904 393930 140956
rect 169570 140836 169576 140888
rect 169628 140876 169634 140888
rect 394142 140876 394148 140888
rect 169628 140848 394148 140876
rect 169628 140836 169634 140848
rect 394142 140836 394148 140848
rect 394200 140836 394206 140888
rect 170030 140768 170036 140820
rect 170088 140808 170094 140820
rect 400214 140808 400220 140820
rect 170088 140780 400220 140808
rect 170088 140768 170094 140780
rect 400214 140768 400220 140780
rect 400272 140808 400278 140820
rect 401226 140808 401232 140820
rect 400272 140780 401232 140808
rect 400272 140768 400278 140780
rect 401226 140768 401232 140780
rect 401284 140768 401290 140820
rect 397914 140700 397920 140752
rect 397972 140740 397978 140752
rect 410150 140740 410156 140752
rect 397972 140712 410156 140740
rect 397972 140700 397978 140712
rect 410150 140700 410156 140712
rect 410208 140700 410214 140752
rect 394234 140604 394240 140616
rect 393286 140576 394240 140604
rect 169938 140292 169944 140344
rect 169996 140332 170002 140344
rect 393286 140332 393314 140576
rect 394234 140564 394240 140576
rect 394292 140604 394298 140616
rect 403618 140604 403624 140616
rect 394292 140576 403624 140604
rect 394292 140564 394298 140576
rect 403618 140564 403624 140576
rect 403676 140564 403682 140616
rect 169996 140304 393314 140332
rect 169996 140292 170002 140304
rect 398190 140292 398196 140344
rect 398248 140332 398254 140344
rect 410058 140332 410064 140344
rect 398248 140304 410064 140332
rect 398248 140292 398254 140304
rect 410058 140292 410064 140304
rect 410116 140292 410122 140344
rect 167546 140224 167552 140276
rect 167604 140264 167610 140276
rect 392670 140264 392676 140276
rect 167604 140236 392676 140264
rect 167604 140224 167610 140236
rect 392670 140224 392676 140236
rect 392728 140224 392734 140276
rect 398006 140224 398012 140276
rect 398064 140264 398070 140276
rect 409874 140264 409880 140276
rect 398064 140236 409880 140264
rect 398064 140224 398070 140236
rect 409874 140224 409880 140236
rect 409932 140224 409938 140276
rect 168374 140156 168380 140208
rect 168432 140196 168438 140208
rect 394142 140196 394148 140208
rect 168432 140168 394148 140196
rect 168432 140156 168438 140168
rect 394142 140156 394148 140168
rect 394200 140196 394206 140208
rect 407758 140196 407764 140208
rect 394200 140168 407764 140196
rect 394200 140156 394206 140168
rect 407758 140156 407764 140168
rect 407816 140156 407822 140208
rect 167454 140088 167460 140140
rect 167512 140128 167518 140140
rect 395430 140128 395436 140140
rect 167512 140100 395436 140128
rect 167512 140088 167518 140100
rect 395430 140088 395436 140100
rect 395488 140088 395494 140140
rect 398098 140088 398104 140140
rect 398156 140128 398162 140140
rect 409966 140128 409972 140140
rect 398156 140100 409972 140128
rect 398156 140088 398162 140100
rect 409966 140088 409972 140100
rect 410024 140088 410030 140140
rect 167822 140020 167828 140072
rect 167880 140060 167886 140072
rect 395522 140060 395528 140072
rect 167880 140032 395528 140060
rect 167880 140020 167886 140032
rect 395522 140020 395528 140032
rect 395580 140020 395586 140072
rect 396074 140020 396080 140072
rect 396132 140060 396138 140072
rect 396718 140060 396724 140072
rect 396132 140032 396724 140060
rect 396132 140020 396138 140032
rect 396718 140020 396724 140032
rect 396776 140020 396782 140072
rect 398282 140020 398288 140072
rect 398340 140060 398346 140072
rect 410242 140060 410248 140072
rect 398340 140032 410248 140060
rect 398340 140020 398346 140032
rect 410242 140020 410248 140032
rect 410300 140020 410306 140072
rect 169294 139952 169300 140004
rect 169352 139992 169358 140004
rect 396534 139992 396540 140004
rect 169352 139964 396540 139992
rect 169352 139952 169358 139964
rect 396534 139952 396540 139964
rect 396592 139992 396598 140004
rect 403802 139992 403808 140004
rect 396592 139964 403808 139992
rect 396592 139952 396598 139964
rect 403802 139952 403808 139964
rect 403860 139952 403866 140004
rect 168006 139884 168012 139936
rect 168064 139924 168070 139936
rect 395154 139924 395160 139936
rect 168064 139896 395160 139924
rect 168064 139884 168070 139896
rect 395154 139884 395160 139896
rect 395212 139924 395218 139936
rect 395614 139924 395620 139936
rect 395212 139896 395620 139924
rect 395212 139884 395218 139896
rect 395614 139884 395620 139896
rect 395672 139884 395678 139936
rect 396810 139884 396816 139936
rect 396868 139924 396874 139936
rect 403710 139924 403716 139936
rect 396868 139896 403716 139924
rect 396868 139884 396874 139896
rect 403710 139884 403716 139896
rect 403768 139884 403774 139936
rect 167914 139816 167920 139868
rect 167972 139856 167978 139868
rect 396074 139856 396080 139868
rect 167972 139828 396080 139856
rect 167972 139816 167978 139828
rect 396074 139816 396080 139828
rect 396132 139816 396138 139868
rect 169386 139748 169392 139800
rect 169444 139788 169450 139800
rect 398190 139788 398196 139800
rect 169444 139760 398196 139788
rect 169444 139748 169450 139760
rect 398190 139748 398196 139760
rect 398248 139748 398254 139800
rect 398834 139748 398840 139800
rect 398892 139788 398898 139800
rect 400122 139788 400128 139800
rect 398892 139760 400128 139788
rect 398892 139748 398898 139760
rect 400122 139748 400128 139760
rect 400180 139748 400186 139800
rect 169110 139680 169116 139732
rect 169168 139720 169174 139732
rect 398006 139720 398012 139732
rect 169168 139692 398012 139720
rect 169168 139680 169174 139692
rect 398006 139680 398012 139692
rect 398064 139680 398070 139732
rect 168282 139612 168288 139664
rect 168340 139652 168346 139664
rect 398098 139652 398104 139664
rect 168340 139624 398104 139652
rect 168340 139612 168346 139624
rect 398098 139612 398104 139624
rect 398156 139612 398162 139664
rect 166902 139544 166908 139596
rect 166960 139584 166966 139596
rect 396626 139584 396632 139596
rect 166960 139556 396632 139584
rect 166960 139544 166966 139556
rect 396626 139544 396632 139556
rect 396684 139584 396690 139596
rect 401134 139584 401140 139596
rect 396684 139556 401140 139584
rect 396684 139544 396690 139556
rect 401134 139544 401140 139556
rect 401192 139544 401198 139596
rect 165522 139476 165528 139528
rect 165580 139516 165586 139528
rect 396810 139516 396816 139528
rect 165580 139488 396816 139516
rect 165580 139476 165586 139488
rect 396810 139476 396816 139488
rect 396868 139476 396874 139528
rect 167638 139408 167644 139460
rect 167696 139448 167702 139460
rect 398834 139448 398840 139460
rect 167696 139420 398840 139448
rect 167696 139408 167702 139420
rect 398834 139408 398840 139420
rect 398892 139408 398898 139460
rect 400582 137844 400588 137896
rect 400640 137884 400646 137896
rect 401042 137884 401048 137896
rect 400640 137856 401048 137884
rect 400640 137844 400646 137856
rect 401042 137844 401048 137856
rect 401100 137844 401106 137896
rect 167546 136076 167552 136128
rect 167604 136116 167610 136128
rect 168006 136116 168012 136128
rect 167604 136088 168012 136116
rect 167604 136076 167610 136088
rect 168006 136076 168012 136088
rect 168064 136076 168070 136128
rect 167546 135940 167552 135992
rect 167604 135980 167610 135992
rect 168374 135980 168380 135992
rect 167604 135952 168380 135980
rect 167604 135940 167610 135952
rect 168374 135940 168380 135952
rect 168432 135940 168438 135992
rect 305638 135192 305644 135244
rect 305696 135232 305702 135244
rect 397454 135232 397460 135244
rect 305696 135204 397460 135232
rect 305696 135192 305702 135204
rect 397454 135192 397460 135204
rect 397512 135192 397518 135244
rect 167822 134172 167828 134224
rect 167880 134212 167886 134224
rect 168190 134212 168196 134224
rect 167880 134184 168196 134212
rect 167880 134172 167886 134184
rect 168190 134172 168196 134184
rect 168248 134172 168254 134224
rect 167546 134036 167552 134088
rect 167604 134076 167610 134088
rect 167822 134076 167828 134088
rect 167604 134048 167828 134076
rect 167604 134036 167610 134048
rect 167822 134036 167828 134048
rect 167880 134036 167886 134088
rect 309778 133832 309784 133884
rect 309836 133872 309842 133884
rect 397454 133872 397460 133884
rect 309836 133844 397460 133872
rect 309836 133832 309842 133844
rect 397454 133832 397460 133844
rect 397512 133832 397518 133884
rect 347774 129684 347780 129736
rect 347832 129724 347838 129736
rect 397454 129724 397460 129736
rect 347832 129696 397460 129724
rect 347832 129684 347838 129696
rect 397454 129684 397460 129696
rect 397512 129684 397518 129736
rect 393866 128324 393872 128376
rect 393924 128364 393930 128376
rect 398374 128364 398380 128376
rect 393924 128336 398380 128364
rect 393924 128324 393930 128336
rect 398374 128324 398380 128336
rect 398432 128324 398438 128376
rect 562318 126896 562324 126948
rect 562376 126936 562382 126948
rect 579706 126936 579712 126948
rect 562376 126908 579712 126936
rect 562376 126896 562382 126908
rect 579706 126896 579712 126908
rect 579764 126896 579770 126948
rect 375006 126624 375012 126676
rect 375064 126664 375070 126676
rect 376018 126664 376024 126676
rect 375064 126636 376024 126664
rect 375064 126624 375070 126636
rect 376018 126624 376024 126636
rect 376076 126624 376082 126676
rect 287054 125536 287060 125588
rect 287112 125576 287118 125588
rect 397454 125576 397460 125588
rect 287112 125548 397460 125576
rect 287112 125536 287118 125548
rect 397454 125536 397460 125548
rect 397512 125536 397518 125588
rect 372614 124176 372620 124228
rect 372672 124216 372678 124228
rect 375006 124216 375012 124228
rect 372672 124188 375012 124216
rect 372672 124176 372678 124188
rect 375006 124176 375012 124188
rect 375064 124176 375070 124228
rect 349798 124108 349804 124160
rect 349856 124148 349862 124160
rect 397454 124148 397460 124160
rect 349856 124120 397460 124148
rect 349856 124108 349862 124120
rect 397454 124108 397460 124120
rect 397512 124108 397518 124160
rect 392762 123428 392768 123480
rect 392820 123468 392826 123480
rect 397914 123468 397920 123480
rect 392820 123440 397920 123468
rect 392820 123428 392826 123440
rect 397914 123428 397920 123440
rect 397972 123428 397978 123480
rect 371878 123088 371884 123140
rect 371936 123128 371942 123140
rect 372614 123128 372620 123140
rect 371936 123100 372620 123128
rect 371936 123088 371942 123100
rect 372614 123088 372620 123100
rect 372672 123088 372678 123140
rect 400582 121388 400588 121440
rect 400640 121428 400646 121440
rect 400950 121428 400956 121440
rect 400640 121400 400956 121428
rect 400640 121388 400646 121400
rect 400950 121388 400956 121400
rect 401008 121388 401014 121440
rect 286318 120028 286324 120080
rect 286376 120068 286382 120080
rect 397454 120068 397460 120080
rect 286376 120040 397460 120068
rect 286376 120028 286382 120040
rect 397454 120028 397460 120040
rect 397512 120028 397518 120080
rect 395614 118668 395620 118720
rect 395672 118708 395678 118720
rect 396074 118708 396080 118720
rect 395672 118680 396080 118708
rect 395672 118668 395678 118680
rect 396074 118668 396080 118680
rect 396132 118668 396138 118720
rect 396626 118600 396632 118652
rect 396684 118640 396690 118652
rect 398098 118640 398104 118652
rect 396684 118612 398104 118640
rect 396684 118600 396690 118612
rect 398098 118600 398104 118612
rect 398156 118600 398162 118652
rect 551278 113092 551284 113144
rect 551336 113132 551342 113144
rect 579706 113132 579712 113144
rect 551336 113104 579712 113132
rect 551336 113092 551342 113104
rect 579706 113092 579712 113104
rect 579764 113092 579770 113144
rect 396534 113024 396540 113076
rect 396592 113064 396598 113076
rect 397546 113064 397552 113076
rect 396592 113036 397552 113064
rect 396592 113024 396598 113036
rect 397546 113024 397552 113036
rect 397604 113024 397610 113076
rect 395154 106224 395160 106276
rect 395212 106264 395218 106276
rect 399570 106264 399576 106276
rect 395212 106236 399576 106264
rect 395212 106224 395218 106236
rect 399570 106224 399576 106236
rect 399628 106224 399634 106276
rect 393774 104796 393780 104848
rect 393832 104836 393838 104848
rect 397454 104836 397460 104848
rect 393832 104808 397460 104836
rect 393832 104796 393838 104808
rect 397454 104796 397460 104808
rect 397512 104796 397518 104848
rect 394050 102076 394056 102128
rect 394108 102116 394114 102128
rect 397454 102116 397460 102128
rect 394108 102088 397460 102116
rect 394108 102076 394114 102088
rect 397454 102076 397460 102088
rect 397512 102076 397518 102128
rect 394142 99288 394148 99340
rect 394200 99328 394206 99340
rect 397454 99328 397460 99340
rect 394200 99300 397460 99328
rect 394200 99288 394206 99300
rect 397454 99288 397460 99300
rect 397512 99288 397518 99340
rect 371878 98036 371884 98048
rect 368492 98008 371884 98036
rect 367738 97928 367744 97980
rect 367796 97968 367802 97980
rect 368492 97968 368520 98008
rect 371878 97996 371884 98008
rect 371936 97996 371942 98048
rect 367796 97940 368520 97968
rect 367796 97928 367802 97940
rect 395430 97928 395436 97980
rect 395488 97968 395494 97980
rect 398190 97968 398196 97980
rect 395488 97940 398196 97968
rect 395488 97928 395494 97940
rect 398190 97928 398196 97940
rect 398248 97928 398254 97980
rect 165522 96568 165528 96620
rect 165580 96608 165586 96620
rect 166994 96608 167000 96620
rect 165580 96580 167000 96608
rect 165580 96568 165586 96580
rect 166994 96568 167000 96580
rect 167052 96568 167058 96620
rect 394234 95140 394240 95192
rect 394292 95180 394298 95192
rect 397454 95180 397460 95192
rect 394292 95152 397460 95180
rect 394292 95140 394298 95152
rect 397454 95140 397460 95152
rect 397512 95140 397518 95192
rect 392578 92420 392584 92472
rect 392636 92460 392642 92472
rect 397454 92460 397460 92472
rect 392636 92432 397460 92460
rect 392636 92420 392642 92432
rect 397454 92420 397460 92432
rect 397512 92420 397518 92472
rect 364978 91060 364984 91112
rect 365036 91100 365042 91112
rect 367738 91100 367744 91112
rect 365036 91072 367744 91100
rect 365036 91060 365042 91072
rect 367738 91060 367744 91072
rect 367796 91060 367802 91112
rect 395614 90992 395620 91044
rect 395672 91032 395678 91044
rect 397914 91032 397920 91044
rect 395672 91004 397920 91032
rect 395672 90992 395678 91004
rect 397914 90992 397920 91004
rect 397972 90992 397978 91044
rect 392670 89632 392676 89684
rect 392728 89672 392734 89684
rect 397454 89672 397460 89684
rect 392728 89644 397460 89672
rect 392728 89632 392734 89644
rect 397454 89632 397460 89644
rect 397512 89632 397518 89684
rect 395706 88272 395712 88324
rect 395764 88312 395770 88324
rect 398834 88312 398840 88324
rect 395764 88284 398840 88312
rect 395764 88272 395770 88284
rect 398834 88272 398840 88284
rect 398892 88272 398898 88324
rect 395522 86912 395528 86964
rect 395580 86952 395586 86964
rect 397730 86952 397736 86964
rect 395580 86924 397736 86952
rect 395580 86912 395586 86924
rect 397730 86912 397736 86924
rect 397788 86912 397794 86964
rect 544378 86912 544384 86964
rect 544436 86952 544442 86964
rect 579982 86952 579988 86964
rect 544436 86924 579988 86952
rect 544436 86912 544442 86924
rect 579982 86912 579988 86924
rect 580040 86912 580046 86964
rect 395246 85484 395252 85536
rect 395304 85524 395310 85536
rect 397546 85524 397552 85536
rect 395304 85496 397552 85524
rect 395304 85484 395310 85496
rect 397546 85484 397552 85496
rect 397604 85484 397610 85536
rect 360194 83988 360200 84040
rect 360252 84028 360258 84040
rect 364978 84028 364984 84040
rect 360252 84000 364984 84028
rect 360252 83988 360258 84000
rect 364978 83988 364984 84000
rect 365036 83988 365042 84040
rect 392578 82084 392584 82136
rect 392636 82124 392642 82136
rect 392946 82124 392952 82136
rect 392636 82096 392952 82124
rect 392636 82084 392642 82096
rect 392946 82084 392952 82096
rect 393004 82124 393010 82136
rect 397454 82124 397460 82136
rect 393004 82096 397460 82124
rect 393004 82084 393010 82096
rect 397454 82084 397460 82096
rect 397512 82084 397518 82136
rect 356698 81404 356704 81456
rect 356756 81444 356762 81456
rect 360194 81444 360200 81456
rect 356756 81416 360200 81444
rect 356756 81404 356762 81416
rect 360194 81404 360200 81416
rect 360252 81404 360258 81456
rect 395890 79636 395896 79688
rect 395948 79676 395954 79688
rect 398190 79676 398196 79688
rect 395948 79648 398196 79676
rect 395948 79636 395954 79648
rect 398190 79636 398196 79648
rect 398248 79636 398254 79688
rect 394326 78548 394332 78600
rect 394384 78588 394390 78600
rect 397454 78588 397460 78600
rect 394384 78560 397460 78588
rect 394384 78548 394390 78560
rect 397454 78548 397460 78560
rect 397512 78548 397518 78600
rect 396902 75216 396908 75268
rect 396960 75256 396966 75268
rect 398098 75256 398104 75268
rect 396960 75228 398104 75256
rect 396960 75216 396966 75228
rect 398098 75216 398104 75228
rect 398156 75216 398162 75268
rect 395430 71816 395436 71868
rect 395488 71856 395494 71868
rect 397914 71856 397920 71868
rect 395488 71828 397920 71856
rect 395488 71816 395494 71828
rect 397914 71816 397920 71828
rect 397972 71816 397978 71868
rect 355318 68280 355324 68332
rect 355376 68320 355382 68332
rect 356698 68320 356704 68332
rect 355376 68292 356704 68320
rect 355376 68280 355382 68292
rect 356698 68280 356704 68292
rect 356756 68280 356762 68332
rect 392670 66852 392676 66904
rect 392728 66892 392734 66904
rect 393038 66892 393044 66904
rect 392728 66864 393044 66892
rect 392728 66852 392734 66864
rect 393038 66852 393044 66864
rect 393096 66892 393102 66904
rect 397454 66892 397460 66904
rect 393096 66864 397460 66892
rect 393096 66852 393102 66864
rect 397454 66852 397460 66864
rect 397512 66852 397518 66904
rect 165522 64948 165528 65000
rect 165580 64988 165586 65000
rect 168282 64988 168288 65000
rect 165580 64960 168288 64988
rect 165580 64948 165586 64960
rect 168282 64948 168288 64960
rect 168340 64948 168346 65000
rect 280798 57196 280804 57248
rect 280856 57236 280862 57248
rect 395982 57236 395988 57248
rect 280856 57208 395988 57236
rect 280856 57196 280862 57208
rect 395982 57196 395988 57208
rect 396040 57236 396046 57248
rect 397454 57236 397460 57248
rect 396040 57208 397460 57236
rect 396040 57196 396046 57208
rect 397454 57196 397460 57208
rect 397512 57196 397518 57248
rect 355318 56624 355324 56636
rect 354646 56596 355324 56624
rect 351914 56516 351920 56568
rect 351972 56556 351978 56568
rect 354646 56556 354674 56596
rect 355318 56584 355324 56596
rect 355376 56584 355382 56636
rect 351972 56528 354674 56556
rect 351972 56516 351978 56528
rect 398006 56176 398012 56228
rect 398064 56216 398070 56228
rect 399110 56216 399116 56228
rect 398064 56188 399116 56216
rect 398064 56176 398070 56188
rect 399110 56176 399116 56188
rect 399168 56176 399174 56228
rect 282178 54476 282184 54528
rect 282236 54516 282242 54528
rect 396994 54516 397000 54528
rect 282236 54488 397000 54516
rect 282236 54476 282242 54488
rect 396994 54476 397000 54488
rect 397052 54476 397058 54528
rect 347498 53796 347504 53848
rect 347556 53836 347562 53848
rect 351914 53836 351920 53848
rect 347556 53808 351920 53836
rect 347556 53796 347562 53808
rect 351914 53796 351920 53808
rect 351972 53796 351978 53848
rect 282822 51008 282828 51060
rect 282880 51048 282886 51060
rect 347498 51048 347504 51060
rect 282880 51020 347504 51048
rect 282880 51008 282886 51020
rect 347498 51008 347504 51020
rect 347556 51008 347562 51060
rect 279418 48968 279424 49020
rect 279476 49008 279482 49020
rect 397086 49008 397092 49020
rect 279476 48980 397092 49008
rect 279476 48968 279482 48980
rect 397086 48968 397092 48980
rect 397144 49008 397150 49020
rect 397454 49008 397460 49020
rect 397144 48980 397460 49008
rect 397144 48968 397150 48980
rect 397454 48968 397460 48980
rect 397512 48968 397518 49020
rect 282270 47540 282276 47592
rect 282328 47580 282334 47592
rect 397454 47580 397460 47592
rect 282328 47552 397460 47580
rect 282328 47540 282334 47552
rect 397454 47540 397460 47552
rect 397512 47540 397518 47592
rect 398742 46860 398748 46912
rect 398800 46900 398806 46912
rect 399018 46900 399024 46912
rect 398800 46872 399024 46900
rect 398800 46860 398806 46872
rect 399018 46860 399024 46872
rect 399076 46860 399082 46912
rect 518158 46860 518164 46912
rect 518216 46900 518222 46912
rect 580166 46900 580172 46912
rect 518216 46872 580172 46900
rect 518216 46860 518222 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 168098 44140 168104 44192
rect 168156 44180 168162 44192
rect 169018 44180 169024 44192
rect 168156 44152 169024 44180
rect 168156 44140 168162 44152
rect 169018 44140 169024 44152
rect 169076 44140 169082 44192
rect 280890 43392 280896 43444
rect 280948 43432 280954 43444
rect 397178 43432 397184 43444
rect 280948 43404 397184 43432
rect 280948 43392 280954 43404
rect 397178 43392 397184 43404
rect 397236 43392 397242 43444
rect 167822 42032 167828 42084
rect 167880 42072 167886 42084
rect 169202 42072 169208 42084
rect 167880 42044 169208 42072
rect 167880 42032 167886 42044
rect 169202 42032 169208 42044
rect 169260 42032 169266 42084
rect 167730 41692 167736 41744
rect 167788 41732 167794 41744
rect 169110 41732 169116 41744
rect 167788 41704 169116 41732
rect 167788 41692 167794 41704
rect 169110 41692 169116 41704
rect 169168 41692 169174 41744
rect 279510 41420 279516 41472
rect 279568 41460 279574 41472
rect 397454 41460 397460 41472
rect 279568 41432 397460 41460
rect 279568 41420 279574 41432
rect 397454 41420 397460 41432
rect 397512 41420 397518 41472
rect 280982 40672 280988 40724
rect 281040 40712 281046 40724
rect 394510 40712 394516 40724
rect 281040 40684 394516 40712
rect 281040 40672 281046 40684
rect 394510 40672 394516 40684
rect 394568 40712 394574 40724
rect 397454 40712 397460 40724
rect 394568 40684 397460 40712
rect 394568 40672 394574 40684
rect 397454 40672 397460 40684
rect 397512 40672 397518 40724
rect 397730 40672 397736 40724
rect 397788 40712 397794 40724
rect 398742 40712 398748 40724
rect 397788 40684 398748 40712
rect 397788 40672 397794 40684
rect 398742 40672 398748 40684
rect 398800 40672 398806 40724
rect 168006 39992 168012 40044
rect 168064 40032 168070 40044
rect 169294 40032 169300 40044
rect 168064 40004 169300 40032
rect 168064 39992 168070 40004
rect 169294 39992 169300 40004
rect 169352 39992 169358 40044
rect 281074 39312 281080 39364
rect 281132 39352 281138 39364
rect 397270 39352 397276 39364
rect 281132 39324 397276 39352
rect 281132 39312 281138 39324
rect 397270 39312 397276 39324
rect 397328 39352 397334 39364
rect 397454 39352 397460 39364
rect 397328 39324 397460 39352
rect 397328 39312 397334 39324
rect 397454 39312 397460 39324
rect 397512 39312 397518 39364
rect 278958 37272 278964 37324
rect 279016 37312 279022 37324
rect 397546 37312 397552 37324
rect 279016 37284 397552 37312
rect 279016 37272 279022 37284
rect 397546 37272 397552 37284
rect 397604 37272 397610 37324
rect 167914 37204 167920 37256
rect 167972 37244 167978 37256
rect 168926 37244 168932 37256
rect 167972 37216 168932 37244
rect 167972 37204 167978 37216
rect 168926 37204 168932 37216
rect 168984 37204 168990 37256
rect 509234 37204 509240 37256
rect 509292 37244 509298 37256
rect 509510 37244 509516 37256
rect 509292 37216 509516 37244
rect 509292 37204 509298 37216
rect 509510 37204 509516 37216
rect 509568 37204 509574 37256
rect 281166 36524 281172 36576
rect 281224 36564 281230 36576
rect 335354 36564 335360 36576
rect 281224 36536 335360 36564
rect 281224 36524 281230 36536
rect 335354 36524 335360 36536
rect 335412 36524 335418 36576
rect 279970 34484 279976 34536
rect 280028 34524 280034 34536
rect 399754 34524 399760 34536
rect 280028 34496 399760 34524
rect 280028 34484 280034 34496
rect 399754 34484 399760 34496
rect 399812 34484 399818 34536
rect 168926 33464 168932 33516
rect 168984 33504 168990 33516
rect 169570 33504 169576 33516
rect 168984 33476 169576 33504
rect 168984 33464 168990 33476
rect 169570 33464 169576 33476
rect 169628 33464 169634 33516
rect 168098 33260 168104 33312
rect 168156 33300 168162 33312
rect 169662 33300 169668 33312
rect 168156 33272 169668 33300
rect 168156 33260 168162 33272
rect 169662 33260 169668 33272
rect 169720 33260 169726 33312
rect 279326 32376 279332 32428
rect 279384 32416 279390 32428
rect 394602 32416 394608 32428
rect 279384 32388 394608 32416
rect 279384 32376 279390 32388
rect 394602 32376 394608 32388
rect 394660 32416 394666 32428
rect 397454 32416 397460 32428
rect 394660 32388 397460 32416
rect 394660 32376 394666 32388
rect 397454 32376 397460 32388
rect 397512 32376 397518 32428
rect 165522 31696 165528 31748
rect 165580 31736 165586 31748
rect 398466 31736 398472 31748
rect 165580 31708 398472 31736
rect 165580 31696 165586 31708
rect 398466 31696 398472 31708
rect 398524 31696 398530 31748
rect 169386 31628 169392 31680
rect 169444 31668 169450 31680
rect 398650 31668 398656 31680
rect 169444 31640 398656 31668
rect 169444 31628 169450 31640
rect 398650 31628 398656 31640
rect 398708 31628 398714 31680
rect 169478 31560 169484 31612
rect 169536 31600 169542 31612
rect 398558 31600 398564 31612
rect 169536 31572 398564 31600
rect 169536 31560 169542 31572
rect 398558 31560 398564 31572
rect 398616 31560 398622 31612
rect 391934 31492 391940 31544
rect 391992 31532 391998 31544
rect 393222 31532 393228 31544
rect 391992 31504 393228 31532
rect 391992 31492 391998 31504
rect 393222 31492 393228 31504
rect 393280 31532 393286 31544
rect 397454 31532 397460 31544
rect 393280 31504 397460 31532
rect 393280 31492 393286 31504
rect 397454 31492 397460 31504
rect 397512 31492 397518 31544
rect 280062 31016 280068 31068
rect 280120 31056 280126 31068
rect 391934 31056 391940 31068
rect 280120 31028 391940 31056
rect 280120 31016 280126 31028
rect 391934 31016 391940 31028
rect 391992 31016 391998 31068
rect 169662 30268 169668 30320
rect 169720 30308 169726 30320
rect 398098 30308 398104 30320
rect 169720 30280 398104 30308
rect 169720 30268 169726 30280
rect 398098 30268 398104 30280
rect 398156 30268 398162 30320
rect 169938 30200 169944 30252
rect 169996 30240 170002 30252
rect 397730 30240 397736 30252
rect 169996 30212 397736 30240
rect 169996 30200 170002 30212
rect 397730 30200 397736 30212
rect 397788 30200 397794 30252
rect 169846 30132 169852 30184
rect 169904 30172 169910 30184
rect 397914 30172 397920 30184
rect 169904 30144 397920 30172
rect 169904 30132 169910 30144
rect 397914 30132 397920 30144
rect 397972 30132 397978 30184
rect 169018 30064 169024 30116
rect 169076 30104 169082 30116
rect 392578 30104 392584 30116
rect 169076 30076 392584 30104
rect 169076 30064 169082 30076
rect 392578 30064 392584 30076
rect 392636 30064 392642 30116
rect 168006 29996 168012 30048
rect 168064 30036 168070 30048
rect 281074 30036 281080 30048
rect 168064 30008 281080 30036
rect 168064 29996 168070 30008
rect 281074 29996 281080 30008
rect 281132 29996 281138 30048
rect 167178 29928 167184 29980
rect 167236 29968 167242 29980
rect 280890 29968 280896 29980
rect 167236 29940 280896 29968
rect 167236 29928 167242 29940
rect 280890 29928 280896 29940
rect 280948 29928 280954 29980
rect 168190 29860 168196 29912
rect 168248 29900 168254 29912
rect 278958 29900 278964 29912
rect 168248 29872 278964 29900
rect 168248 29860 168254 29872
rect 278958 29860 278964 29872
rect 279016 29860 279022 29912
rect 167822 29792 167828 29844
rect 167880 29832 167886 29844
rect 279510 29832 279516 29844
rect 167880 29804 279516 29832
rect 167880 29792 167886 29804
rect 279510 29792 279516 29804
rect 279568 29792 279574 29844
rect 170398 29724 170404 29776
rect 170456 29764 170462 29776
rect 280062 29764 280068 29776
rect 170456 29736 280068 29764
rect 170456 29724 170462 29736
rect 280062 29724 280068 29736
rect 280120 29724 280126 29776
rect 168282 29656 168288 29708
rect 168340 29696 168346 29708
rect 279970 29696 279976 29708
rect 168340 29668 279976 29696
rect 168340 29656 168346 29668
rect 279970 29656 279976 29668
rect 280028 29656 280034 29708
rect 167546 29588 167552 29640
rect 167604 29628 167610 29640
rect 279418 29628 279424 29640
rect 167604 29600 279424 29628
rect 167604 29588 167610 29600
rect 279418 29588 279424 29600
rect 279476 29588 279482 29640
rect 446858 29248 446864 29300
rect 446916 29288 446922 29300
rect 522298 29288 522304 29300
rect 446916 29260 522304 29288
rect 446916 29248 446922 29260
rect 522298 29248 522304 29260
rect 522356 29248 522362 29300
rect 438394 29180 438400 29232
rect 438452 29220 438458 29232
rect 520918 29220 520924 29232
rect 438452 29192 520924 29220
rect 438452 29180 438458 29192
rect 520918 29180 520924 29192
rect 520976 29180 520982 29232
rect 208302 29112 208308 29164
rect 208360 29152 208366 29164
rect 289078 29152 289084 29164
rect 208360 29124 289084 29152
rect 208360 29112 208366 29124
rect 289078 29112 289084 29124
rect 289136 29112 289142 29164
rect 429930 29112 429936 29164
rect 429988 29152 429994 29164
rect 560938 29152 560944 29164
rect 429988 29124 560944 29152
rect 429988 29112 429994 29124
rect 560938 29112 560944 29124
rect 560996 29112 561002 29164
rect 216490 29044 216496 29096
rect 216548 29084 216554 29096
rect 519538 29084 519544 29096
rect 216548 29056 519544 29084
rect 216548 29044 216554 29056
rect 519538 29044 519544 29056
rect 519596 29044 519602 29096
rect 183002 28976 183008 29028
rect 183060 29016 183066 29028
rect 515398 29016 515404 29028
rect 183060 28988 515404 29016
rect 183060 28976 183066 28988
rect 515398 28976 515404 28988
rect 515456 28976 515462 29028
rect 169110 28908 169116 28960
rect 169168 28948 169174 28960
rect 398374 28948 398380 28960
rect 169168 28920 398380 28948
rect 169168 28908 169174 28920
rect 398374 28908 398380 28920
rect 398432 28908 398438 28960
rect 506106 28908 506112 28960
rect 506164 28948 506170 28960
rect 510706 28948 510712 28960
rect 506164 28920 510712 28948
rect 506164 28908 506170 28920
rect 510706 28908 510712 28920
rect 510764 28908 510770 28960
rect 167270 28840 167276 28892
rect 167328 28880 167334 28892
rect 398190 28880 398196 28892
rect 167328 28852 398196 28880
rect 167328 28840 167334 28852
rect 398190 28840 398196 28852
rect 398248 28840 398254 28892
rect 497642 28840 497648 28892
rect 497700 28880 497706 28892
rect 509418 28880 509424 28892
rect 497700 28852 509424 28880
rect 497700 28840 497706 28852
rect 509418 28840 509424 28852
rect 509476 28840 509482 28892
rect 169570 28772 169576 28824
rect 169628 28812 169634 28824
rect 399202 28812 399208 28824
rect 169628 28784 399208 28812
rect 169628 28772 169634 28784
rect 399202 28772 399208 28784
rect 399260 28772 399266 28824
rect 413002 28772 413008 28824
rect 413060 28812 413066 28824
rect 554038 28812 554044 28824
rect 413060 28784 554044 28812
rect 413060 28772 413066 28784
rect 554038 28772 554044 28784
rect 554096 28772 554102 28824
rect 168834 28704 168840 28756
rect 168892 28744 168898 28756
rect 398282 28744 398288 28756
rect 168892 28716 398288 28744
rect 168892 28704 168898 28716
rect 398282 28704 398288 28716
rect 398340 28704 398346 28756
rect 421466 28704 421472 28756
rect 421524 28744 421530 28756
rect 549898 28744 549904 28756
rect 421524 28716 549904 28744
rect 421524 28704 421530 28716
rect 549898 28704 549904 28716
rect 549956 28704 549962 28756
rect 395338 28636 395344 28688
rect 395396 28676 395402 28688
rect 480346 28676 480352 28688
rect 395396 28648 480352 28676
rect 395396 28636 395402 28648
rect 480346 28636 480352 28648
rect 480404 28636 480410 28688
rect 489178 28636 489184 28688
rect 489236 28676 489242 28688
rect 509326 28676 509332 28688
rect 489236 28648 509332 28676
rect 489236 28636 489242 28648
rect 509326 28636 509332 28648
rect 509384 28636 509390 28688
rect 395798 28568 395804 28620
rect 395856 28608 395862 28620
rect 463142 28608 463148 28620
rect 395856 28580 463148 28608
rect 395856 28568 395862 28580
rect 463142 28568 463148 28580
rect 463200 28568 463206 28620
rect 169294 28500 169300 28552
rect 169352 28540 169358 28552
rect 396718 28540 396724 28552
rect 169352 28512 396724 28540
rect 169352 28500 169358 28512
rect 396718 28500 396724 28512
rect 396776 28500 396782 28552
rect 404170 28500 404176 28552
rect 404228 28540 404234 28552
rect 558178 28540 558184 28552
rect 404228 28512 558184 28540
rect 404228 28500 404234 28512
rect 558178 28500 558184 28512
rect 558236 28500 558242 28552
rect 169202 28432 169208 28484
rect 169260 28472 169266 28484
rect 395430 28472 395436 28484
rect 169260 28444 395436 28472
rect 169260 28432 169266 28444
rect 395430 28432 395436 28444
rect 395488 28432 395494 28484
rect 169754 28364 169760 28416
rect 169812 28404 169818 28416
rect 392670 28404 392676 28416
rect 169812 28376 392676 28404
rect 169812 28364 169818 28376
rect 392670 28364 392676 28376
rect 392728 28364 392734 28416
rect 28902 28296 28908 28348
rect 28960 28336 28966 28348
rect 224954 28336 224960 28348
rect 28960 28308 224960 28336
rect 28960 28296 28966 28308
rect 224954 28296 224960 28308
rect 225012 28296 225018 28348
rect 250714 28296 250720 28348
rect 250772 28336 250778 28348
rect 281166 28336 281172 28348
rect 250772 28308 281172 28336
rect 250772 28296 250778 28308
rect 281166 28296 281172 28308
rect 281224 28296 281230 28348
rect 307754 28296 307760 28348
rect 307812 28336 307818 28348
rect 472066 28336 472072 28348
rect 307812 28308 472072 28336
rect 307812 28296 307818 28308
rect 472066 28296 472072 28308
rect 472124 28296 472130 28348
rect 259178 28228 259184 28280
rect 259236 28268 259242 28280
rect 389818 28268 389824 28280
rect 259236 28240 389824 28268
rect 259236 28228 259242 28240
rect 389818 28228 389824 28240
rect 389876 28228 389882 28280
rect 167362 28160 167368 28212
rect 167420 28200 167426 28212
rect 282178 28200 282184 28212
rect 167420 28172 282184 28200
rect 167420 28160 167426 28172
rect 282178 28160 282184 28172
rect 282236 28160 282242 28212
rect 167454 28092 167460 28144
rect 167512 28132 167518 28144
rect 282270 28132 282276 28144
rect 167512 28104 282276 28132
rect 167512 28092 167518 28104
rect 282270 28092 282276 28104
rect 282328 28092 282334 28144
rect 171042 28024 171048 28076
rect 171100 28064 171106 28076
rect 266998 28064 267004 28076
rect 171100 28036 267004 28064
rect 171100 28024 171106 28036
rect 266998 28024 267004 28036
rect 267056 28024 267062 28076
rect 275922 28024 275928 28076
rect 275980 28064 275986 28076
rect 319438 28064 319444 28076
rect 275980 28036 319444 28064
rect 275980 28024 275986 28036
rect 319438 28024 319444 28036
rect 319496 28024 319502 28076
rect 174538 27956 174544 28008
rect 174596 27996 174602 28008
rect 555418 27996 555424 28008
rect 174596 27968 555424 27996
rect 174596 27956 174602 27968
rect 555418 27956 555424 27968
rect 555476 27956 555482 28008
rect 168926 27888 168932 27940
rect 168984 27928 168990 27940
rect 398006 27928 398012 27940
rect 168984 27900 398012 27928
rect 168984 27888 168990 27900
rect 398006 27888 398012 27900
rect 398064 27888 398070 27940
rect 284938 6808 284944 6860
rect 284996 6848 285002 6860
rect 580166 6848 580172 6860
rect 284996 6820 580172 6848
rect 284996 6808 285002 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
<< via1 >>
rect 242900 536800 242952 536852
rect 396632 536800 396684 536852
rect 237380 535440 237432 535492
rect 396632 535440 396684 535492
rect 231860 532788 231912 532840
rect 396724 532788 396776 532840
rect 226340 532720 226392 532772
rect 396632 532720 396684 532772
rect 222200 530000 222252 530052
rect 396724 530000 396776 530052
rect 213920 529932 213972 529984
rect 396632 529932 396684 529984
rect 207020 527144 207072 527196
rect 396632 527144 396684 527196
rect 191840 509260 191892 509312
rect 396356 509260 396408 509312
rect 190460 507832 190512 507884
rect 396632 507832 396684 507884
rect 48136 498856 48188 498908
rect 177304 498856 177356 498908
rect 49424 498788 49476 498840
rect 338120 498788 338172 498840
rect 457444 498040 457496 498092
rect 462320 498040 462372 498092
rect 49332 497768 49384 497820
rect 53840 497768 53892 497820
rect 116860 497428 116912 497480
rect 133144 497428 133196 497480
rect 113548 497360 113600 497412
rect 131856 497360 131908 497412
rect 92296 497292 92348 497344
rect 131764 497292 131816 497344
rect 89536 497224 89588 497276
rect 130476 497224 130528 497276
rect 85948 497156 86000 497208
rect 130384 497156 130436 497208
rect 118608 497088 118660 497140
rect 189816 497088 189868 497140
rect 86500 497020 86552 497072
rect 189724 497020 189776 497072
rect 410524 497020 410576 497072
rect 432144 497020 432196 497072
rect 81256 496952 81308 497004
rect 185584 496952 185636 497004
rect 432604 496952 432656 497004
rect 456800 496952 456852 497004
rect 79876 496884 79928 496936
rect 188344 496884 188396 496936
rect 284944 496884 284996 496936
rect 426440 496884 426492 496936
rect 427084 496884 427136 496936
rect 430580 496884 430632 496936
rect 494704 496884 494756 496936
rect 498200 496884 498252 496936
rect 73344 496816 73396 496868
rect 75184 496816 75236 496868
rect 78312 496816 78364 496868
rect 79324 496816 79376 496868
rect 103428 496816 103480 496868
rect 150900 496816 150952 496868
rect 150992 496816 151044 496868
rect 359464 496816 359516 496868
rect 424324 496816 424376 496868
rect 426532 496816 426584 496868
rect 428464 496816 428516 496868
rect 433340 496816 433392 496868
rect 479524 496816 479576 496868
rect 495440 496816 495492 496868
rect 497464 496816 497516 496868
rect 505100 496816 505152 496868
rect 96344 496136 96396 496188
rect 184204 496136 184256 496188
rect 47952 496068 48004 496120
rect 163504 496068 163556 496120
rect 193220 496068 193272 496120
rect 415400 496068 415452 496120
rect 255320 494776 255372 494828
rect 455788 494776 455840 494828
rect 49516 494708 49568 494760
rect 340880 494708 340932 494760
rect 106096 493348 106148 493400
rect 177396 493348 177448 493400
rect 47860 493280 47912 493332
rect 175924 493280 175976 493332
rect 209780 493280 209832 493332
rect 433432 493280 433484 493332
rect 89168 491920 89220 491972
rect 166264 491920 166316 491972
rect 195980 491920 196032 491972
rect 427912 491920 427964 491972
rect 91192 490560 91244 490612
rect 170404 490560 170456 490612
rect 204904 490560 204956 490612
rect 419632 490560 419684 490612
rect 88156 489132 88208 489184
rect 162124 489132 162176 489184
rect 216680 489132 216732 489184
rect 434812 489132 434864 489184
rect 74356 487772 74408 487824
rect 155224 487772 155276 487824
rect 211804 487772 211856 487824
rect 419540 487772 419592 487824
rect 101956 486480 102008 486532
rect 176016 486480 176068 486532
rect 198740 486480 198792 486532
rect 422300 486480 422352 486532
rect 48044 486412 48096 486464
rect 409880 486412 409932 486464
rect 252560 485120 252612 485172
rect 433524 485120 433576 485172
rect 96436 485052 96488 485104
rect 383660 485052 383712 485104
rect 263600 483624 263652 483676
rect 437572 483624 437624 483676
rect 281540 482332 281592 482384
rect 443092 482332 443144 482384
rect 75184 482264 75236 482316
rect 331220 482264 331272 482316
rect 104716 480904 104768 480956
rect 182824 480904 182876 480956
rect 205640 480904 205692 480956
rect 423680 480904 423732 480956
rect 302240 479544 302292 479596
rect 449992 479544 450044 479596
rect 133788 479476 133840 479528
rect 389180 479476 389232 479528
rect 110328 478116 110380 478168
rect 181444 478116 181496 478168
rect 273260 478116 273312 478168
rect 441712 478116 441764 478168
rect 288440 476824 288492 476876
rect 445852 476824 445904 476876
rect 108856 476756 108908 476808
rect 407764 476756 407816 476808
rect 298100 475328 298152 475380
rect 448612 475328 448664 475380
rect 305000 474036 305052 474088
rect 451280 474036 451332 474088
rect 77208 473968 77260 474020
rect 342904 473968 342956 474020
rect 291200 472676 291252 472728
rect 447232 472676 447284 472728
rect 81256 472608 81308 472660
rect 356060 472608 356112 472660
rect 212540 471248 212592 471300
rect 425060 471248 425112 471300
rect 309140 469820 309192 469872
rect 452752 469820 452804 469872
rect 230480 467100 230532 467152
rect 427820 467100 427872 467152
rect 316040 465672 316092 465724
rect 454684 465672 454736 465724
rect 245660 457444 245712 457496
rect 410524 457444 410576 457496
rect 236000 454656 236052 454708
rect 429200 454656 429252 454708
rect 224960 453296 225012 453348
rect 424324 453296 424376 453348
rect 325700 451936 325752 451988
rect 458272 451936 458324 451988
rect 157248 451868 157300 451920
rect 410708 451868 410760 451920
rect 219440 450576 219492 450628
rect 284944 450576 284996 450628
rect 322940 450576 322992 450628
rect 432604 450576 432656 450628
rect 154488 450508 154540 450560
rect 409236 450508 409288 450560
rect 318800 449216 318852 449268
rect 456892 449216 456944 449268
rect 103336 449148 103388 449200
rect 410616 449148 410668 449200
rect 311900 447856 311952 447908
rect 454040 447856 454092 447908
rect 102048 447788 102100 447840
rect 411996 447788 412048 447840
rect 295340 446428 295392 446480
rect 448520 446428 448572 446480
rect 100668 446360 100720 446412
rect 410432 446360 410484 446412
rect 324320 445068 324372 445120
rect 497464 445068 497516 445120
rect 93676 445000 93728 445052
rect 378140 445000 378192 445052
rect 321560 443708 321612 443760
rect 502340 443708 502392 443760
rect 99196 443640 99248 443692
rect 411904 443640 411956 443692
rect 317420 442280 317472 442332
rect 500960 442280 501012 442332
rect 97908 442212 97960 442264
rect 411812 442212 411864 442264
rect 310888 440920 310940 440972
rect 479524 440920 479576 440972
rect 99288 440852 99340 440904
rect 357992 440852 358044 440904
rect 314660 439560 314712 439612
rect 494704 439560 494756 439612
rect 104808 439492 104860 439544
rect 410156 439492 410208 439544
rect 307852 438200 307904 438252
rect 492680 438200 492732 438252
rect 143448 438132 143500 438184
rect 394700 438132 394752 438184
rect 303896 436840 303948 436892
rect 489920 436840 489972 436892
rect 142068 436772 142120 436824
rect 409420 436772 409472 436824
rect 88248 436704 88300 436756
rect 411720 436704 411772 436756
rect 269120 435412 269172 435464
rect 465080 435412 465132 435464
rect 85488 435344 85540 435396
rect 411260 435344 411312 435396
rect 262220 434052 262272 434104
rect 460940 434052 460992 434104
rect 81164 433984 81216 434036
rect 335360 433984 335412 434036
rect 265440 432692 265492 432744
rect 457444 432692 457496 432744
rect 111708 432624 111760 432676
rect 410524 432624 410576 432676
rect 82728 432556 82780 432608
rect 411352 432556 411404 432608
rect 258448 431332 258500 431384
rect 458180 431332 458232 431384
rect 108948 431264 109000 431316
rect 410248 431264 410300 431316
rect 96528 431196 96580 431248
rect 411628 431196 411680 431248
rect 560944 430584 560996 430636
rect 580172 430584 580224 430636
rect 251456 429972 251508 430024
rect 452660 429972 452712 430024
rect 93768 429904 93820 429956
rect 411444 429904 411496 429956
rect 47768 429836 47820 429888
rect 409972 429836 410024 429888
rect 397368 428612 397420 428664
rect 445760 428612 445812 428664
rect 200856 428544 200908 428596
rect 416780 428544 416832 428596
rect 67548 428476 67600 428528
rect 410064 428476 410116 428528
rect 49608 428408 49660 428460
rect 411536 428408 411588 428460
rect 284576 427388 284628 427440
rect 444380 427388 444432 427440
rect 277584 427320 277636 427372
rect 441620 427320 441672 427372
rect 270592 427252 270644 427304
rect 440332 427252 440384 427304
rect 267096 427184 267148 427236
rect 438860 427184 438912 427236
rect 260288 427116 260340 427168
rect 436100 427116 436152 427168
rect 84016 427048 84068 427100
rect 359372 427048 359424 427100
rect 256792 426232 256844 426284
rect 434720 426232 434772 426284
rect 248512 426164 248564 426216
rect 449900 426164 449952 426216
rect 218612 426096 218664 426148
rect 420920 426096 420972 426148
rect 244464 426028 244516 426080
rect 447140 426028 447192 426080
rect 239312 425960 239364 426012
rect 445944 425960 445996 426012
rect 233976 425892 234028 425944
rect 443000 425892 443052 425944
rect 229100 425824 229152 425876
rect 440240 425824 440292 425876
rect 223580 425756 223632 425808
rect 437480 425756 437532 425808
rect 198004 425688 198056 425740
rect 418160 425688 418212 425740
rect 300676 424940 300728 424992
rect 488540 424940 488592 424992
rect 297640 424872 297692 424924
rect 485780 424872 485832 424924
rect 290648 424804 290700 424856
rect 480260 424804 480312 424856
rect 293868 424736 293920 424788
rect 483020 424736 483072 424788
rect 283656 424668 283708 424720
rect 474740 424668 474792 424720
rect 286968 424600 287020 424652
rect 477500 424600 477552 424652
rect 276664 424532 276716 424584
rect 470600 424532 470652 424584
rect 279976 424464 280028 424516
rect 473360 424464 473412 424516
rect 273168 424396 273220 424448
rect 467840 424396 467892 424448
rect 78588 424328 78640 424380
rect 185676 424328 185728 424380
rect 203248 424328 203300 424380
rect 430672 424328 430724 424380
rect 73068 423580 73120 423632
rect 218612 423580 218664 423632
rect 342904 423580 342956 423632
rect 344100 423580 344152 423632
rect 407764 423580 407816 423632
rect 408684 423580 408736 423632
rect 71688 423512 71740 423564
rect 211804 423512 211856 423564
rect 70308 423444 70360 423496
rect 204904 423444 204956 423496
rect 68928 423376 68980 423428
rect 198004 423376 198056 423428
rect 363880 423240 363932 423292
rect 410340 423240 410392 423292
rect 250536 423172 250588 423224
rect 428464 423172 428516 423224
rect 241336 423104 241388 423156
rect 427084 423104 427136 423156
rect 146208 423036 146260 423088
rect 396540 423036 396592 423088
rect 79324 422968 79376 423020
rect 330116 422968 330168 423020
rect 359464 422968 359516 423020
rect 403532 422968 403584 423020
rect 126888 422900 126940 422952
rect 382556 422900 382608 422952
rect 365628 422832 365680 422884
rect 419540 422832 419592 422884
rect 398748 422764 398800 422816
rect 412732 422764 412784 422816
rect 386236 422696 386288 422748
rect 412640 422696 412692 422748
rect 374368 422628 374420 422680
rect 416136 422628 416188 422680
rect 405648 422560 405700 422612
rect 418988 422560 419040 422612
rect 334256 422492 334308 422544
rect 351092 422492 351144 422544
rect 362224 422492 362276 422544
rect 416044 422492 416096 422544
rect 351736 422424 351788 422476
rect 360108 422424 360160 422476
rect 377864 422424 377916 422476
rect 431316 422424 431368 422476
rect 186228 422356 186280 422408
rect 347780 422356 347832 422408
rect 353208 422356 353260 422408
rect 420184 422356 420236 422408
rect 188896 422288 188948 422340
rect 368572 422288 368624 422340
rect 407672 422220 407724 422272
rect 435364 422288 435416 422340
rect 360108 421540 360160 421592
rect 552020 421540 552072 421592
rect 186964 421472 187016 421524
rect 552204 421472 552256 421524
rect 388352 421404 388404 421456
rect 418804 421404 418856 421456
rect 376208 421336 376260 421388
rect 417424 421336 417476 421388
rect 355232 421268 355284 421320
rect 413284 421268 413336 421320
rect 346308 421200 346360 421252
rect 413560 421200 413612 421252
rect 349896 421132 349948 421184
rect 429200 421132 429252 421184
rect 169760 421064 169812 421116
rect 391204 421064 391256 421116
rect 393688 421064 393740 421116
rect 438124 421064 438176 421116
rect 329104 420996 329156 421048
rect 551284 420996 551336 421048
rect 402336 420928 402388 420980
rect 414756 420928 414808 420980
rect 367376 420316 367428 420368
rect 482284 420316 482336 420368
rect 187516 420248 187568 420300
rect 413376 420248 413428 420300
rect 190368 420180 190420 420232
rect 413468 420180 413520 420232
rect 187056 420112 187108 420164
rect 414664 420112 414716 420164
rect 190736 420044 190788 420096
rect 414848 420044 414900 420096
rect 187332 419976 187384 420028
rect 421656 419976 421708 420028
rect 187148 419908 187200 419960
rect 424416 419908 424468 419960
rect 187240 419840 187292 419892
rect 428556 419840 428608 419892
rect 372528 419772 372580 419824
rect 550640 419772 550692 419824
rect 131948 419704 132000 419756
rect 425888 419704 425940 419756
rect 189356 419636 189408 419688
rect 494520 419636 494572 419688
rect 189080 419568 189132 419620
rect 552296 419568 552348 419620
rect 187424 419500 187476 419552
rect 552112 419500 552164 419552
rect 107568 419432 107620 419484
rect 186320 419432 186372 419484
rect 412088 418888 412140 418940
rect 413836 418888 413888 418940
rect 412640 418752 412692 418804
rect 506756 418752 506808 418804
rect 549904 418140 549956 418192
rect 580172 418140 580224 418192
rect 412732 417392 412784 417444
rect 531320 417392 531372 417444
rect 412088 416848 412140 416900
rect 413652 416848 413704 416900
rect 75828 416032 75880 416084
rect 178684 416032 178736 416084
rect 187424 414128 187476 414180
rect 173164 413992 173216 414044
rect 186320 413992 186372 414044
rect 187424 413924 187476 413976
rect 186964 413788 187016 413840
rect 187240 413788 187292 413840
rect 106188 413244 106240 413296
rect 180064 413244 180116 413296
rect 139308 412564 139360 412616
rect 186320 412564 186372 412616
rect 413560 411952 413612 412004
rect 470140 411952 470192 412004
rect 414848 411884 414900 411936
rect 543740 411884 543792 411936
rect 439504 411340 439556 411392
rect 445760 411340 445812 411392
rect 418896 411272 418948 411324
rect 458272 411272 458324 411324
rect 136548 411204 136600 411256
rect 186412 411204 186464 411256
rect 171048 409844 171100 409896
rect 186320 409844 186372 409896
rect 417516 409844 417568 409896
rect 519084 409844 519136 409896
rect 413652 409776 413704 409828
rect 437480 409776 437532 409828
rect 95148 409096 95200 409148
rect 188436 409096 188488 409148
rect 414756 408416 414808 408468
rect 437480 408416 437532 408468
rect 91008 407736 91060 407788
rect 188528 407736 188580 407788
rect 129648 407056 129700 407108
rect 186320 407056 186372 407108
rect 413468 407056 413520 407108
rect 437480 407056 437532 407108
rect 66168 406376 66220 406428
rect 164884 406376 164936 406428
rect 84108 404948 84160 405000
rect 189908 404948 189960 405000
rect 124128 404268 124180 404320
rect 186320 404268 186372 404320
rect 413376 404268 413428 404320
rect 437480 404268 437532 404320
rect 1308 401616 1360 401668
rect 53840 401616 53892 401668
rect 54944 401616 54996 401668
rect 104900 401616 104952 401668
rect 190000 401616 190052 401668
rect 432604 401616 432656 401668
rect 437480 401616 437532 401668
rect 121368 401548 121420 401600
rect 186320 401548 186372 401600
rect 48228 400868 48280 400920
rect 184296 400868 184348 400920
rect 413468 400188 413520 400240
rect 437480 400188 437532 400240
rect 131212 398828 131264 398880
rect 144184 398828 144236 398880
rect 425704 398828 425756 398880
rect 437480 398828 437532 398880
rect 414664 398760 414716 398812
rect 437572 398760 437624 398812
rect 131212 397468 131264 397520
rect 142804 397468 142856 397520
rect 131212 396176 131264 396228
rect 140228 396176 140280 396228
rect 131488 396108 131540 396160
rect 141516 396108 141568 396160
rect 131304 396040 131356 396092
rect 183008 396040 183060 396092
rect 162124 395972 162176 396024
rect 186320 395972 186372 396024
rect 131212 394748 131264 394800
rect 162216 394748 162268 394800
rect 131304 394680 131356 394732
rect 174544 394680 174596 394732
rect 131212 393388 131264 393440
rect 160744 393388 160796 393440
rect 132040 393320 132092 393372
rect 181536 393320 181588 393372
rect 177396 393252 177448 393304
rect 186320 393252 186372 393304
rect 413284 393252 413336 393304
rect 437480 393252 437532 393304
rect 132040 392028 132092 392080
rect 137468 392028 137520 392080
rect 131212 391960 131264 392012
rect 159364 391960 159416 392012
rect 176016 391892 176068 391944
rect 186320 391892 186372 391944
rect 413376 391212 413428 391264
rect 437572 391212 437624 391264
rect 131212 390600 131264 390652
rect 134708 390600 134760 390652
rect 131488 390532 131540 390584
rect 152556 390532 152608 390584
rect 411996 390260 412048 390312
rect 413468 390260 413520 390312
rect 131304 389784 131356 389836
rect 165068 389784 165120 389836
rect 131120 389308 131172 389360
rect 134524 389308 134576 389360
rect 131212 389240 131264 389292
rect 134616 389240 134668 389292
rect 131488 389172 131540 389224
rect 177488 389172 177540 389224
rect 435456 389172 435508 389224
rect 437756 389172 437808 389224
rect 166264 389104 166316 389156
rect 186412 389104 186464 389156
rect 170404 389036 170456 389088
rect 186320 389036 186372 389088
rect 131212 387880 131264 387932
rect 133512 387880 133564 387932
rect 131304 387812 131356 387864
rect 157984 387812 158036 387864
rect 131212 386588 131264 386640
rect 133420 386588 133472 386640
rect 131120 386384 131172 386436
rect 184480 386384 184532 386436
rect 155224 386316 155276 386368
rect 186320 386316 186372 386368
rect 417700 385636 417752 385688
rect 437480 385636 437532 385688
rect 131120 385160 131172 385212
rect 141424 385160 141476 385212
rect 131212 385092 131264 385144
rect 155316 385092 155368 385144
rect 131304 385024 131356 385076
rect 156696 385024 156748 385076
rect 131212 383732 131264 383784
rect 147036 383732 147088 383784
rect 430120 383732 430172 383784
rect 437480 383732 437532 383784
rect 131120 383664 131172 383716
rect 182916 383664 182968 383716
rect 411812 383664 411864 383716
rect 438216 383664 438268 383716
rect 131120 382304 131172 382356
rect 133328 382304 133380 382356
rect 131212 382236 131264 382288
rect 176200 382236 176252 382288
rect 435824 382236 435876 382288
rect 437940 382236 437992 382288
rect 132224 381012 132276 381064
rect 138664 381012 138716 381064
rect 131212 380944 131264 380996
rect 180156 380944 180208 380996
rect 131488 380876 131540 380928
rect 184388 380876 184440 380928
rect 411720 380876 411772 380928
rect 416780 380876 416832 380928
rect 428832 380876 428884 380928
rect 437480 380876 437532 380928
rect 144184 380808 144236 380860
rect 186412 380808 186464 380860
rect 131212 379584 131264 379636
rect 151176 379584 151228 379636
rect 131488 379516 131540 379568
rect 173348 379516 173400 379568
rect 413284 379516 413336 379568
rect 437480 379516 437532 379568
rect 142804 379448 142856 379500
rect 186320 379448 186372 379500
rect 131120 378292 131172 378344
rect 142896 378292 142948 378344
rect 131212 378224 131264 378276
rect 146944 378224 146996 378276
rect 131304 378156 131356 378208
rect 178868 378156 178920 378208
rect 554044 378156 554096 378208
rect 580172 378156 580224 378208
rect 131948 378088 132000 378140
rect 186320 378088 186372 378140
rect 131212 376796 131264 376848
rect 137376 376796 137428 376848
rect 131120 376728 131172 376780
rect 166264 376728 166316 376780
rect 422944 376728 422996 376780
rect 437480 376728 437532 376780
rect 141516 376660 141568 376712
rect 186320 376660 186372 376712
rect 131488 375436 131540 375488
rect 144184 375436 144236 375488
rect 131212 375368 131264 375420
rect 181628 375368 181680 375420
rect 421932 375368 421984 375420
rect 437480 375368 437532 375420
rect 140228 375300 140280 375352
rect 186320 375300 186372 375352
rect 183008 375232 183060 375284
rect 186412 375232 186464 375284
rect 432972 374280 433024 374332
rect 437480 374280 437532 374332
rect 131212 374144 131264 374196
rect 140136 374144 140188 374196
rect 131120 374076 131172 374128
rect 140044 374076 140096 374128
rect 131212 374008 131264 374060
rect 156604 374008 156656 374060
rect 162216 373940 162268 373992
rect 186320 373940 186372 373992
rect 131212 372648 131264 372700
rect 142804 372648 142856 372700
rect 131488 372580 131540 372632
rect 170404 372580 170456 372632
rect 174544 372512 174596 372564
rect 186320 372512 186372 372564
rect 131212 371288 131264 371340
rect 137284 371288 137336 371340
rect 426072 371288 426124 371340
rect 437480 371288 437532 371340
rect 131120 371220 131172 371272
rect 164976 371220 165028 371272
rect 411260 371220 411312 371272
rect 439688 371220 439740 371272
rect 160744 371152 160796 371204
rect 186320 371152 186372 371204
rect 181536 371084 181588 371136
rect 186412 371084 186464 371136
rect 131212 369928 131264 369980
rect 162124 369928 162176 369980
rect 131120 369860 131172 369912
rect 177396 369860 177448 369912
rect 424600 369860 424652 369912
rect 437480 369860 437532 369912
rect 159364 369792 159416 369844
rect 186320 369792 186372 369844
rect 131488 368568 131540 368620
rect 152464 368568 152516 368620
rect 131212 368500 131264 368552
rect 174544 368500 174596 368552
rect 137468 368432 137520 368484
rect 186320 368432 186372 368484
rect 131212 367208 131264 367260
rect 135904 367208 135956 367260
rect 131120 367140 131172 367192
rect 160744 367140 160796 367192
rect 131212 367072 131264 367124
rect 176016 367072 176068 367124
rect 431592 367072 431644 367124
rect 437480 367072 437532 367124
rect 134708 367004 134760 367056
rect 186412 367004 186464 367056
rect 165068 366936 165120 366988
rect 186320 366936 186372 366988
rect 131212 365712 131264 365764
rect 163688 365712 163740 365764
rect 432880 365712 432932 365764
rect 437480 365712 437532 365764
rect 152556 365644 152608 365696
rect 186320 365644 186372 365696
rect 433984 364556 434036 364608
rect 437480 364556 437532 364608
rect 131120 364420 131172 364472
rect 169116 364420 169168 364472
rect 131212 364352 131264 364404
rect 181536 364352 181588 364404
rect 558184 364352 558236 364404
rect 580172 364352 580224 364404
rect 134524 364284 134576 364336
rect 186320 364284 186372 364336
rect 131120 363060 131172 363112
rect 133236 363060 133288 363112
rect 131212 362992 131264 363044
rect 152740 362992 152792 363044
rect 131488 362924 131540 362976
rect 159364 362924 159416 362976
rect 415308 362924 415360 362976
rect 437480 362924 437532 362976
rect 177488 362856 177540 362908
rect 186320 362856 186372 362908
rect 132224 362176 132276 362228
rect 173256 362176 173308 362228
rect 131212 361632 131264 361684
rect 148508 361632 148560 361684
rect 131120 361564 131172 361616
rect 178776 361564 178828 361616
rect 134616 361496 134668 361548
rect 186320 361496 186372 361548
rect 157984 361428 158036 361480
rect 186412 361428 186464 361480
rect 131120 360272 131172 360324
rect 134524 360272 134576 360324
rect 131212 360204 131264 360256
rect 158260 360204 158312 360256
rect 414848 360204 414900 360256
rect 437480 360204 437532 360256
rect 133512 360136 133564 360188
rect 186320 360136 186372 360188
rect 411260 359320 411312 359372
rect 412916 359320 412968 359372
rect 132040 358844 132092 358896
rect 165160 358844 165212 358896
rect 131212 358776 131264 358828
rect 177580 358776 177632 358828
rect 184480 358708 184532 358760
rect 187424 358708 187476 358760
rect 131120 357484 131172 357536
rect 166448 357484 166500 357536
rect 131212 357416 131264 357468
rect 183100 357416 183152 357468
rect 414756 357416 414808 357468
rect 437480 357416 437532 357468
rect 133420 357348 133472 357400
rect 186320 357348 186372 357400
rect 156696 357280 156748 357332
rect 186412 357280 186464 357332
rect 131212 356192 131264 356244
rect 138848 356192 138900 356244
rect 131120 356124 131172 356176
rect 145748 356124 145800 356176
rect 131304 356056 131356 356108
rect 158168 356056 158220 356108
rect 428740 356056 428792 356108
rect 437480 356056 437532 356108
rect 141424 355988 141476 356040
rect 186320 355988 186372 356040
rect 131212 354764 131264 354816
rect 141516 354764 141568 354816
rect 131304 354696 131356 354748
rect 156788 354696 156840 354748
rect 427084 354696 427136 354748
rect 437480 354696 437532 354748
rect 155316 354628 155368 354680
rect 186320 354628 186372 354680
rect 131212 353336 131264 353388
rect 155500 353336 155552 353388
rect 131120 353268 131172 353320
rect 184572 353268 184624 353320
rect 424508 353268 424560 353320
rect 437480 353268 437532 353320
rect 147036 353200 147088 353252
rect 186320 353200 186372 353252
rect 182916 353132 182968 353184
rect 186412 353132 186464 353184
rect 411260 353132 411312 353184
rect 413376 353132 413428 353184
rect 131212 352044 131264 352096
rect 141700 352044 141752 352096
rect 131120 351976 131172 352028
rect 144460 351976 144512 352028
rect 131488 351908 131540 351960
rect 148416 351908 148468 351960
rect 133328 351840 133380 351892
rect 186320 351840 186372 351892
rect 131120 350616 131172 350668
rect 141608 350616 141660 350668
rect 131212 350548 131264 350600
rect 176108 350548 176160 350600
rect 420368 350548 420420 350600
rect 437480 350548 437532 350600
rect 176200 350480 176252 350532
rect 186320 350480 186372 350532
rect 131212 349188 131264 349240
rect 147220 349188 147272 349240
rect 131120 349120 131172 349172
rect 174728 349120 174780 349172
rect 435640 349120 435692 349172
rect 437480 349120 437532 349172
rect 138664 349052 138716 349104
rect 186320 349052 186372 349104
rect 184388 348984 184440 349036
rect 186412 348984 186464 349036
rect 131212 348304 131264 348356
rect 134892 348304 134944 348356
rect 131488 347828 131540 347880
rect 134800 347828 134852 347880
rect 131304 347760 131356 347812
rect 145656 347760 145708 347812
rect 423128 347760 423180 347812
rect 437480 347760 437532 347812
rect 180156 347692 180208 347744
rect 186320 347692 186372 347744
rect 131212 346468 131264 346520
rect 162308 346468 162360 346520
rect 131120 346400 131172 346452
rect 180248 346400 180300 346452
rect 430028 346400 430080 346452
rect 437480 346400 437532 346452
rect 151176 346332 151228 346384
rect 186320 346332 186372 346384
rect 131212 345176 131264 345228
rect 143080 345176 143132 345228
rect 131120 345108 131172 345160
rect 155408 345108 155460 345160
rect 131212 345040 131264 345092
rect 170588 345040 170640 345092
rect 429936 345040 429988 345092
rect 437480 345040 437532 345092
rect 173348 344972 173400 345024
rect 186320 344972 186372 345024
rect 131304 343680 131356 343732
rect 153844 343680 153896 343732
rect 411260 343680 411312 343732
rect 413008 343680 413060 343732
rect 131212 343612 131264 343664
rect 173440 343612 173492 343664
rect 142896 343544 142948 343596
rect 186320 343544 186372 343596
rect 178868 343476 178920 343528
rect 186412 343476 186464 343528
rect 131212 342320 131264 342372
rect 144368 342320 144420 342372
rect 423036 342320 423088 342372
rect 437480 342320 437532 342372
rect 131488 342252 131540 342304
rect 159548 342252 159600 342304
rect 411260 342252 411312 342304
rect 439780 342252 439832 342304
rect 146944 342184 146996 342236
rect 186320 342184 186372 342236
rect 131212 341028 131264 341080
rect 149704 341028 149756 341080
rect 131304 340960 131356 341012
rect 160928 340960 160980 341012
rect 131120 340892 131172 340944
rect 178868 340892 178920 340944
rect 166264 340824 166316 340876
rect 186320 340824 186372 340876
rect 132040 340144 132092 340196
rect 180340 340144 180392 340196
rect 131304 339532 131356 339584
rect 137560 339532 137612 339584
rect 131212 339464 131264 339516
rect 166356 339464 166408 339516
rect 435548 339464 435600 339516
rect 437848 339464 437900 339516
rect 137376 339396 137428 339448
rect 186320 339396 186372 339448
rect 181628 339328 181680 339380
rect 186412 339328 186464 339380
rect 131212 338172 131264 338224
rect 137468 338172 137520 338224
rect 131120 338104 131172 338156
rect 152648 338104 152700 338156
rect 417608 338104 417660 338156
rect 437480 338104 437532 338156
rect 144184 338036 144236 338088
rect 186320 338036 186372 338088
rect 411260 338036 411312 338088
rect 417700 338036 417752 338088
rect 131212 336880 131264 336932
rect 147036 336880 147088 336932
rect 132040 336812 132092 336864
rect 151268 336812 151320 336864
rect 131488 336744 131540 336796
rect 181628 336744 181680 336796
rect 425980 336744 426032 336796
rect 437480 336744 437532 336796
rect 140136 336676 140188 336728
rect 186320 336676 186372 336728
rect 131212 335384 131264 335436
rect 140228 335384 140280 335436
rect 131120 335316 131172 335368
rect 147128 335316 147180 335368
rect 140044 335248 140096 335300
rect 186320 335248 186372 335300
rect 156604 335180 156656 335232
rect 186412 335180 186464 335232
rect 132224 334024 132276 334076
rect 142988 334024 143040 334076
rect 131212 333956 131264 334008
rect 163596 333956 163648 334008
rect 142804 333888 142856 333940
rect 186320 333888 186372 333940
rect 131120 332732 131172 332784
rect 140136 332732 140188 332784
rect 131304 332664 131356 332716
rect 142896 332664 142948 332716
rect 131212 332596 131264 332648
rect 183008 332596 183060 332648
rect 419172 332596 419224 332648
rect 437480 332596 437532 332648
rect 170404 332528 170456 332580
rect 186320 332528 186372 332580
rect 132224 331304 132276 331356
rect 140044 331304 140096 331356
rect 131488 331236 131540 331288
rect 170496 331236 170548 331288
rect 416228 331236 416280 331288
rect 437480 331236 437532 331288
rect 137284 331168 137336 331220
rect 186412 331168 186464 331220
rect 164976 331100 165028 331152
rect 186320 331100 186372 331152
rect 417700 330488 417752 330540
rect 437572 330488 437624 330540
rect 132224 329944 132276 329996
rect 133512 329944 133564 329996
rect 131120 329876 131172 329928
rect 159456 329876 159508 329928
rect 431500 329876 431552 329928
rect 437480 329876 437532 329928
rect 131212 329808 131264 329860
rect 165068 329808 165120 329860
rect 411260 329808 411312 329860
rect 439596 329808 439648 329860
rect 131948 329740 132000 329792
rect 186320 329740 186372 329792
rect 131212 328516 131264 328568
rect 152556 328516 152608 328568
rect 131304 328448 131356 328500
rect 174636 328448 174688 328500
rect 421840 328448 421892 328500
rect 437480 328448 437532 328500
rect 177396 328380 177448 328432
rect 186320 328380 186372 328432
rect 131120 327156 131172 327208
rect 166264 327156 166316 327208
rect 131212 327088 131264 327140
rect 184480 327088 184532 327140
rect 162124 327020 162176 327072
rect 186320 327020 186372 327072
rect 174544 326952 174596 327004
rect 186412 326952 186464 327004
rect 427176 326340 427228 326392
rect 438492 326340 438544 326392
rect 132224 325796 132276 325848
rect 160836 325796 160888 325848
rect 131212 325728 131264 325780
rect 158076 325728 158128 325780
rect 131304 325660 131356 325712
rect 133420 325660 133472 325712
rect 411260 325660 411312 325712
rect 431224 325660 431276 325712
rect 152464 325592 152516 325644
rect 186320 325592 186372 325644
rect 131488 324368 131540 324420
rect 151176 324368 151228 324420
rect 131212 324300 131264 324352
rect 169024 324300 169076 324352
rect 411260 324300 411312 324352
rect 439872 324300 439924 324352
rect 551376 324300 551428 324352
rect 580172 324300 580224 324352
rect 135904 324232 135956 324284
rect 186320 324232 186372 324284
rect 131488 323076 131540 323128
rect 137376 323076 137428 323128
rect 131120 323008 131172 323060
rect 156696 323008 156748 323060
rect 131212 322940 131264 322992
rect 177488 322940 177540 322992
rect 160744 322872 160796 322924
rect 186320 322872 186372 322924
rect 176016 322804 176068 322856
rect 186412 322804 186464 322856
rect 417792 322192 417844 322244
rect 438400 322192 438452 322244
rect 131212 321648 131264 321700
rect 144276 321648 144328 321700
rect 131120 321580 131172 321632
rect 155316 321580 155368 321632
rect 173256 321512 173308 321564
rect 186320 321512 186372 321564
rect 420276 320832 420328 320884
rect 437480 320832 437532 320884
rect 131120 320220 131172 320272
rect 162216 320220 162268 320272
rect 131212 320152 131264 320204
rect 176016 320152 176068 320204
rect 163688 320084 163740 320136
rect 186320 320084 186372 320136
rect 132224 318860 132276 318912
rect 156604 318860 156656 318912
rect 131212 318792 131264 318844
rect 173256 318792 173308 318844
rect 429844 318792 429896 318844
rect 437480 318792 437532 318844
rect 169116 318724 169168 318776
rect 186320 318724 186372 318776
rect 131488 317432 131540 317484
rect 174544 317432 174596 317484
rect 411260 317432 411312 317484
rect 425796 317432 425848 317484
rect 159364 317364 159416 317416
rect 186320 317364 186372 317416
rect 431960 317364 432012 317416
rect 438308 317364 438360 317416
rect 181536 317296 181588 317348
rect 186412 317296 186464 317348
rect 132224 316072 132276 316124
rect 133328 316072 133380 316124
rect 131212 316004 131264 316056
rect 155224 316004 155276 316056
rect 411260 316004 411312 316056
rect 428464 316004 428516 316056
rect 133236 315936 133288 315988
rect 186320 315936 186372 315988
rect 131488 314712 131540 314764
rect 138756 314712 138808 314764
rect 131212 314644 131264 314696
rect 180156 314644 180208 314696
rect 419080 314644 419132 314696
rect 437480 314644 437532 314696
rect 152740 314576 152792 314628
rect 186320 314576 186372 314628
rect 131304 313896 131356 313948
rect 170404 313896 170456 313948
rect 131212 313352 131264 313404
rect 152464 313352 152516 313404
rect 131120 313284 131172 313336
rect 157984 313284 158036 313336
rect 411260 313284 411312 313336
rect 421564 313284 421616 313336
rect 421748 313284 421800 313336
rect 437480 313284 437532 313336
rect 148508 313216 148560 313268
rect 186412 313216 186464 313268
rect 178776 313148 178828 313200
rect 186320 313148 186372 313200
rect 131120 311924 131172 311976
rect 148324 311924 148376 311976
rect 131212 311856 131264 311908
rect 164976 311856 165028 311908
rect 411260 311856 411312 311908
rect 424324 311856 424376 311908
rect 434076 311856 434128 311908
rect 438768 311856 438820 311908
rect 556804 311856 556856 311908
rect 580172 311856 580224 311908
rect 134524 311788 134576 311840
rect 186320 311788 186372 311840
rect 131488 310564 131540 310616
rect 159364 310564 159416 310616
rect 131212 310496 131264 310548
rect 182916 310496 182968 310548
rect 414664 310496 414716 310548
rect 437480 310496 437532 310548
rect 180340 310428 180392 310480
rect 186320 310428 186372 310480
rect 131304 309748 131356 309800
rect 184388 309748 184440 309800
rect 420920 309748 420972 309800
rect 431960 309748 432012 309800
rect 131120 309612 131172 309664
rect 134708 309612 134760 309664
rect 131212 309136 131264 309188
rect 141424 309136 141476 309188
rect 411260 309136 411312 309188
rect 420920 309136 420972 309188
rect 158260 309068 158312 309120
rect 186320 309068 186372 309120
rect 410524 309068 410576 309120
rect 417792 309068 417844 309120
rect 165160 309000 165212 309052
rect 186412 309000 186464 309052
rect 131212 307912 131264 307964
rect 134616 307912 134668 307964
rect 131120 307844 131172 307896
rect 145564 307844 145616 307896
rect 131488 307776 131540 307828
rect 160744 307776 160796 307828
rect 432696 307776 432748 307828
rect 437480 307776 437532 307828
rect 177580 307708 177632 307760
rect 186320 307708 186372 307760
rect 424692 307028 424744 307080
rect 438400 307028 438452 307080
rect 131120 306416 131172 306468
rect 142804 306416 142856 306468
rect 131212 306348 131264 306400
rect 177396 306348 177448 306400
rect 166448 306280 166500 306332
rect 186320 306280 186372 306332
rect 409972 306280 410024 306332
rect 430120 306280 430172 306332
rect 131488 305124 131540 305176
rect 178776 305124 178828 305176
rect 131120 305056 131172 305108
rect 137284 305056 137336 305108
rect 131212 304988 131264 305040
rect 133236 304988 133288 305040
rect 428648 304988 428700 305040
rect 437480 304988 437532 305040
rect 158168 304920 158220 304972
rect 186412 304920 186464 304972
rect 183100 304852 183152 304904
rect 186688 304852 186740 304904
rect 421012 304240 421064 304292
rect 435824 304240 435876 304292
rect 131304 303696 131356 303748
rect 144184 303696 144236 303748
rect 131212 303628 131264 303680
rect 181536 303628 181588 303680
rect 411260 303628 411312 303680
rect 421012 303628 421064 303680
rect 435732 303628 435784 303680
rect 438676 303628 438728 303680
rect 145748 303560 145800 303612
rect 186320 303560 186372 303612
rect 131120 302268 131172 302320
rect 135904 302268 135956 302320
rect 131212 302200 131264 302252
rect 162124 302200 162176 302252
rect 432788 302200 432840 302252
rect 438032 302200 438084 302252
rect 138848 302132 138900 302184
rect 186320 302132 186372 302184
rect 411536 302132 411588 302184
rect 428832 302132 428884 302184
rect 431408 301452 431460 301504
rect 437572 301452 437624 301504
rect 131212 300908 131264 300960
rect 138664 300908 138716 300960
rect 131488 300840 131540 300892
rect 146944 300840 146996 300892
rect 156788 300772 156840 300824
rect 186320 300772 186372 300824
rect 410524 300772 410576 300824
rect 413284 300772 413336 300824
rect 439780 300772 439832 300824
rect 552204 300772 552256 300824
rect 439872 300704 439924 300756
rect 550548 300704 550600 300756
rect 428832 300092 428884 300144
rect 438584 300092 438636 300144
rect 131120 299888 131172 299940
rect 134524 299888 134576 299940
rect 141516 299412 141568 299464
rect 186320 299412 186372 299464
rect 184572 299344 184624 299396
rect 186412 299344 186464 299396
rect 522304 298120 522356 298172
rect 580172 298120 580224 298172
rect 155500 298052 155552 298104
rect 186320 298052 186372 298104
rect 418988 298052 419040 298104
rect 545488 298052 545540 298104
rect 421656 297984 421708 298036
rect 528744 297984 528796 298036
rect 411260 297916 411312 297968
rect 422944 297916 422996 297968
rect 431316 297916 431368 297968
rect 520280 297916 520332 297968
rect 428556 297848 428608 297900
rect 512000 297848 512052 297900
rect 424416 297780 424468 297832
rect 503168 297780 503220 297832
rect 425888 297712 425940 297764
rect 494704 297712 494756 297764
rect 132132 297372 132184 297424
rect 141516 297372 141568 297424
rect 141700 296624 141752 296676
rect 186320 296624 186372 296676
rect 410156 296624 410208 296676
rect 421932 296624 421984 296676
rect 422944 295944 422996 295996
rect 438400 295944 438452 295996
rect 477500 295944 477552 295996
rect 544384 295944 544436 295996
rect 144460 295264 144512 295316
rect 186320 295264 186372 295316
rect 148416 295196 148468 295248
rect 186412 295196 186464 295248
rect 420184 294652 420236 294704
rect 512000 294652 512052 294704
rect 416136 294584 416188 294636
rect 512184 294584 512236 294636
rect 141608 293904 141660 293956
rect 186320 293904 186372 293956
rect 439688 293904 439740 293956
rect 441620 293904 441672 293956
rect 419632 293224 419684 293276
rect 432972 293224 433024 293276
rect 411260 292544 411312 292596
rect 419632 292544 419684 292596
rect 176108 292476 176160 292528
rect 186320 292476 186372 292528
rect 419632 291864 419684 291916
rect 437020 291864 437072 291916
rect 131948 291796 132000 291848
rect 176200 291796 176252 291848
rect 416044 291796 416096 291848
rect 512092 291796 512144 291848
rect 411260 291184 411312 291236
rect 419632 291184 419684 291236
rect 147220 291116 147272 291168
rect 186412 291116 186464 291168
rect 174728 291048 174780 291100
rect 186320 291048 186372 291100
rect 134892 289756 134944 289808
rect 186320 289756 186372 289808
rect 415400 289076 415452 289128
rect 426072 289076 426124 289128
rect 411260 288396 411312 288448
rect 415400 288396 415452 288448
rect 145656 288328 145708 288380
rect 186320 288328 186372 288380
rect 411260 287036 411312 287088
rect 418160 287036 418212 287088
rect 424600 287036 424652 287088
rect 134800 286968 134852 287020
rect 186320 286968 186372 287020
rect 180248 286900 180300 286952
rect 186412 286900 186464 286952
rect 162308 285608 162360 285660
rect 186320 285608 186372 285660
rect 419816 284928 419868 284980
rect 431592 284928 431644 284980
rect 411260 284316 411312 284368
rect 419816 284316 419868 284368
rect 143080 284248 143132 284300
rect 186320 284248 186372 284300
rect 418252 283636 418304 283688
rect 432880 283636 432932 283688
rect 414940 283568 414992 283620
rect 438492 283568 438544 283620
rect 411260 282888 411312 282940
rect 418252 282888 418304 282940
rect 155408 282820 155460 282872
rect 186320 282820 186372 282872
rect 170588 282752 170640 282804
rect 186412 282752 186464 282804
rect 153844 281460 153896 281512
rect 186320 281460 186372 281512
rect 418344 280780 418396 280832
rect 433984 280780 434036 280832
rect 411260 280168 411312 280220
rect 418344 280168 418396 280220
rect 173440 280100 173492 280152
rect 186320 280100 186372 280152
rect 132040 279420 132092 279472
rect 173348 279420 173400 279472
rect 411260 279420 411312 279472
rect 415308 279420 415360 279472
rect 416872 279420 416924 279472
rect 144368 278672 144420 278724
rect 186320 278672 186372 278724
rect 159548 277312 159600 277364
rect 186320 277312 186372 277364
rect 178868 277244 178920 277296
rect 186412 277244 186464 277296
rect 411260 276836 411312 276888
rect 414020 276836 414072 276888
rect 414848 276836 414900 276888
rect 160928 275952 160980 276004
rect 186320 275952 186372 276004
rect 416688 275272 416740 275324
rect 436928 275272 436980 275324
rect 411260 274660 411312 274712
rect 415492 274660 415544 274712
rect 416688 274660 416740 274712
rect 149704 274592 149756 274644
rect 186320 274592 186372 274644
rect 137560 273164 137612 273216
rect 186320 273164 186372 273216
rect 411260 273164 411312 273216
rect 413100 273164 413152 273216
rect 414756 273164 414808 273216
rect 166356 273096 166408 273148
rect 186412 273096 186464 273148
rect 515404 271872 515456 271924
rect 579804 271872 579856 271924
rect 152648 271804 152700 271856
rect 186320 271804 186372 271856
rect 416688 271124 416740 271176
rect 428740 271124 428792 271176
rect 411260 270512 411312 270564
rect 415584 270512 415636 270564
rect 416688 270512 416740 270564
rect 137468 270444 137520 270496
rect 186320 270444 186372 270496
rect 151268 269016 151320 269068
rect 186320 269016 186372 269068
rect 181628 268948 181680 269000
rect 186412 268948 186464 269000
rect 416964 268336 417016 268388
rect 427084 268336 427136 268388
rect 411260 267724 411312 267776
rect 416964 267724 417016 267776
rect 147036 267656 147088 267708
rect 186320 267656 186372 267708
rect 411260 266976 411312 267028
rect 414112 266976 414164 267028
rect 424508 266976 424560 267028
rect 147128 266296 147180 266348
rect 186320 266296 186372 266348
rect 140228 264868 140280 264920
rect 186320 264868 186372 264920
rect 163596 264800 163648 264852
rect 186412 264800 186464 264852
rect 411260 263576 411312 263628
rect 415676 263576 415728 263628
rect 420368 263576 420420 263628
rect 142988 263508 143040 263560
rect 186320 263508 186372 263560
rect 411260 262828 411312 262880
rect 414204 262828 414256 262880
rect 435640 262828 435692 262880
rect 140136 262148 140188 262200
rect 186320 262148 186372 262200
rect 142896 260788 142948 260840
rect 186320 260788 186372 260840
rect 411260 259428 411312 259480
rect 417056 259428 417108 259480
rect 423128 259428 423180 259480
rect 140044 259360 140096 259412
rect 186320 259360 186372 259412
rect 183008 259292 183060 259344
rect 186412 259292 186464 259344
rect 411260 258680 411312 258732
rect 414296 258680 414348 258732
rect 430028 258680 430080 258732
rect 555424 258068 555476 258120
rect 580172 258068 580224 258120
rect 170496 258000 170548 258052
rect 186320 258000 186372 258052
rect 159456 256640 159508 256692
rect 186320 256640 186372 256692
rect 417332 255960 417384 256012
rect 429936 255960 429988 256012
rect 430028 255960 430080 256012
rect 438308 255960 438360 256012
rect 411260 255280 411312 255332
rect 417148 255280 417200 255332
rect 417332 255280 417384 255332
rect 133512 255212 133564 255264
rect 186320 255212 186372 255264
rect 165068 255144 165120 255196
rect 186412 255144 186464 255196
rect 411260 254532 411312 254584
rect 414388 254532 414440 254584
rect 423036 254532 423088 254584
rect 152556 253852 152608 253904
rect 186320 253852 186372 253904
rect 174636 252492 174688 252544
rect 186320 252492 186372 252544
rect 410800 252492 410852 252544
rect 427176 252492 427228 252544
rect 166264 251132 166316 251184
rect 186320 251132 186372 251184
rect 184480 251064 184532 251116
rect 186412 251064 186464 251116
rect 411260 250452 411312 250504
rect 411628 250452 411680 250504
rect 435548 250452 435600 250504
rect 160836 249704 160888 249756
rect 186320 249704 186372 249756
rect 133420 248344 133472 248396
rect 186320 248344 186372 248396
rect 411812 247664 411864 247716
rect 417608 247664 417660 247716
rect 158076 246984 158128 247036
rect 186320 246984 186372 247036
rect 169024 246916 169076 246968
rect 186412 246916 186464 246968
rect 417332 246304 417384 246356
rect 425980 246304 426032 246356
rect 411260 245624 411312 245676
rect 417332 245624 417384 245676
rect 151176 245556 151228 245608
rect 186320 245556 186372 245608
rect 520924 244264 520976 244316
rect 579804 244264 579856 244316
rect 156696 244196 156748 244248
rect 186320 244196 186372 244248
rect 410800 244196 410852 244248
rect 417700 244196 417752 244248
rect 137376 242836 137428 242888
rect 186320 242836 186372 242888
rect 411260 241816 411312 241868
rect 414480 241816 414532 241868
rect 419172 241816 419224 241868
rect 155316 241408 155368 241460
rect 186412 241408 186464 241460
rect 177488 241340 177540 241392
rect 186320 241340 186372 241392
rect 144276 240048 144328 240100
rect 186320 240048 186372 240100
rect 411260 240048 411312 240100
rect 416228 240048 416280 240100
rect 162216 238688 162268 238740
rect 186320 238688 186372 238740
rect 416688 238008 416740 238060
rect 431500 238008 431552 238060
rect 411260 237396 411312 237448
rect 415768 237396 415820 237448
rect 416688 237396 416740 237448
rect 176016 237328 176068 237380
rect 186320 237328 186372 237380
rect 409420 237328 409472 237380
rect 421840 237328 421892 237380
rect 176200 237260 176252 237312
rect 186412 237260 186464 237312
rect 156604 235900 156656 235952
rect 186320 235900 186372 235952
rect 173256 234540 173308 234592
rect 186320 234540 186372 234592
rect 411260 233248 411312 233300
rect 415860 233248 415912 233300
rect 420276 233248 420328 233300
rect 141516 233180 141568 233232
rect 186320 233180 186372 233232
rect 469220 233180 469272 233232
rect 579988 233180 580040 233232
rect 174544 233112 174596 233164
rect 186412 233112 186464 233164
rect 133328 231752 133380 231804
rect 186320 231752 186372 231804
rect 411352 231072 411404 231124
rect 412088 231072 412140 231124
rect 434076 231072 434128 231124
rect 155224 230392 155276 230444
rect 186320 230392 186372 230444
rect 415952 229712 416004 229764
rect 428832 229712 428884 229764
rect 411260 229100 411312 229152
rect 415952 229100 416004 229152
rect 138756 229032 138808 229084
rect 186320 229032 186372 229084
rect 180156 228964 180208 229016
rect 186412 228964 186464 229016
rect 409512 227740 409564 227792
rect 414940 227740 414992 227792
rect 170404 227672 170456 227724
rect 186320 227672 186372 227724
rect 157984 226244 158036 226296
rect 186320 226244 186372 226296
rect 411536 225564 411588 225616
rect 424692 225564 424744 225616
rect 152464 224884 152516 224936
rect 186320 224884 186372 224936
rect 184388 224816 184440 224868
rect 186412 224816 186464 224868
rect 415308 224204 415360 224256
rect 429844 224204 429896 224256
rect 411260 223592 411312 223644
rect 414572 223592 414624 223644
rect 415308 223592 415360 223644
rect 148324 223524 148376 223576
rect 186320 223524 186372 223576
rect 164976 222096 165028 222148
rect 186320 222096 186372 222148
rect 410800 222096 410852 222148
rect 435732 222096 435784 222148
rect 159364 220736 159416 220788
rect 186412 220736 186464 220788
rect 182916 220668 182968 220720
rect 186504 220668 186556 220720
rect 411996 220056 412048 220108
rect 419080 220056 419132 220108
rect 134708 219376 134760 219428
rect 186320 219376 186372 219428
rect 460940 219376 460992 219428
rect 580172 219376 580224 219428
rect 141424 217948 141476 218000
rect 186320 217948 186372 218000
rect 411260 217268 411312 217320
rect 414756 217268 414808 217320
rect 421748 217268 421800 217320
rect 145564 216588 145616 216640
rect 186320 216588 186372 216640
rect 412088 216588 412140 216640
rect 432788 216588 432840 216640
rect 134616 215228 134668 215280
rect 186412 215228 186464 215280
rect 160744 215160 160796 215212
rect 186320 215160 186372 215212
rect 142804 213868 142856 213920
rect 186320 213868 186372 213920
rect 411260 213324 411312 213376
rect 414664 213324 414716 213376
rect 177396 212440 177448 212492
rect 186320 212440 186372 212492
rect 411260 211760 411312 211812
rect 413192 211760 413244 211812
rect 432696 211760 432748 211812
rect 137284 211080 137336 211132
rect 186320 211080 186372 211132
rect 178776 211012 178828 211064
rect 186412 211012 186464 211064
rect 133236 209720 133288 209772
rect 186320 209720 186372 209772
rect 411628 209040 411680 209092
rect 431408 209040 431460 209092
rect 144184 208292 144236 208344
rect 186320 208292 186372 208344
rect 411352 207612 411404 207664
rect 428648 207612 428700 207664
rect 135904 206932 135956 206984
rect 186320 206932 186372 206984
rect 181536 206864 181588 206916
rect 186412 206864 186464 206916
rect 519544 205640 519596 205692
rect 580172 205640 580224 205692
rect 162124 205572 162176 205624
rect 186320 205572 186372 205624
rect 413928 204892 413980 204944
rect 436836 204892 436888 204944
rect 411260 204280 411312 204332
rect 413376 204280 413428 204332
rect 413928 204280 413980 204332
rect 146944 204212 146996 204264
rect 186320 204212 186372 204264
rect 415308 203532 415360 203584
rect 430028 203532 430080 203584
rect 411260 203056 411312 203108
rect 414848 203056 414900 203108
rect 415308 203056 415360 203108
rect 138664 202784 138716 202836
rect 186412 202784 186464 202836
rect 173348 202716 173400 202768
rect 186320 202716 186372 202768
rect 412640 202104 412692 202156
rect 536840 202104 536892 202156
rect 134524 201424 134576 201476
rect 186320 201424 186372 201476
rect 411260 200744 411312 200796
rect 422944 200744 422996 200796
rect 401048 199996 401100 200048
rect 412272 199996 412324 200048
rect 405004 199928 405056 199980
rect 415400 199928 415452 199980
rect 400956 199860 401008 199912
rect 411444 199860 411496 199912
rect 399576 199792 399628 199844
rect 412180 199792 412232 199844
rect 407764 199724 407816 199776
rect 419816 199724 419868 199776
rect 398380 199656 398432 199708
rect 410432 199656 410484 199708
rect 194600 199588 194652 199640
rect 195612 199588 195664 199640
rect 399208 199588 399260 199640
rect 411812 199588 411864 199640
rect 406384 199520 406436 199572
rect 419724 199520 419776 199572
rect 393228 199452 393280 199504
rect 411260 199452 411312 199504
rect 261852 199384 261904 199436
rect 552020 199384 552072 199436
rect 189724 199112 189776 199164
rect 239588 199112 239640 199164
rect 188344 199044 188396 199096
rect 259644 199044 259696 199096
rect 189816 198976 189868 199028
rect 327540 198976 327592 199028
rect 185584 198908 185636 198960
rect 271972 198908 272024 198960
rect 296168 198908 296220 198960
rect 436744 198908 436796 198960
rect 131856 198840 131908 198892
rect 311992 198840 312044 198892
rect 133144 198772 133196 198824
rect 319628 198772 319680 198824
rect 344192 198772 344244 198824
rect 425704 198772 425756 198824
rect 190000 198704 190052 198756
rect 194600 198704 194652 198756
rect 208216 198704 208268 198756
rect 435456 198704 435508 198756
rect 182824 198636 182876 198688
rect 379612 198636 379664 198688
rect 397368 198636 397420 198688
rect 413376 198636 413428 198688
rect 184204 198568 184256 198620
rect 351460 198568 351512 198620
rect 368112 198568 368164 198620
rect 432604 198568 432656 198620
rect 188436 198500 188488 198552
rect 339500 198500 339552 198552
rect 364248 198500 364300 198552
rect 412640 198500 412692 198552
rect 188528 198432 188580 198484
rect 323492 198432 323544 198484
rect 397276 198432 397328 198484
rect 413192 198432 413244 198484
rect 163504 198364 163556 198416
rect 267740 198364 267792 198416
rect 397184 198364 397236 198416
rect 414756 198364 414808 198416
rect 184296 198296 184348 198348
rect 279516 198296 279568 198348
rect 395804 198296 395856 198348
rect 414112 198296 414164 198348
rect 177304 198228 177356 198280
rect 255596 198228 255648 198280
rect 395896 198228 395948 198280
rect 414388 198228 414440 198280
rect 175924 198160 175976 198212
rect 243636 198160 243688 198212
rect 395712 198160 395764 198212
rect 414296 198160 414348 198212
rect 185676 198092 185728 198144
rect 247500 198092 247552 198144
rect 395436 198092 395488 198144
rect 178684 198024 178736 198076
rect 235540 198024 235592 198076
rect 323584 198024 323636 198076
rect 395620 198024 395672 198076
rect 396724 198092 396776 198144
rect 415492 198092 415544 198144
rect 414204 198024 414256 198076
rect 164884 197956 164936 198008
rect 219532 197956 219584 198008
rect 224224 197956 224276 198008
rect 261852 197956 261904 198008
rect 264152 197956 264204 198008
rect 280252 197956 280304 198008
rect 319444 197956 319496 198008
rect 391572 197956 391624 198008
rect 395528 197956 395580 198008
rect 415584 197956 415636 198008
rect 189908 197888 189960 197940
rect 227720 197888 227772 197940
rect 403624 197888 403676 197940
rect 418344 197888 418396 197940
rect 188896 197820 188948 197872
rect 212540 197820 212592 197872
rect 399760 197820 399812 197872
rect 411352 197820 411404 197872
rect 186228 197752 186280 197804
rect 200120 197752 200172 197804
rect 400864 197752 400916 197804
rect 411720 197752 411772 197804
rect 395620 197344 395672 197396
rect 395804 197344 395856 197396
rect 148968 197276 149020 197328
rect 383660 197276 383712 197328
rect 151084 197208 151136 197260
rect 375564 197208 375616 197260
rect 131028 197140 131080 197192
rect 355508 197140 355560 197192
rect 131764 197072 131816 197124
rect 331588 197072 331640 197124
rect 130476 197004 130528 197056
rect 315580 197004 315632 197056
rect 130384 196936 130436 196988
rect 303620 196936 303672 196988
rect 397828 196800 397880 196852
rect 409328 196800 409380 196852
rect 398748 196732 398800 196784
rect 410340 196732 410392 196784
rect 399116 196664 399168 196716
rect 411904 196664 411956 196716
rect 399024 196596 399076 196648
rect 411996 196596 412048 196648
rect 397000 195916 397052 195968
rect 415952 195916 416004 195968
rect 395988 195848 396040 195900
rect 415860 195848 415912 195900
rect 394424 195780 394476 195832
rect 414480 195780 414532 195832
rect 396908 195712 396960 195764
rect 417148 195712 417200 195764
rect 392676 195644 392728 195696
rect 413100 195644 413152 195696
rect 392584 195576 392636 195628
rect 414020 195576 414072 195628
rect 393136 195508 393188 195560
rect 415768 195508 415820 195560
rect 394332 195440 394384 195492
rect 417056 195440 417108 195492
rect 392952 195372 393004 195424
rect 415676 195372 415728 195424
rect 393044 195304 393096 195356
rect 417240 195304 417292 195356
rect 400128 195236 400180 195288
rect 503720 195236 503772 195288
rect 397092 195168 397144 195220
rect 414572 195168 414624 195220
rect 403808 195100 403860 195152
rect 421012 195100 421064 195152
rect 403716 195032 403768 195084
rect 418252 195032 418304 195084
rect 204168 193808 204220 193860
rect 284944 193808 284996 193860
rect 452660 193128 452712 193180
rect 580172 193128 580224 193180
rect 401232 192924 401284 192976
rect 419632 192924 419684 192976
rect 394608 192856 394660 192908
rect 414848 192856 414900 192908
rect 401140 192788 401192 192840
rect 420920 192788 420972 192840
rect 394516 192720 394568 192772
rect 414664 192720 414716 192772
rect 392768 192652 392820 192704
rect 416872 192652 416924 192704
rect 393964 192584 394016 192636
rect 418160 192584 418212 192636
rect 389824 192516 389876 192568
rect 416780 192516 416832 192568
rect 189264 192448 189316 192500
rect 224960 192448 225012 192500
rect 282184 192448 282236 192500
rect 413008 192448 413060 192500
rect 400680 191836 400732 191888
rect 404268 191836 404320 191888
rect 188712 191156 188764 191208
rect 236000 191156 236052 191208
rect 187148 191088 187200 191140
rect 509240 191088 509292 191140
rect 189172 189728 189224 189780
rect 248420 189728 248472 189780
rect 282368 189728 282420 189780
rect 412916 189728 412968 189780
rect 169852 188300 169904 188352
rect 407120 188300 407172 188352
rect 397460 187688 397512 187740
rect 400680 187688 400732 187740
rect 187240 186940 187292 186992
rect 286324 186940 286376 186992
rect 187516 184152 187568 184204
rect 395344 184152 395396 184204
rect 390560 182860 390612 182912
rect 397460 182860 397512 182912
rect 188804 182792 188856 182844
rect 466460 182792 466512 182844
rect 387340 181024 387392 181076
rect 390560 181024 390612 181076
rect 186872 180072 186924 180124
rect 309784 180072 309836 180124
rect 443000 179324 443052 179376
rect 580172 179324 580224 179376
rect 274640 178644 274692 178696
rect 349804 178644 349856 178696
rect 187608 177284 187660 177336
rect 305644 177284 305696 177336
rect 384304 175176 384356 175228
rect 387340 175176 387392 175228
rect 382280 168376 382332 168428
rect 384304 168376 384356 168428
rect 289084 165588 289136 165640
rect 580172 165588 580224 165640
rect 381544 164772 381596 164824
rect 382280 164772 382332 164824
rect 187332 155184 187384 155236
rect 510896 155184 510948 155236
rect 379520 154300 379572 154352
rect 381544 154300 381596 154352
rect 428464 153824 428516 153876
rect 580632 153824 580684 153876
rect 431224 153144 431276 153196
rect 580172 153144 580224 153196
rect 170220 152464 170272 152516
rect 371240 152464 371292 152516
rect 168932 151036 168984 151088
rect 282920 151036 282972 151088
rect 424324 151036 424376 151088
rect 580540 151036 580592 151088
rect 188988 149676 189040 149728
rect 281540 149676 281592 149728
rect 282276 149676 282328 149728
rect 412824 149676 412876 149728
rect 421564 149676 421616 149728
rect 580356 149676 580408 149728
rect 168840 148316 168892 148368
rect 299480 148316 299532 148368
rect 425796 148316 425848 148368
rect 580264 148316 580316 148368
rect 406016 146956 406068 147008
rect 439504 146956 439556 147008
rect 439596 146956 439648 147008
rect 512276 146956 512328 147008
rect 211160 146888 211212 146940
rect 280160 146888 280212 146940
rect 282460 146888 282512 146940
rect 412732 146888 412784 146940
rect 485780 146888 485832 146940
rect 562324 146888 562376 146940
rect 377312 146208 377364 146260
rect 379520 146276 379572 146328
rect 169208 145528 169260 145580
rect 215300 145528 215352 145580
rect 398472 144236 398524 144288
rect 410524 144236 410576 144288
rect 189080 144168 189132 144220
rect 580448 144168 580500 144220
rect 194600 143488 194652 143540
rect 195060 143488 195112 143540
rect 418896 143488 418948 143540
rect 192576 143420 192628 143472
rect 406016 143420 406068 143472
rect 188344 142876 188396 142928
rect 195060 142876 195112 142928
rect 398564 142876 398616 142928
rect 409420 142876 409472 142928
rect 417424 142876 417476 142928
rect 454684 142876 454736 142928
rect 176200 142808 176252 142860
rect 191840 142808 191892 142860
rect 192576 142808 192628 142860
rect 274272 142808 274324 142860
rect 323584 142808 323636 142860
rect 376024 142808 376076 142860
rect 377312 142808 377364 142860
rect 399392 142808 399444 142860
rect 411536 142808 411588 142860
rect 418804 142808 418856 142860
rect 479156 142808 479208 142860
rect 20 142672 72 142724
rect 1308 142672 1360 142724
rect 1308 142196 1360 142248
rect 176200 142196 176252 142248
rect 1400 142128 1452 142180
rect 188344 142128 188396 142180
rect 398656 141720 398708 141772
rect 409512 141720 409564 141772
rect 394148 141652 394200 141704
rect 405004 141652 405056 141704
rect 399300 141584 399352 141636
rect 411628 141584 411680 141636
rect 438216 141584 438268 141636
rect 509332 141584 509384 141636
rect 394240 141516 394292 141568
rect 406384 141516 406436 141568
rect 438124 141516 438176 141568
rect 509424 141516 509476 141568
rect 395804 141448 395856 141500
rect 419540 141448 419592 141500
rect 435364 141448 435416 141500
rect 510712 141448 510764 141500
rect 198740 141380 198792 141432
rect 518164 141380 518216 141432
rect 168196 141040 168248 141092
rect 173164 141040 173216 141092
rect 170128 140972 170180 141024
rect 393780 140972 393832 141024
rect 394240 140972 394292 141024
rect 169668 140904 169720 140956
rect 393872 140904 393924 140956
rect 169576 140836 169628 140888
rect 394148 140836 394200 140888
rect 170036 140768 170088 140820
rect 400220 140768 400272 140820
rect 401232 140768 401284 140820
rect 397920 140700 397972 140752
rect 410156 140700 410208 140752
rect 169944 140292 169996 140344
rect 394240 140564 394292 140616
rect 403624 140564 403676 140616
rect 398196 140292 398248 140344
rect 410064 140292 410116 140344
rect 167552 140224 167604 140276
rect 392676 140224 392728 140276
rect 398012 140224 398064 140276
rect 409880 140224 409932 140276
rect 168380 140156 168432 140208
rect 394148 140156 394200 140208
rect 407764 140156 407816 140208
rect 167460 140088 167512 140140
rect 395436 140088 395488 140140
rect 398104 140088 398156 140140
rect 409972 140088 410024 140140
rect 167828 140020 167880 140072
rect 395528 140020 395580 140072
rect 396080 140020 396132 140072
rect 396724 140020 396776 140072
rect 398288 140020 398340 140072
rect 410248 140020 410300 140072
rect 169300 139952 169352 140004
rect 396540 139952 396592 140004
rect 403808 139952 403860 140004
rect 168012 139884 168064 139936
rect 395160 139884 395212 139936
rect 395620 139884 395672 139936
rect 396816 139884 396868 139936
rect 403716 139884 403768 139936
rect 167920 139816 167972 139868
rect 396080 139816 396132 139868
rect 169392 139748 169444 139800
rect 398196 139748 398248 139800
rect 398840 139748 398892 139800
rect 400128 139748 400180 139800
rect 169116 139680 169168 139732
rect 398012 139680 398064 139732
rect 168288 139612 168340 139664
rect 398104 139612 398156 139664
rect 166908 139544 166960 139596
rect 396632 139544 396684 139596
rect 401140 139544 401192 139596
rect 165528 139476 165580 139528
rect 396816 139476 396868 139528
rect 167644 139408 167696 139460
rect 398840 139408 398892 139460
rect 400588 137844 400640 137896
rect 401048 137844 401100 137896
rect 167552 136076 167604 136128
rect 168012 136076 168064 136128
rect 167552 135940 167604 135992
rect 168380 135940 168432 135992
rect 305644 135192 305696 135244
rect 397460 135192 397512 135244
rect 167828 134172 167880 134224
rect 168196 134172 168248 134224
rect 167552 134036 167604 134088
rect 167828 134036 167880 134088
rect 309784 133832 309836 133884
rect 397460 133832 397512 133884
rect 347780 129684 347832 129736
rect 397460 129684 397512 129736
rect 393872 128324 393924 128376
rect 398380 128324 398432 128376
rect 562324 126896 562376 126948
rect 579712 126896 579764 126948
rect 375012 126624 375064 126676
rect 376024 126624 376076 126676
rect 287060 125536 287112 125588
rect 397460 125536 397512 125588
rect 372620 124176 372672 124228
rect 375012 124176 375064 124228
rect 349804 124108 349856 124160
rect 397460 124108 397512 124160
rect 392768 123428 392820 123480
rect 397920 123428 397972 123480
rect 371884 123088 371936 123140
rect 372620 123088 372672 123140
rect 400588 121388 400640 121440
rect 400956 121388 401008 121440
rect 286324 120028 286376 120080
rect 397460 120028 397512 120080
rect 395620 118668 395672 118720
rect 396080 118668 396132 118720
rect 396632 118600 396684 118652
rect 398104 118600 398156 118652
rect 551284 113092 551336 113144
rect 579712 113092 579764 113144
rect 396540 113024 396592 113076
rect 397552 113024 397604 113076
rect 395160 106224 395212 106276
rect 399576 106224 399628 106276
rect 393780 104796 393832 104848
rect 397460 104796 397512 104848
rect 394056 102076 394108 102128
rect 397460 102076 397512 102128
rect 394148 99288 394200 99340
rect 397460 99288 397512 99340
rect 367744 97928 367796 97980
rect 371884 97996 371936 98048
rect 395436 97928 395488 97980
rect 398196 97928 398248 97980
rect 165528 96568 165580 96620
rect 167000 96568 167052 96620
rect 394240 95140 394292 95192
rect 397460 95140 397512 95192
rect 392584 92420 392636 92472
rect 397460 92420 397512 92472
rect 364984 91060 365036 91112
rect 367744 91060 367796 91112
rect 395620 90992 395672 91044
rect 397920 90992 397972 91044
rect 392676 89632 392728 89684
rect 397460 89632 397512 89684
rect 395712 88272 395764 88324
rect 398840 88272 398892 88324
rect 395528 86912 395580 86964
rect 397736 86912 397788 86964
rect 544384 86912 544436 86964
rect 579988 86912 580040 86964
rect 395252 85484 395304 85536
rect 397552 85484 397604 85536
rect 360200 83988 360252 84040
rect 364984 83988 365036 84040
rect 392584 82084 392636 82136
rect 392952 82084 393004 82136
rect 397460 82084 397512 82136
rect 356704 81404 356756 81456
rect 360200 81404 360252 81456
rect 395896 79636 395948 79688
rect 398196 79636 398248 79688
rect 394332 78548 394384 78600
rect 397460 78548 397512 78600
rect 396908 75216 396960 75268
rect 398104 75216 398156 75268
rect 395436 71816 395488 71868
rect 397920 71816 397972 71868
rect 355324 68280 355376 68332
rect 356704 68280 356756 68332
rect 392676 66852 392728 66904
rect 393044 66852 393096 66904
rect 397460 66852 397512 66904
rect 165528 64948 165580 65000
rect 168288 64948 168340 65000
rect 280804 57196 280856 57248
rect 395988 57196 396040 57248
rect 397460 57196 397512 57248
rect 351920 56516 351972 56568
rect 355324 56584 355376 56636
rect 398012 56176 398064 56228
rect 399116 56176 399168 56228
rect 282184 54476 282236 54528
rect 397000 54476 397052 54528
rect 347504 53796 347556 53848
rect 351920 53796 351972 53848
rect 282828 51008 282880 51060
rect 347504 51008 347556 51060
rect 279424 48968 279476 49020
rect 397092 48968 397144 49020
rect 397460 48968 397512 49020
rect 282276 47540 282328 47592
rect 397460 47540 397512 47592
rect 398748 46860 398800 46912
rect 399024 46860 399076 46912
rect 518164 46860 518216 46912
rect 580172 46860 580224 46912
rect 168104 44140 168156 44192
rect 169024 44140 169076 44192
rect 280896 43392 280948 43444
rect 397184 43392 397236 43444
rect 167828 42032 167880 42084
rect 169208 42032 169260 42084
rect 167736 41692 167788 41744
rect 169116 41692 169168 41744
rect 279516 41420 279568 41472
rect 397460 41420 397512 41472
rect 280988 40672 281040 40724
rect 394516 40672 394568 40724
rect 397460 40672 397512 40724
rect 397736 40672 397788 40724
rect 398748 40672 398800 40724
rect 168012 39992 168064 40044
rect 169300 39992 169352 40044
rect 281080 39312 281132 39364
rect 397276 39312 397328 39364
rect 397460 39312 397512 39364
rect 278964 37272 279016 37324
rect 397552 37272 397604 37324
rect 167920 37204 167972 37256
rect 168932 37204 168984 37256
rect 509240 37204 509292 37256
rect 509516 37204 509568 37256
rect 281172 36524 281224 36576
rect 335360 36524 335412 36576
rect 279976 34484 280028 34536
rect 399760 34484 399812 34536
rect 168932 33464 168984 33516
rect 169576 33464 169628 33516
rect 168104 33260 168156 33312
rect 169668 33260 169720 33312
rect 279332 32376 279384 32428
rect 394608 32376 394660 32428
rect 397460 32376 397512 32428
rect 165528 31696 165580 31748
rect 398472 31696 398524 31748
rect 169392 31628 169444 31680
rect 398656 31628 398708 31680
rect 169484 31560 169536 31612
rect 398564 31560 398616 31612
rect 391940 31492 391992 31544
rect 393228 31492 393280 31544
rect 397460 31492 397512 31544
rect 280068 31016 280120 31068
rect 391940 31016 391992 31068
rect 169668 30268 169720 30320
rect 398104 30268 398156 30320
rect 169944 30200 169996 30252
rect 397736 30200 397788 30252
rect 169852 30132 169904 30184
rect 397920 30132 397972 30184
rect 169024 30064 169076 30116
rect 392584 30064 392636 30116
rect 168012 29996 168064 30048
rect 281080 29996 281132 30048
rect 167184 29928 167236 29980
rect 280896 29928 280948 29980
rect 168196 29860 168248 29912
rect 278964 29860 279016 29912
rect 167828 29792 167880 29844
rect 279516 29792 279568 29844
rect 170404 29724 170456 29776
rect 280068 29724 280120 29776
rect 168288 29656 168340 29708
rect 279976 29656 280028 29708
rect 167552 29588 167604 29640
rect 279424 29588 279476 29640
rect 446864 29248 446916 29300
rect 522304 29248 522356 29300
rect 438400 29180 438452 29232
rect 520924 29180 520976 29232
rect 208308 29112 208360 29164
rect 289084 29112 289136 29164
rect 429936 29112 429988 29164
rect 560944 29112 560996 29164
rect 216496 29044 216548 29096
rect 519544 29044 519596 29096
rect 183008 28976 183060 29028
rect 515404 28976 515456 29028
rect 169116 28908 169168 28960
rect 398380 28908 398432 28960
rect 506112 28908 506164 28960
rect 510712 28908 510764 28960
rect 167276 28840 167328 28892
rect 398196 28840 398248 28892
rect 497648 28840 497700 28892
rect 509424 28840 509476 28892
rect 169576 28772 169628 28824
rect 399208 28772 399260 28824
rect 413008 28772 413060 28824
rect 554044 28772 554096 28824
rect 168840 28704 168892 28756
rect 398288 28704 398340 28756
rect 421472 28704 421524 28756
rect 549904 28704 549956 28756
rect 395344 28636 395396 28688
rect 480352 28636 480404 28688
rect 489184 28636 489236 28688
rect 509332 28636 509384 28688
rect 395804 28568 395856 28620
rect 463148 28568 463200 28620
rect 169300 28500 169352 28552
rect 396724 28500 396776 28552
rect 404176 28500 404228 28552
rect 558184 28500 558236 28552
rect 169208 28432 169260 28484
rect 395436 28432 395488 28484
rect 169760 28364 169812 28416
rect 392676 28364 392728 28416
rect 28908 28296 28960 28348
rect 224960 28296 225012 28348
rect 250720 28296 250772 28348
rect 281172 28296 281224 28348
rect 307760 28296 307812 28348
rect 472072 28296 472124 28348
rect 259184 28228 259236 28280
rect 389824 28228 389876 28280
rect 167368 28160 167420 28212
rect 282184 28160 282236 28212
rect 167460 28092 167512 28144
rect 282276 28092 282328 28144
rect 171048 28024 171100 28076
rect 267004 28024 267056 28076
rect 275928 28024 275980 28076
rect 319444 28024 319496 28076
rect 174544 27956 174596 28008
rect 555424 27956 555476 28008
rect 168932 27888 168984 27940
rect 398012 27888 398064 27940
rect 284944 6808 284996 6860
rect 580172 6808 580224 6860
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 48042 536888 48098 536897
rect 396630 536888 396686 536897
rect 48042 536823 48098 536832
rect 242900 536852 242952 536858
rect 47950 533760 48006 533769
rect 47950 533695 48006 533704
rect 47858 531040 47914 531049
rect 47858 530975 47914 530984
rect 47766 508056 47822 508065
rect 47766 507991 47822 508000
rect 47780 429894 47808 507991
rect 47872 493338 47900 530975
rect 47964 496126 47992 533695
rect 47952 496120 48004 496126
rect 47952 496062 48004 496068
rect 47860 493332 47912 493338
rect 47860 493274 47912 493280
rect 48056 486470 48084 536823
rect 396630 536823 396632 536832
rect 242900 536794 242952 536800
rect 396684 536823 396686 536832
rect 396632 536794 396684 536800
rect 48226 535936 48282 535945
rect 48226 535871 48282 535880
rect 48134 532808 48190 532817
rect 48134 532743 48190 532752
rect 48148 498914 48176 532743
rect 48136 498908 48188 498914
rect 48136 498850 48188 498856
rect 48044 486464 48096 486470
rect 48044 486406 48096 486412
rect 47768 429888 47820 429894
rect 47768 429830 47820 429836
rect 1308 401668 1360 401674
rect 1308 401610 1360 401616
rect 1320 142730 1348 401610
rect 48240 400926 48268 535871
rect 237380 535492 237432 535498
rect 237380 535434 237432 535440
rect 231860 532840 231912 532846
rect 231860 532782 231912 532788
rect 226340 532772 226392 532778
rect 226340 532714 226392 532720
rect 222200 530052 222252 530058
rect 49514 529986 49570 529995
rect 222200 529994 222252 530000
rect 49514 529921 49570 529930
rect 213920 529984 213972 529990
rect 213920 529926 213972 529932
rect 49422 528218 49478 528227
rect 49422 528153 49478 528162
rect 49330 508328 49386 508337
rect 49330 508263 49386 508272
rect 49344 497826 49372 508263
rect 49436 498846 49464 528153
rect 49424 498840 49476 498846
rect 49424 498782 49476 498788
rect 49332 497820 49384 497826
rect 49332 497762 49384 497768
rect 49528 494766 49556 529921
rect 207020 527196 207072 527202
rect 207020 527138 207072 527144
rect 49606 509994 49662 510003
rect 49606 509929 49662 509938
rect 49516 494760 49568 494766
rect 49516 494702 49568 494708
rect 49620 428466 49648 509929
rect 191840 509312 191892 509318
rect 191840 509254 191892 509260
rect 190460 507884 190512 507890
rect 190460 507826 190512 507832
rect 177304 498908 177356 498914
rect 177304 498850 177356 498856
rect 67546 498128 67602 498137
rect 67546 498063 67602 498072
rect 73342 498128 73398 498137
rect 73342 498063 73398 498072
rect 74354 498128 74410 498137
rect 74354 498063 74410 498072
rect 78586 498128 78642 498137
rect 78586 498063 78642 498072
rect 79874 498128 79930 498137
rect 79874 498063 79930 498072
rect 81254 498128 81310 498137
rect 81254 498063 81310 498072
rect 85946 498128 86002 498137
rect 85946 498063 86002 498072
rect 86498 498128 86554 498137
rect 86498 498063 86554 498072
rect 89534 498128 89590 498137
rect 89534 498063 89590 498072
rect 92294 498128 92350 498137
rect 92294 498063 92350 498072
rect 96526 498128 96582 498137
rect 96526 498063 96582 498072
rect 103426 498128 103482 498137
rect 103426 498063 103482 498072
rect 104806 498128 104862 498137
rect 104806 498063 104862 498072
rect 113546 498128 113602 498137
rect 113546 498063 113602 498072
rect 116858 498128 116914 498137
rect 116858 498063 116914 498072
rect 118606 498128 118662 498137
rect 118606 498063 118662 498072
rect 121366 498128 121422 498137
rect 121366 498063 121422 498072
rect 126886 498128 126942 498137
rect 126886 498063 126942 498072
rect 129646 498128 129702 498137
rect 129646 498063 129702 498072
rect 146206 498128 146262 498137
rect 146206 498063 146262 498072
rect 150990 498128 151046 498137
rect 150990 498063 151046 498072
rect 154486 498128 154542 498137
rect 154486 498063 154542 498072
rect 53840 497820 53892 497826
rect 53840 497762 53892 497768
rect 49608 428460 49660 428466
rect 49608 428402 49660 428408
rect 53852 401674 53880 497762
rect 66166 496904 66222 496913
rect 66166 496839 66222 496848
rect 66180 406434 66208 496839
rect 67560 428534 67588 498063
rect 73066 497448 73122 497457
rect 73066 497383 73122 497392
rect 68926 496904 68982 496913
rect 68926 496839 68982 496848
rect 70306 496904 70362 496913
rect 70306 496839 70362 496848
rect 71686 496904 71742 496913
rect 71686 496839 71742 496848
rect 67548 428528 67600 428534
rect 67548 428470 67600 428476
rect 68940 423434 68968 496839
rect 70320 423502 70348 496839
rect 71700 423570 71728 496839
rect 73080 423638 73108 497383
rect 73356 496874 73384 498063
rect 73344 496868 73396 496874
rect 73344 496810 73396 496816
rect 74368 487830 74396 498063
rect 75826 496904 75882 496913
rect 75184 496868 75236 496874
rect 75826 496839 75882 496848
rect 77206 496904 77262 496913
rect 77206 496839 77262 496848
rect 78310 496904 78366 496913
rect 78310 496839 78312 496848
rect 75184 496810 75236 496816
rect 74356 487824 74408 487830
rect 74356 487766 74408 487772
rect 75196 482322 75224 496810
rect 75184 482316 75236 482322
rect 75184 482258 75236 482264
rect 73068 423632 73120 423638
rect 73068 423574 73120 423580
rect 71688 423564 71740 423570
rect 71688 423506 71740 423512
rect 70308 423496 70360 423502
rect 70308 423438 70360 423444
rect 68928 423428 68980 423434
rect 68928 423370 68980 423376
rect 75840 416090 75868 496839
rect 77220 474026 77248 496839
rect 78364 496839 78366 496848
rect 78312 496810 78364 496816
rect 77208 474020 77260 474026
rect 77208 473962 77260 473968
rect 78600 424386 78628 498063
rect 79888 496942 79916 498063
rect 81162 497040 81218 497049
rect 81268 497010 81296 498063
rect 85960 497214 85988 498063
rect 85948 497208 86000 497214
rect 85948 497150 86000 497156
rect 86512 497078 86540 498063
rect 89548 497282 89576 498063
rect 92308 497350 92336 498063
rect 96342 497856 96398 497865
rect 96342 497791 96398 497800
rect 92296 497344 92348 497350
rect 92296 497286 92348 497292
rect 89536 497276 89588 497282
rect 89536 497218 89588 497224
rect 86500 497072 86552 497078
rect 84014 497040 84070 497049
rect 81162 496975 81218 496984
rect 81256 497004 81308 497010
rect 79876 496936 79928 496942
rect 79876 496878 79928 496884
rect 79324 496868 79376 496874
rect 79324 496810 79376 496816
rect 78588 424380 78640 424386
rect 78588 424322 78640 424328
rect 79336 423026 79364 496810
rect 81176 434042 81204 496975
rect 86500 497014 86552 497020
rect 88154 497040 88210 497049
rect 84014 496975 84070 496984
rect 88154 496975 88210 496984
rect 93674 497040 93730 497049
rect 93674 496975 93730 496984
rect 81256 496946 81308 496952
rect 81254 496904 81310 496913
rect 81254 496839 81310 496848
rect 82726 496904 82782 496913
rect 82726 496839 82782 496848
rect 81268 472666 81296 496839
rect 81256 472660 81308 472666
rect 81256 472602 81308 472608
rect 81164 434036 81216 434042
rect 81164 433978 81216 433984
rect 82740 432614 82768 496839
rect 82728 432608 82780 432614
rect 82728 432550 82780 432556
rect 84028 427106 84056 496975
rect 84106 496904 84162 496913
rect 84106 496839 84162 496848
rect 85486 496904 85542 496913
rect 85486 496839 85542 496848
rect 84016 427100 84068 427106
rect 84016 427042 84068 427048
rect 79324 423020 79376 423026
rect 79324 422962 79376 422968
rect 75828 416084 75880 416090
rect 75828 416026 75880 416032
rect 66168 406428 66220 406434
rect 66168 406370 66220 406376
rect 84120 405006 84148 496839
rect 85500 435402 85528 496839
rect 88168 489190 88196 496975
rect 88246 496904 88302 496913
rect 88246 496839 88302 496848
rect 89166 496904 89222 496913
rect 89166 496839 89222 496848
rect 91006 496904 91062 496913
rect 91006 496839 91062 496848
rect 91190 496904 91246 496913
rect 91190 496839 91246 496848
rect 88156 489184 88208 489190
rect 88156 489126 88208 489132
rect 88260 436762 88288 496839
rect 89180 491978 89208 496839
rect 89168 491972 89220 491978
rect 89168 491914 89220 491920
rect 88248 436756 88300 436762
rect 88248 436698 88300 436704
rect 85488 435396 85540 435402
rect 85488 435338 85540 435344
rect 91020 407794 91048 496839
rect 91204 490618 91232 496839
rect 91192 490612 91244 490618
rect 91192 490554 91244 490560
rect 93688 445058 93716 496975
rect 93766 496904 93822 496913
rect 93766 496839 93822 496848
rect 95146 496904 95202 496913
rect 95146 496839 95202 496848
rect 93676 445052 93728 445058
rect 93676 444994 93728 445000
rect 93780 429962 93808 496839
rect 93768 429956 93820 429962
rect 93768 429898 93820 429904
rect 95160 409154 95188 496839
rect 96356 496194 96384 497791
rect 96434 497040 96490 497049
rect 96434 496975 96490 496984
rect 96344 496188 96396 496194
rect 96344 496130 96396 496136
rect 96448 485110 96476 496975
rect 96436 485104 96488 485110
rect 96436 485046 96488 485052
rect 96540 431254 96568 498063
rect 99286 497040 99342 497049
rect 99286 496975 99342 496984
rect 101954 497040 102010 497049
rect 101954 496975 102010 496984
rect 97906 496904 97962 496913
rect 97906 496839 97962 496848
rect 99194 496904 99250 496913
rect 99194 496839 99250 496848
rect 97920 442270 97948 496839
rect 99208 443698 99236 496839
rect 99196 443692 99248 443698
rect 99196 443634 99248 443640
rect 97908 442264 97960 442270
rect 97908 442206 97960 442212
rect 99300 440910 99328 496975
rect 100666 496904 100722 496913
rect 100666 496839 100722 496848
rect 100680 446418 100708 496839
rect 101968 486538 101996 496975
rect 102046 496904 102102 496913
rect 102046 496839 102102 496848
rect 103334 496904 103390 496913
rect 103440 496874 103468 498063
rect 104714 496904 104770 496913
rect 103334 496839 103390 496848
rect 103428 496868 103480 496874
rect 101956 486532 102008 486538
rect 101956 486474 102008 486480
rect 102060 447846 102088 496839
rect 103348 449206 103376 496839
rect 104714 496839 104770 496848
rect 103428 496810 103480 496816
rect 104728 480962 104756 496839
rect 104716 480956 104768 480962
rect 104716 480898 104768 480904
rect 103336 449200 103388 449206
rect 103336 449142 103388 449148
rect 102048 447840 102100 447846
rect 102048 447782 102100 447788
rect 100668 446412 100720 446418
rect 100668 446354 100720 446360
rect 99288 440904 99340 440910
rect 99288 440846 99340 440852
rect 104820 439550 104848 498063
rect 113560 497418 113588 498063
rect 116872 497486 116900 498063
rect 116860 497480 116912 497486
rect 116860 497422 116912 497428
rect 113548 497412 113600 497418
rect 113548 497354 113600 497360
rect 118620 497146 118648 498063
rect 118608 497140 118660 497146
rect 118608 497082 118660 497088
rect 106094 497040 106150 497049
rect 106094 496975 106150 496984
rect 108854 497040 108910 497049
rect 108854 496975 108910 496984
rect 106108 493406 106136 496975
rect 106186 496904 106242 496913
rect 106186 496839 106242 496848
rect 107566 496904 107622 496913
rect 107566 496839 107622 496848
rect 106096 493400 106148 493406
rect 106096 493342 106148 493348
rect 104808 439544 104860 439550
rect 104808 439486 104860 439492
rect 96528 431248 96580 431254
rect 96528 431190 96580 431196
rect 106200 413302 106228 496839
rect 107580 419490 107608 496839
rect 108868 476814 108896 496975
rect 108946 496904 109002 496913
rect 108946 496839 109002 496848
rect 110326 496904 110382 496913
rect 110326 496839 110382 496848
rect 111706 496904 111762 496913
rect 111706 496839 111762 496848
rect 108856 476808 108908 476814
rect 108856 476750 108908 476756
rect 108960 431322 108988 496839
rect 110340 478174 110368 496839
rect 110328 478168 110380 478174
rect 110328 478110 110380 478116
rect 111720 432682 111748 496839
rect 111708 432676 111760 432682
rect 111708 432618 111760 432624
rect 108948 431316 109000 431322
rect 108948 431258 109000 431264
rect 107568 419484 107620 419490
rect 107568 419426 107620 419432
rect 106188 413296 106240 413302
rect 106188 413238 106240 413244
rect 95148 409148 95200 409154
rect 95148 409090 95200 409096
rect 91008 407788 91060 407794
rect 91008 407730 91060 407736
rect 84108 405000 84160 405006
rect 84108 404942 84160 404948
rect 53840 401668 53892 401674
rect 53840 401610 53892 401616
rect 54944 401668 54996 401674
rect 54944 401610 54996 401616
rect 104900 401668 104952 401674
rect 104900 401610 104952 401616
rect 48228 400920 48280 400926
rect 48228 400862 48280 400868
rect 54956 399976 54984 401610
rect 104912 399976 104940 401610
rect 121380 401606 121408 498063
rect 124126 496904 124182 496913
rect 124126 496839 124182 496848
rect 124140 404326 124168 496839
rect 126900 422958 126928 498063
rect 126888 422952 126940 422958
rect 126888 422894 126940 422900
rect 129660 407114 129688 498063
rect 133144 497480 133196 497486
rect 133144 497422 133196 497428
rect 131856 497412 131908 497418
rect 131856 497354 131908 497360
rect 131764 497344 131816 497350
rect 131764 497286 131816 497292
rect 130476 497276 130528 497282
rect 130476 497218 130528 497224
rect 130384 497208 130436 497214
rect 130384 497150 130436 497156
rect 129648 407108 129700 407114
rect 129648 407050 129700 407056
rect 124128 404320 124180 404326
rect 124128 404262 124180 404268
rect 121368 401600 121420 401606
rect 121368 401542 121420 401548
rect 28906 350024 28962 350033
rect 28906 349959 28962 349968
rect 20 142724 72 142730
rect 20 142666 72 142672
rect 1308 142724 1360 142730
rect 1308 142666 1360 142672
rect 32 16574 60 142666
rect 1320 142254 1348 142666
rect 1308 142248 1360 142254
rect 1308 142190 1360 142196
rect 1400 142180 1452 142186
rect 1400 142122 1452 142128
rect 32 16546 152 16574
rect 124 354 152 16546
rect 542 354 654 480
rect 124 326 654 354
rect 1412 354 1440 142122
rect 28920 28354 28948 349959
rect 78692 300002 79994 300030
rect 78692 28937 78720 300002
rect 130396 196994 130424 497150
rect 130488 197062 130516 497218
rect 131026 496904 131082 496913
rect 131026 496839 131082 496848
rect 131040 197198 131068 496839
rect 131210 399120 131266 399129
rect 131210 399055 131266 399064
rect 131224 398886 131252 399055
rect 131212 398880 131264 398886
rect 131212 398822 131264 398828
rect 131210 398576 131266 398585
rect 131210 398511 131266 398520
rect 131224 397526 131252 398511
rect 131212 397520 131264 397526
rect 131212 397462 131264 397468
rect 131486 397352 131542 397361
rect 131486 397287 131542 397296
rect 131302 396808 131358 396817
rect 131302 396743 131358 396752
rect 131210 396264 131266 396273
rect 131210 396199 131212 396208
rect 131264 396199 131266 396208
rect 131212 396170 131264 396176
rect 131316 396098 131344 396743
rect 131500 396166 131528 397287
rect 131488 396160 131540 396166
rect 131488 396102 131540 396108
rect 131304 396092 131356 396098
rect 131304 396034 131356 396040
rect 131210 395584 131266 395593
rect 131210 395519 131266 395528
rect 131224 394806 131252 395519
rect 131302 395040 131358 395049
rect 131302 394975 131358 394984
rect 131212 394800 131264 394806
rect 131212 394742 131264 394748
rect 131316 394738 131344 394975
rect 131304 394732 131356 394738
rect 131304 394674 131356 394680
rect 131210 394496 131266 394505
rect 131210 394431 131266 394440
rect 131224 393446 131252 394431
rect 131212 393440 131264 393446
rect 131212 393382 131264 393388
rect 131210 393272 131266 393281
rect 131210 393207 131266 393216
rect 131224 392018 131252 393207
rect 131302 392184 131358 392193
rect 131302 392119 131358 392128
rect 131212 392012 131264 392018
rect 131212 391954 131264 391960
rect 131210 391504 131266 391513
rect 131210 391439 131266 391448
rect 131224 390658 131252 391439
rect 131212 390652 131264 390658
rect 131212 390594 131264 390600
rect 131118 390416 131174 390425
rect 131118 390351 131174 390360
rect 131132 389366 131160 390351
rect 131316 389842 131344 392119
rect 131486 390960 131542 390969
rect 131486 390895 131542 390904
rect 131500 390590 131528 390895
rect 131488 390584 131540 390590
rect 131488 390526 131540 390532
rect 131486 389872 131542 389881
rect 131304 389836 131356 389842
rect 131486 389807 131542 389816
rect 131304 389778 131356 389784
rect 131120 389360 131172 389366
rect 131120 389302 131172 389308
rect 131212 389292 131264 389298
rect 131212 389234 131264 389240
rect 131224 389201 131252 389234
rect 131500 389230 131528 389807
rect 131488 389224 131540 389230
rect 131210 389192 131266 389201
rect 131488 389166 131540 389172
rect 131210 389127 131266 389136
rect 131302 388648 131358 388657
rect 131302 388583 131358 388592
rect 131210 388104 131266 388113
rect 131210 388039 131266 388048
rect 131224 387938 131252 388039
rect 131212 387932 131264 387938
rect 131212 387874 131264 387880
rect 131316 387870 131344 388583
rect 131304 387864 131356 387870
rect 131304 387806 131356 387812
rect 131118 387424 131174 387433
rect 131118 387359 131174 387368
rect 131132 386442 131160 387359
rect 131210 386880 131266 386889
rect 131210 386815 131266 386824
rect 131224 386646 131252 386815
rect 131212 386640 131264 386646
rect 131212 386582 131264 386588
rect 131120 386436 131172 386442
rect 131120 386378 131172 386384
rect 131302 386336 131358 386345
rect 131302 386271 131358 386280
rect 131118 385792 131174 385801
rect 131118 385727 131174 385736
rect 131132 385218 131160 385727
rect 131120 385212 131172 385218
rect 131120 385154 131172 385160
rect 131212 385144 131264 385150
rect 131210 385112 131212 385121
rect 131264 385112 131266 385121
rect 131316 385082 131344 386271
rect 131210 385047 131266 385056
rect 131304 385076 131356 385082
rect 131304 385018 131356 385024
rect 131118 384568 131174 384577
rect 131118 384503 131174 384512
rect 131132 383722 131160 384503
rect 131210 384024 131266 384033
rect 131210 383959 131266 383968
rect 131224 383790 131252 383959
rect 131212 383784 131264 383790
rect 131212 383726 131264 383732
rect 131120 383716 131172 383722
rect 131120 383658 131172 383664
rect 131118 383480 131174 383489
rect 131118 383415 131174 383424
rect 131132 382362 131160 383415
rect 131210 382800 131266 382809
rect 131210 382735 131266 382744
rect 131120 382356 131172 382362
rect 131120 382298 131172 382304
rect 131224 382294 131252 382735
rect 131212 382288 131264 382294
rect 131212 382230 131264 382236
rect 131486 382256 131542 382265
rect 131486 382191 131542 382200
rect 131210 381032 131266 381041
rect 131210 380967 131212 380976
rect 131264 380967 131266 380976
rect 131212 380938 131264 380944
rect 131500 380934 131528 382191
rect 131488 380928 131540 380934
rect 131488 380870 131540 380876
rect 131210 380488 131266 380497
rect 131210 380423 131266 380432
rect 131224 379642 131252 380423
rect 131486 379944 131542 379953
rect 131486 379879 131542 379888
rect 131212 379636 131264 379642
rect 131212 379578 131264 379584
rect 131500 379574 131528 379879
rect 131488 379568 131540 379574
rect 131488 379510 131540 379516
rect 131118 379400 131174 379409
rect 131118 379335 131174 379344
rect 131132 378350 131160 379335
rect 131302 378720 131358 378729
rect 131302 378655 131358 378664
rect 131120 378344 131172 378350
rect 131120 378286 131172 378292
rect 131212 378276 131264 378282
rect 131212 378218 131264 378224
rect 131224 378185 131252 378218
rect 131316 378214 131344 378655
rect 131304 378208 131356 378214
rect 131210 378176 131266 378185
rect 131304 378150 131356 378156
rect 131210 378111 131266 378120
rect 131118 377632 131174 377641
rect 131118 377567 131174 377576
rect 131132 376786 131160 377567
rect 131210 377088 131266 377097
rect 131210 377023 131266 377032
rect 131224 376854 131252 377023
rect 131212 376848 131264 376854
rect 131212 376790 131264 376796
rect 131120 376780 131172 376786
rect 131120 376722 131172 376728
rect 131210 376408 131266 376417
rect 131210 376343 131266 376352
rect 131224 375426 131252 376343
rect 131486 375864 131542 375873
rect 131486 375799 131542 375808
rect 131500 375494 131528 375799
rect 131488 375488 131540 375494
rect 131488 375430 131540 375436
rect 131212 375420 131264 375426
rect 131212 375362 131264 375368
rect 131210 375320 131266 375329
rect 131210 375255 131266 375264
rect 131118 374640 131174 374649
rect 131118 374575 131174 374584
rect 131132 374134 131160 374575
rect 131224 374202 131252 375255
rect 131212 374196 131264 374202
rect 131212 374138 131264 374144
rect 131120 374128 131172 374134
rect 131120 374070 131172 374076
rect 131210 374096 131266 374105
rect 131210 374031 131212 374040
rect 131264 374031 131266 374040
rect 131212 374002 131264 374008
rect 131210 373552 131266 373561
rect 131210 373487 131266 373496
rect 131224 372706 131252 373487
rect 131486 373008 131542 373017
rect 131486 372943 131542 372952
rect 131212 372700 131264 372706
rect 131212 372642 131264 372648
rect 131500 372638 131528 372943
rect 131488 372632 131540 372638
rect 131488 372574 131540 372580
rect 131118 372328 131174 372337
rect 131118 372263 131174 372272
rect 131132 371278 131160 372263
rect 131210 371784 131266 371793
rect 131210 371719 131266 371728
rect 131224 371346 131252 371719
rect 131212 371340 131264 371346
rect 131212 371282 131264 371288
rect 131120 371272 131172 371278
rect 131120 371214 131172 371220
rect 131118 370696 131174 370705
rect 131118 370631 131174 370640
rect 131132 369918 131160 370631
rect 131210 370016 131266 370025
rect 131210 369951 131212 369960
rect 131264 369951 131266 369960
rect 131212 369922 131264 369928
rect 131120 369912 131172 369918
rect 131120 369854 131172 369860
rect 131210 369472 131266 369481
rect 131210 369407 131266 369416
rect 131224 368558 131252 369407
rect 131486 368928 131542 368937
rect 131486 368863 131542 368872
rect 131500 368626 131528 368863
rect 131488 368620 131540 368626
rect 131488 368562 131540 368568
rect 131212 368552 131264 368558
rect 131212 368494 131264 368500
rect 131210 368248 131266 368257
rect 131210 368183 131266 368192
rect 131118 367704 131174 367713
rect 131118 367639 131174 367648
rect 131132 367198 131160 367639
rect 131224 367266 131252 368183
rect 131212 367260 131264 367266
rect 131212 367202 131264 367208
rect 131120 367192 131172 367198
rect 131120 367134 131172 367140
rect 131210 367160 131266 367169
rect 131210 367095 131212 367104
rect 131264 367095 131266 367104
rect 131212 367066 131264 367072
rect 131210 365936 131266 365945
rect 131210 365871 131266 365880
rect 131224 365770 131252 365871
rect 131212 365764 131264 365770
rect 131212 365706 131264 365712
rect 131118 365392 131174 365401
rect 131118 365327 131174 365336
rect 131132 364478 131160 365327
rect 131210 364848 131266 364857
rect 131210 364783 131266 364792
rect 131120 364472 131172 364478
rect 131120 364414 131172 364420
rect 131224 364410 131252 364783
rect 131212 364404 131264 364410
rect 131212 364346 131264 364352
rect 131486 364304 131542 364313
rect 131486 364239 131542 364248
rect 131118 363624 131174 363633
rect 131118 363559 131174 363568
rect 131132 363118 131160 363559
rect 131120 363112 131172 363118
rect 131120 363054 131172 363060
rect 131210 363080 131266 363089
rect 131210 363015 131212 363024
rect 131264 363015 131266 363024
rect 131212 362986 131264 362992
rect 131500 362982 131528 364239
rect 131488 362976 131540 362982
rect 131488 362918 131540 362924
rect 131118 362536 131174 362545
rect 131118 362471 131174 362480
rect 131132 361622 131160 362471
rect 131210 361856 131266 361865
rect 131210 361791 131266 361800
rect 131224 361690 131252 361791
rect 131212 361684 131264 361690
rect 131212 361626 131264 361632
rect 131120 361616 131172 361622
rect 131120 361558 131172 361564
rect 131118 361312 131174 361321
rect 131118 361247 131174 361256
rect 131132 360330 131160 361247
rect 131120 360324 131172 360330
rect 131120 360266 131172 360272
rect 131212 360256 131264 360262
rect 131210 360224 131212 360233
rect 131264 360224 131266 360233
rect 131210 360159 131266 360168
rect 131210 359000 131266 359009
rect 131210 358935 131266 358944
rect 131224 358834 131252 358935
rect 131212 358828 131264 358834
rect 131212 358770 131264 358776
rect 131118 358456 131174 358465
rect 131118 358391 131174 358400
rect 131132 357542 131160 358391
rect 131210 357912 131266 357921
rect 131210 357847 131266 357856
rect 131120 357536 131172 357542
rect 131120 357478 131172 357484
rect 131224 357474 131252 357847
rect 131212 357468 131264 357474
rect 131212 357410 131264 357416
rect 131302 357232 131358 357241
rect 131302 357167 131358 357176
rect 131118 356688 131174 356697
rect 131118 356623 131174 356632
rect 131132 356182 131160 356623
rect 131212 356244 131264 356250
rect 131212 356186 131264 356192
rect 131120 356176 131172 356182
rect 131224 356153 131252 356186
rect 131120 356118 131172 356124
rect 131210 356144 131266 356153
rect 131316 356114 131344 357167
rect 131210 356079 131266 356088
rect 131304 356108 131356 356114
rect 131304 356050 131356 356056
rect 131302 355464 131358 355473
rect 131302 355399 131358 355408
rect 131210 354920 131266 354929
rect 131210 354855 131266 354864
rect 131224 354822 131252 354855
rect 131212 354816 131264 354822
rect 131212 354758 131264 354764
rect 131316 354754 131344 355399
rect 131304 354748 131356 354754
rect 131304 354690 131356 354696
rect 131118 354376 131174 354385
rect 131118 354311 131174 354320
rect 131132 353326 131160 354311
rect 131210 353832 131266 353841
rect 131210 353767 131266 353776
rect 131224 353394 131252 353767
rect 131212 353388 131264 353394
rect 131212 353330 131264 353336
rect 131120 353320 131172 353326
rect 131120 353262 131172 353268
rect 131210 353152 131266 353161
rect 131210 353087 131266 353096
rect 131118 352608 131174 352617
rect 131118 352543 131174 352552
rect 131132 352034 131160 352543
rect 131224 352102 131252 353087
rect 131212 352096 131264 352102
rect 131212 352038 131264 352044
rect 131486 352064 131542 352073
rect 131120 352028 131172 352034
rect 131486 351999 131542 352008
rect 131120 351970 131172 351976
rect 131500 351966 131528 351999
rect 131488 351960 131540 351966
rect 131488 351902 131540 351908
rect 131118 351520 131174 351529
rect 131118 351455 131174 351464
rect 131132 350674 131160 351455
rect 131210 350840 131266 350849
rect 131210 350775 131266 350784
rect 131120 350668 131172 350674
rect 131120 350610 131172 350616
rect 131224 350606 131252 350775
rect 131212 350600 131264 350606
rect 131212 350542 131264 350548
rect 131118 350296 131174 350305
rect 131118 350231 131174 350240
rect 131132 349178 131160 350231
rect 131210 349752 131266 349761
rect 131210 349687 131266 349696
rect 131224 349246 131252 349687
rect 131212 349240 131264 349246
rect 131212 349182 131264 349188
rect 131120 349172 131172 349178
rect 131120 349114 131172 349120
rect 131210 349072 131266 349081
rect 131210 349007 131266 349016
rect 131224 348362 131252 349007
rect 131302 348528 131358 348537
rect 131302 348463 131358 348472
rect 131212 348356 131264 348362
rect 131212 348298 131264 348304
rect 131316 347818 131344 348463
rect 131486 347984 131542 347993
rect 131486 347919 131542 347928
rect 131500 347886 131528 347919
rect 131488 347880 131540 347886
rect 131488 347822 131540 347828
rect 131304 347812 131356 347818
rect 131304 347754 131356 347760
rect 131118 347440 131174 347449
rect 131118 347375 131174 347384
rect 131132 346458 131160 347375
rect 131210 346760 131266 346769
rect 131210 346695 131266 346704
rect 131224 346526 131252 346695
rect 131212 346520 131264 346526
rect 131212 346462 131264 346468
rect 131120 346452 131172 346458
rect 131120 346394 131172 346400
rect 131210 346216 131266 346225
rect 131210 346151 131266 346160
rect 131118 345672 131174 345681
rect 131118 345607 131174 345616
rect 131132 345166 131160 345607
rect 131224 345234 131252 346151
rect 131212 345228 131264 345234
rect 131212 345170 131264 345176
rect 131120 345160 131172 345166
rect 131120 345102 131172 345108
rect 131210 345128 131266 345137
rect 131210 345063 131212 345072
rect 131264 345063 131266 345072
rect 131212 345034 131264 345040
rect 131302 344448 131358 344457
rect 131302 344383 131358 344392
rect 131210 343904 131266 343913
rect 131210 343839 131266 343848
rect 131224 343670 131252 343839
rect 131316 343738 131344 344383
rect 131304 343732 131356 343738
rect 131304 343674 131356 343680
rect 131212 343664 131264 343670
rect 131212 343606 131264 343612
rect 131210 343360 131266 343369
rect 131210 343295 131266 343304
rect 131224 342378 131252 343295
rect 131486 342680 131542 342689
rect 131486 342615 131542 342624
rect 131212 342372 131264 342378
rect 131212 342314 131264 342320
rect 131500 342310 131528 342615
rect 131488 342304 131540 342310
rect 131488 342246 131540 342252
rect 131118 342136 131174 342145
rect 131118 342071 131174 342080
rect 131132 340950 131160 342071
rect 131302 341592 131358 341601
rect 131302 341527 131358 341536
rect 131212 341080 131264 341086
rect 131210 341048 131212 341057
rect 131264 341048 131266 341057
rect 131316 341018 131344 341527
rect 131210 340983 131266 340992
rect 131304 341012 131356 341018
rect 131304 340954 131356 340960
rect 131120 340944 131172 340950
rect 131120 340886 131172 340892
rect 131302 340368 131358 340377
rect 131302 340303 131358 340312
rect 131210 339824 131266 339833
rect 131210 339759 131266 339768
rect 131224 339522 131252 339759
rect 131316 339590 131344 340303
rect 131304 339584 131356 339590
rect 131304 339526 131356 339532
rect 131212 339516 131264 339522
rect 131212 339458 131264 339464
rect 131118 339280 131174 339289
rect 131118 339215 131174 339224
rect 131132 338162 131160 339215
rect 131210 338736 131266 338745
rect 131210 338671 131266 338680
rect 131224 338230 131252 338671
rect 131212 338224 131264 338230
rect 131212 338166 131264 338172
rect 131120 338156 131172 338162
rect 131120 338098 131172 338104
rect 131486 338056 131542 338065
rect 131486 337991 131542 338000
rect 131210 336968 131266 336977
rect 131210 336903 131212 336912
rect 131264 336903 131266 336912
rect 131212 336874 131264 336880
rect 131500 336802 131528 337991
rect 131488 336796 131540 336802
rect 131488 336738 131540 336744
rect 131118 336288 131174 336297
rect 131118 336223 131174 336232
rect 131132 335374 131160 336223
rect 131210 335744 131266 335753
rect 131210 335679 131266 335688
rect 131224 335442 131252 335679
rect 131212 335436 131264 335442
rect 131212 335378 131264 335384
rect 131120 335368 131172 335374
rect 131120 335310 131172 335316
rect 131210 335200 131266 335209
rect 131210 335135 131266 335144
rect 131224 334014 131252 335135
rect 131212 334008 131264 334014
rect 131118 333976 131174 333985
rect 131212 333950 131264 333956
rect 131118 333911 131174 333920
rect 131132 332790 131160 333911
rect 131302 333432 131358 333441
rect 131302 333367 131358 333376
rect 131210 332888 131266 332897
rect 131210 332823 131266 332832
rect 131120 332784 131172 332790
rect 131120 332726 131172 332732
rect 131224 332654 131252 332823
rect 131316 332722 131344 333367
rect 131304 332716 131356 332722
rect 131304 332658 131356 332664
rect 131212 332648 131264 332654
rect 131212 332590 131264 332596
rect 131486 331664 131542 331673
rect 131486 331599 131542 331608
rect 131500 331294 131528 331599
rect 131488 331288 131540 331294
rect 131488 331230 131540 331236
rect 131118 331120 131174 331129
rect 131118 331055 131174 331064
rect 131132 329934 131160 331055
rect 131120 329928 131172 329934
rect 131120 329870 131172 329876
rect 131210 329896 131266 329905
rect 131210 329831 131212 329840
rect 131264 329831 131266 329840
rect 131212 329802 131264 329808
rect 131210 329352 131266 329361
rect 131210 329287 131266 329296
rect 131224 328574 131252 329287
rect 131302 328808 131358 328817
rect 131302 328743 131358 328752
rect 131212 328568 131264 328574
rect 131212 328510 131264 328516
rect 131316 328506 131344 328743
rect 131304 328500 131356 328506
rect 131304 328442 131356 328448
rect 131118 328264 131174 328273
rect 131118 328199 131174 328208
rect 131132 327214 131160 328199
rect 131210 327584 131266 327593
rect 131210 327519 131266 327528
rect 131120 327208 131172 327214
rect 131120 327150 131172 327156
rect 131224 327146 131252 327519
rect 131212 327140 131264 327146
rect 131212 327082 131264 327088
rect 131302 326496 131358 326505
rect 131302 326431 131358 326440
rect 131210 325952 131266 325961
rect 131210 325887 131266 325896
rect 131224 325786 131252 325887
rect 131212 325780 131264 325786
rect 131212 325722 131264 325728
rect 131316 325718 131344 326431
rect 131304 325712 131356 325718
rect 131304 325654 131356 325660
rect 131210 325272 131266 325281
rect 131210 325207 131266 325216
rect 131224 324358 131252 325207
rect 131486 324728 131542 324737
rect 131486 324663 131542 324672
rect 131500 324426 131528 324663
rect 131488 324420 131540 324426
rect 131488 324362 131540 324368
rect 131212 324352 131264 324358
rect 131212 324294 131264 324300
rect 131118 324184 131174 324193
rect 131118 324119 131174 324128
rect 131132 323066 131160 324119
rect 131486 323504 131542 323513
rect 131486 323439 131542 323448
rect 131500 323134 131528 323439
rect 131488 323128 131540 323134
rect 131488 323070 131540 323076
rect 131120 323060 131172 323066
rect 131120 323002 131172 323008
rect 131212 322992 131264 322998
rect 131210 322960 131212 322969
rect 131264 322960 131266 322969
rect 131210 322895 131266 322904
rect 131118 322416 131174 322425
rect 131118 322351 131174 322360
rect 131132 321638 131160 322351
rect 131210 321872 131266 321881
rect 131210 321807 131266 321816
rect 131224 321706 131252 321807
rect 131212 321700 131264 321706
rect 131212 321642 131264 321648
rect 131120 321632 131172 321638
rect 131120 321574 131172 321580
rect 131118 321192 131174 321201
rect 131118 321127 131174 321136
rect 131132 320278 131160 321127
rect 131210 320648 131266 320657
rect 131210 320583 131266 320592
rect 131120 320272 131172 320278
rect 131120 320214 131172 320220
rect 131224 320210 131252 320583
rect 131212 320204 131264 320210
rect 131212 320146 131264 320152
rect 131210 318880 131266 318889
rect 131210 318815 131212 318824
rect 131264 318815 131266 318824
rect 131212 318786 131264 318792
rect 131486 317792 131542 317801
rect 131486 317727 131542 317736
rect 131500 317490 131528 317727
rect 131488 317484 131540 317490
rect 131488 317426 131540 317432
rect 131210 316568 131266 316577
rect 131210 316503 131266 316512
rect 131224 316062 131252 316503
rect 131212 316056 131264 316062
rect 131212 315998 131264 316004
rect 131486 316024 131542 316033
rect 131486 315959 131542 315968
rect 131210 315480 131266 315489
rect 131210 315415 131266 315424
rect 131224 314702 131252 315415
rect 131302 314800 131358 314809
rect 131500 314770 131528 315959
rect 131302 314735 131358 314744
rect 131488 314764 131540 314770
rect 131212 314696 131264 314702
rect 131212 314638 131264 314644
rect 131118 314256 131174 314265
rect 131118 314191 131174 314200
rect 131132 313342 131160 314191
rect 131316 313954 131344 314735
rect 131488 314706 131540 314712
rect 131304 313948 131356 313954
rect 131304 313890 131356 313896
rect 131210 313712 131266 313721
rect 131210 313647 131266 313656
rect 131224 313410 131252 313647
rect 131212 313404 131264 313410
rect 131212 313346 131264 313352
rect 131120 313336 131172 313342
rect 131120 313278 131172 313284
rect 131302 313168 131358 313177
rect 131302 313103 131358 313112
rect 131118 312488 131174 312497
rect 131118 312423 131174 312432
rect 131132 311982 131160 312423
rect 131120 311976 131172 311982
rect 131120 311918 131172 311924
rect 131210 311944 131266 311953
rect 131210 311879 131212 311888
rect 131264 311879 131266 311888
rect 131212 311850 131264 311856
rect 131210 311400 131266 311409
rect 131210 311335 131266 311344
rect 131224 310554 131252 311335
rect 131212 310548 131264 310554
rect 131212 310490 131264 310496
rect 131118 310176 131174 310185
rect 131118 310111 131174 310120
rect 131132 309670 131160 310111
rect 131316 309806 131344 313103
rect 131486 310720 131542 310729
rect 131486 310655 131542 310664
rect 131500 310622 131528 310655
rect 131488 310616 131540 310622
rect 131488 310558 131540 310564
rect 131304 309800 131356 309806
rect 131304 309742 131356 309748
rect 131120 309664 131172 309670
rect 131120 309606 131172 309612
rect 131210 309632 131266 309641
rect 131210 309567 131266 309576
rect 131224 309194 131252 309567
rect 131212 309188 131264 309194
rect 131212 309130 131264 309136
rect 131118 309088 131174 309097
rect 131118 309023 131174 309032
rect 131132 307902 131160 309023
rect 131486 308408 131542 308417
rect 131486 308343 131542 308352
rect 131212 307964 131264 307970
rect 131212 307906 131264 307912
rect 131120 307896 131172 307902
rect 131224 307873 131252 307906
rect 131120 307838 131172 307844
rect 131210 307864 131266 307873
rect 131500 307834 131528 308343
rect 131210 307799 131266 307808
rect 131488 307828 131540 307834
rect 131488 307770 131540 307776
rect 131118 307320 131174 307329
rect 131118 307255 131174 307264
rect 131132 306474 131160 307255
rect 131210 306776 131266 306785
rect 131210 306711 131266 306720
rect 131120 306468 131172 306474
rect 131120 306410 131172 306416
rect 131224 306406 131252 306711
rect 131212 306400 131264 306406
rect 131212 306342 131264 306348
rect 131118 306096 131174 306105
rect 131118 306031 131174 306040
rect 131132 305114 131160 306031
rect 131486 305552 131542 305561
rect 131486 305487 131542 305496
rect 131500 305182 131528 305487
rect 131488 305176 131540 305182
rect 131488 305118 131540 305124
rect 131120 305108 131172 305114
rect 131120 305050 131172 305056
rect 131212 305040 131264 305046
rect 131210 305008 131212 305017
rect 131264 305008 131266 305017
rect 131210 304943 131266 304952
rect 131302 304328 131358 304337
rect 131302 304263 131358 304272
rect 131210 303784 131266 303793
rect 131316 303754 131344 304263
rect 131210 303719 131266 303728
rect 131304 303748 131356 303754
rect 131224 303686 131252 303719
rect 131304 303690 131356 303696
rect 131212 303680 131264 303686
rect 131212 303622 131264 303628
rect 131118 303240 131174 303249
rect 131118 303175 131174 303184
rect 131132 302326 131160 303175
rect 131210 302696 131266 302705
rect 131210 302631 131266 302640
rect 131120 302320 131172 302326
rect 131120 302262 131172 302268
rect 131224 302258 131252 302631
rect 131212 302252 131264 302258
rect 131212 302194 131264 302200
rect 131486 302016 131542 302025
rect 131486 301951 131542 301960
rect 131212 300960 131264 300966
rect 131210 300928 131212 300937
rect 131264 300928 131266 300937
rect 131500 300898 131528 301951
rect 131210 300863 131266 300872
rect 131488 300892 131540 300898
rect 131488 300834 131540 300840
rect 131118 300112 131174 300121
rect 131118 300047 131174 300056
rect 131132 299946 131160 300047
rect 131120 299940 131172 299946
rect 131120 299882 131172 299888
rect 131028 197192 131080 197198
rect 131028 197134 131080 197140
rect 131776 197130 131804 497286
rect 131868 198898 131896 497354
rect 131948 419756 132000 419762
rect 131948 419698 132000 419704
rect 131960 400217 131988 419698
rect 131946 400208 132002 400217
rect 131946 400143 132002 400152
rect 131946 397896 132002 397905
rect 131946 397831 132002 397840
rect 131960 378146 131988 397831
rect 132038 393816 132094 393825
rect 132038 393751 132094 393760
rect 132052 393378 132080 393751
rect 132040 393372 132092 393378
rect 132040 393314 132092 393320
rect 132038 392728 132094 392737
rect 132038 392663 132094 392672
rect 132052 392086 132080 392663
rect 132040 392080 132092 392086
rect 132040 392022 132092 392028
rect 132222 381712 132278 381721
rect 132222 381647 132278 381656
rect 132236 381070 132264 381647
rect 132224 381064 132276 381070
rect 132224 381006 132276 381012
rect 131948 378140 132000 378146
rect 131948 378082 132000 378088
rect 131946 371240 132002 371249
rect 131946 371175 132002 371184
rect 131960 329798 131988 371175
rect 132222 366616 132278 366625
rect 132222 366551 132278 366560
rect 132236 362234 132264 366551
rect 132224 362228 132276 362234
rect 132224 362170 132276 362176
rect 132130 360768 132186 360777
rect 132130 360703 132186 360712
rect 132038 359544 132094 359553
rect 132038 359479 132094 359488
rect 132052 358902 132080 359479
rect 132040 358896 132092 358902
rect 132040 358838 132092 358844
rect 132144 354674 132172 360703
rect 132052 354646 132172 354674
rect 132052 340202 132080 354646
rect 132040 340196 132092 340202
rect 132040 340138 132092 340144
rect 132038 337512 132094 337521
rect 132038 337447 132094 337456
rect 132052 336870 132080 337447
rect 132040 336864 132092 336870
rect 132040 336806 132092 336812
rect 132222 334656 132278 334665
rect 132222 334591 132278 334600
rect 132236 334082 132264 334591
rect 132224 334076 132276 334082
rect 132224 334018 132276 334024
rect 132222 332344 132278 332353
rect 132222 332279 132278 332288
rect 132236 331362 132264 332279
rect 132224 331356 132276 331362
rect 132224 331298 132276 331304
rect 132222 330576 132278 330585
rect 132222 330511 132278 330520
rect 132236 330002 132264 330511
rect 132224 329996 132276 330002
rect 132224 329938 132276 329944
rect 131948 329792 132000 329798
rect 131948 329734 132000 329740
rect 132222 327040 132278 327049
rect 132222 326975 132278 326984
rect 132236 325854 132264 326975
rect 132224 325848 132276 325854
rect 132224 325790 132276 325796
rect 131946 320104 132002 320113
rect 131946 320039 132002 320048
rect 131960 291854 131988 320039
rect 132222 319560 132278 319569
rect 132222 319495 132278 319504
rect 132236 318918 132264 319495
rect 132224 318912 132276 318918
rect 132224 318854 132276 318860
rect 132130 318336 132186 318345
rect 132130 318271 132186 318280
rect 132038 301472 132094 301481
rect 132038 301407 132094 301416
rect 131948 291848 132000 291854
rect 131948 291790 132000 291796
rect 132052 279478 132080 301407
rect 132144 297430 132172 318271
rect 132222 317112 132278 317121
rect 132222 317047 132278 317056
rect 132236 316130 132264 317047
rect 132224 316124 132276 316130
rect 132224 316066 132276 316072
rect 132132 297424 132184 297430
rect 132132 297366 132184 297372
rect 132040 279472 132092 279478
rect 132040 279414 132092 279420
rect 131856 198892 131908 198898
rect 131856 198834 131908 198840
rect 133156 198830 133184 497422
rect 133786 496904 133842 496913
rect 133786 496839 133842 496848
rect 136546 496904 136602 496913
rect 136546 496839 136602 496848
rect 139306 496904 139362 496913
rect 139306 496839 139362 496848
rect 142066 496904 142122 496913
rect 142066 496839 142122 496848
rect 143446 496904 143502 496913
rect 143446 496839 143502 496848
rect 133800 479534 133828 496839
rect 133788 479528 133840 479534
rect 133788 479470 133840 479476
rect 136560 411262 136588 496839
rect 139320 412622 139348 496839
rect 142080 436830 142108 496839
rect 143460 438190 143488 496839
rect 143448 438184 143500 438190
rect 143448 438126 143500 438132
rect 142068 436824 142120 436830
rect 142068 436766 142120 436772
rect 146220 423094 146248 498063
rect 148966 496904 149022 496913
rect 151004 496874 151032 498063
rect 148966 496839 149022 496848
rect 150900 496868 150952 496874
rect 146208 423088 146260 423094
rect 146208 423030 146260 423036
rect 139308 412616 139360 412622
rect 139308 412558 139360 412564
rect 136548 411256 136600 411262
rect 136548 411198 136600 411204
rect 144184 398880 144236 398886
rect 144184 398822 144236 398828
rect 142804 397520 142856 397526
rect 142804 397462 142856 397468
rect 140228 396228 140280 396234
rect 140228 396170 140280 396176
rect 137468 392080 137520 392086
rect 137468 392022 137520 392028
rect 134708 390652 134760 390658
rect 134708 390594 134760 390600
rect 134524 389360 134576 389366
rect 134524 389302 134576 389308
rect 133512 387932 133564 387938
rect 133512 387874 133564 387880
rect 133420 386640 133472 386646
rect 133420 386582 133472 386588
rect 133328 382356 133380 382362
rect 133328 382298 133380 382304
rect 133236 363112 133288 363118
rect 133236 363054 133288 363060
rect 133248 315994 133276 363054
rect 133340 351898 133368 382298
rect 133432 357406 133460 386582
rect 133524 360194 133552 387874
rect 134536 364342 134564 389302
rect 134616 389292 134668 389298
rect 134616 389234 134668 389240
rect 134524 364336 134576 364342
rect 134524 364278 134576 364284
rect 134628 361554 134656 389234
rect 134720 367062 134748 390594
rect 137376 376848 137428 376854
rect 137376 376790 137428 376796
rect 137284 371340 137336 371346
rect 137284 371282 137336 371288
rect 135904 367260 135956 367266
rect 135904 367202 135956 367208
rect 134708 367056 134760 367062
rect 134708 366998 134760 367004
rect 134616 361548 134668 361554
rect 134616 361490 134668 361496
rect 134524 360324 134576 360330
rect 134524 360266 134576 360272
rect 133512 360188 133564 360194
rect 133512 360130 133564 360136
rect 133420 357400 133472 357406
rect 133420 357342 133472 357348
rect 133328 351892 133380 351898
rect 133328 351834 133380 351840
rect 133512 329996 133564 330002
rect 133512 329938 133564 329944
rect 133420 325712 133472 325718
rect 133420 325654 133472 325660
rect 133328 316124 133380 316130
rect 133328 316066 133380 316072
rect 133236 315988 133288 315994
rect 133236 315930 133288 315936
rect 133236 305040 133288 305046
rect 133236 304982 133288 304988
rect 133248 209778 133276 304982
rect 133340 231810 133368 316066
rect 133432 248402 133460 325654
rect 133524 255270 133552 329938
rect 134536 311846 134564 360266
rect 134892 348356 134944 348362
rect 134892 348298 134944 348304
rect 134800 347880 134852 347886
rect 134800 347822 134852 347828
rect 134524 311840 134576 311846
rect 134524 311782 134576 311788
rect 134708 309664 134760 309670
rect 134708 309606 134760 309612
rect 134616 307964 134668 307970
rect 134616 307906 134668 307912
rect 134524 299940 134576 299946
rect 134524 299882 134576 299888
rect 133512 255264 133564 255270
rect 133512 255206 133564 255212
rect 133420 248396 133472 248402
rect 133420 248338 133472 248344
rect 133328 231804 133380 231810
rect 133328 231746 133380 231752
rect 133236 209772 133288 209778
rect 133236 209714 133288 209720
rect 134536 201482 134564 299882
rect 134628 215286 134656 307906
rect 134720 219434 134748 309606
rect 134812 287026 134840 347822
rect 134904 289814 134932 348298
rect 135916 324290 135944 367202
rect 137296 331226 137324 371282
rect 137388 339454 137416 376790
rect 137480 368490 137508 392022
rect 138664 381064 138716 381070
rect 138664 381006 138716 381012
rect 137468 368484 137520 368490
rect 137468 368426 137520 368432
rect 138676 349110 138704 381006
rect 140240 375358 140268 396170
rect 141516 396160 141568 396166
rect 141516 396102 141568 396108
rect 141424 385212 141476 385218
rect 141424 385154 141476 385160
rect 140228 375352 140280 375358
rect 140228 375294 140280 375300
rect 140136 374196 140188 374202
rect 140136 374138 140188 374144
rect 140044 374128 140096 374134
rect 140044 374070 140096 374076
rect 138848 356244 138900 356250
rect 138848 356186 138900 356192
rect 138664 349104 138716 349110
rect 138664 349046 138716 349052
rect 137560 339584 137612 339590
rect 137560 339526 137612 339532
rect 137376 339448 137428 339454
rect 137376 339390 137428 339396
rect 137468 338224 137520 338230
rect 137468 338166 137520 338172
rect 137284 331220 137336 331226
rect 137284 331162 137336 331168
rect 135904 324284 135956 324290
rect 135904 324226 135956 324232
rect 137376 323128 137428 323134
rect 137376 323070 137428 323076
rect 137284 305108 137336 305114
rect 137284 305050 137336 305056
rect 135904 302320 135956 302326
rect 135904 302262 135956 302268
rect 134892 289808 134944 289814
rect 134892 289750 134944 289756
rect 134800 287020 134852 287026
rect 134800 286962 134852 286968
rect 134708 219428 134760 219434
rect 134708 219370 134760 219376
rect 134616 215280 134668 215286
rect 134616 215222 134668 215228
rect 135916 206990 135944 302262
rect 137296 211138 137324 305050
rect 137388 242894 137416 323070
rect 137480 270502 137508 338166
rect 137572 273222 137600 339526
rect 138756 314764 138808 314770
rect 138756 314706 138808 314712
rect 138664 300960 138716 300966
rect 138664 300902 138716 300908
rect 137560 273216 137612 273222
rect 137560 273158 137612 273164
rect 137468 270496 137520 270502
rect 137468 270438 137520 270444
rect 137376 242888 137428 242894
rect 137376 242830 137428 242836
rect 137284 211132 137336 211138
rect 137284 211074 137336 211080
rect 135904 206984 135956 206990
rect 135904 206926 135956 206932
rect 138676 202842 138704 300902
rect 138768 229090 138796 314706
rect 138860 302190 138888 356186
rect 140056 335306 140084 374070
rect 140148 336734 140176 374138
rect 141436 356046 141464 385154
rect 141528 376718 141556 396102
rect 142816 379506 142844 397462
rect 144196 380866 144224 398822
rect 147036 383784 147088 383790
rect 147036 383726 147088 383732
rect 144184 380860 144236 380866
rect 144184 380802 144236 380808
rect 142804 379500 142856 379506
rect 142804 379442 142856 379448
rect 142896 378344 142948 378350
rect 142896 378286 142948 378292
rect 141516 376712 141568 376718
rect 141516 376654 141568 376660
rect 142804 372700 142856 372706
rect 142804 372642 142856 372648
rect 141424 356040 141476 356046
rect 141424 355982 141476 355988
rect 141516 354816 141568 354822
rect 141516 354758 141568 354764
rect 140136 336728 140188 336734
rect 140136 336670 140188 336676
rect 140228 335436 140280 335442
rect 140228 335378 140280 335384
rect 140044 335300 140096 335306
rect 140044 335242 140096 335248
rect 140136 332784 140188 332790
rect 140136 332726 140188 332732
rect 140044 331356 140096 331362
rect 140044 331298 140096 331304
rect 138848 302184 138900 302190
rect 138848 302126 138900 302132
rect 140056 259418 140084 331298
rect 140148 262206 140176 332726
rect 140240 264926 140268 335378
rect 141424 309188 141476 309194
rect 141424 309130 141476 309136
rect 140228 264920 140280 264926
rect 140228 264862 140280 264868
rect 140136 262200 140188 262206
rect 140136 262142 140188 262148
rect 140044 259412 140096 259418
rect 140044 259354 140096 259360
rect 138756 229084 138808 229090
rect 138756 229026 138808 229032
rect 141436 218006 141464 309130
rect 141528 299470 141556 354758
rect 141700 352096 141752 352102
rect 141700 352038 141752 352044
rect 141608 350668 141660 350674
rect 141608 350610 141660 350616
rect 141516 299464 141568 299470
rect 141516 299406 141568 299412
rect 141516 297424 141568 297430
rect 141516 297366 141568 297372
rect 141528 233238 141556 297366
rect 141620 293962 141648 350610
rect 141712 296682 141740 352038
rect 142816 333946 142844 372642
rect 142908 343602 142936 378286
rect 146944 378276 146996 378282
rect 146944 378218 146996 378224
rect 144184 375488 144236 375494
rect 144184 375430 144236 375436
rect 143080 345228 143132 345234
rect 143080 345170 143132 345176
rect 142896 343596 142948 343602
rect 142896 343538 142948 343544
rect 142988 334076 143040 334082
rect 142988 334018 143040 334024
rect 142804 333940 142856 333946
rect 142804 333882 142856 333888
rect 142896 332716 142948 332722
rect 142896 332658 142948 332664
rect 142804 306468 142856 306474
rect 142804 306410 142856 306416
rect 141700 296676 141752 296682
rect 141700 296618 141752 296624
rect 141608 293956 141660 293962
rect 141608 293898 141660 293904
rect 141516 233232 141568 233238
rect 141516 233174 141568 233180
rect 141424 218000 141476 218006
rect 141424 217942 141476 217948
rect 142816 213926 142844 306410
rect 142908 260846 142936 332658
rect 143000 263566 143028 334018
rect 143092 284306 143120 345170
rect 144196 338094 144224 375430
rect 145748 356176 145800 356182
rect 145748 356118 145800 356124
rect 144460 352028 144512 352034
rect 144460 351970 144512 351976
rect 144368 342372 144420 342378
rect 144368 342314 144420 342320
rect 144184 338088 144236 338094
rect 144184 338030 144236 338036
rect 144276 321700 144328 321706
rect 144276 321642 144328 321648
rect 144184 303748 144236 303754
rect 144184 303690 144236 303696
rect 143080 284300 143132 284306
rect 143080 284242 143132 284248
rect 142988 263560 143040 263566
rect 142988 263502 143040 263508
rect 142896 260840 142948 260846
rect 142896 260782 142948 260788
rect 142804 213920 142856 213926
rect 142804 213862 142856 213868
rect 144196 208350 144224 303690
rect 144288 240106 144316 321642
rect 144380 278730 144408 342314
rect 144472 295322 144500 351970
rect 145656 347812 145708 347818
rect 145656 347754 145708 347760
rect 145564 307896 145616 307902
rect 145564 307838 145616 307844
rect 144460 295316 144512 295322
rect 144460 295258 144512 295264
rect 144368 278724 144420 278730
rect 144368 278666 144420 278672
rect 144276 240100 144328 240106
rect 144276 240042 144328 240048
rect 145576 216646 145604 307838
rect 145668 288386 145696 347754
rect 145760 303618 145788 356118
rect 146956 342242 146984 378218
rect 147048 353258 147076 383726
rect 148508 361684 148560 361690
rect 148508 361626 148560 361632
rect 147036 353252 147088 353258
rect 147036 353194 147088 353200
rect 148416 351960 148468 351966
rect 148416 351902 148468 351908
rect 147220 349240 147272 349246
rect 147220 349182 147272 349188
rect 146944 342236 146996 342242
rect 146944 342178 146996 342184
rect 147036 336932 147088 336938
rect 147036 336874 147088 336880
rect 145748 303612 145800 303618
rect 145748 303554 145800 303560
rect 146944 300892 146996 300898
rect 146944 300834 146996 300840
rect 145656 288380 145708 288386
rect 145656 288322 145708 288328
rect 145564 216640 145616 216646
rect 145564 216582 145616 216588
rect 144184 208344 144236 208350
rect 144184 208286 144236 208292
rect 146956 204270 146984 300834
rect 147048 267714 147076 336874
rect 147128 335368 147180 335374
rect 147128 335310 147180 335316
rect 147036 267708 147088 267714
rect 147036 267650 147088 267656
rect 147140 266354 147168 335310
rect 147232 291174 147260 349182
rect 148324 311976 148376 311982
rect 148324 311918 148376 311924
rect 147220 291168 147272 291174
rect 147220 291110 147272 291116
rect 147128 266348 147180 266354
rect 147128 266290 147180 266296
rect 148336 223582 148364 311918
rect 148428 295254 148456 351902
rect 148520 313274 148548 361626
rect 148508 313268 148560 313274
rect 148508 313210 148560 313216
rect 148416 295248 148468 295254
rect 148416 295190 148468 295196
rect 148324 223576 148376 223582
rect 148324 223518 148376 223524
rect 146944 204264 146996 204270
rect 146944 204206 146996 204212
rect 138664 202836 138716 202842
rect 138664 202778 138716 202784
rect 134524 201476 134576 201482
rect 134524 201418 134576 201424
rect 133144 198824 133196 198830
rect 133144 198766 133196 198772
rect 148980 197334 149008 496839
rect 150900 496810 150952 496816
rect 150992 496868 151044 496874
rect 150992 496810 151044 496816
rect 150912 489914 150940 496810
rect 150912 489886 151124 489914
rect 149704 341080 149756 341086
rect 149704 341022 149756 341028
rect 149716 274650 149744 341022
rect 149704 274644 149756 274650
rect 149704 274586 149756 274592
rect 148968 197328 149020 197334
rect 148968 197270 149020 197276
rect 151096 197266 151124 489886
rect 154500 450566 154528 498063
rect 157246 496904 157302 496913
rect 157246 496839 157302 496848
rect 155224 487824 155276 487830
rect 155224 487766 155276 487772
rect 154488 450560 154540 450566
rect 154488 450502 154540 450508
rect 152556 390584 152608 390590
rect 152556 390526 152608 390532
rect 151176 379636 151228 379642
rect 151176 379578 151228 379584
rect 151188 346390 151216 379578
rect 152464 368620 152516 368626
rect 152464 368562 152516 368568
rect 151176 346384 151228 346390
rect 151176 346326 151228 346332
rect 151268 336864 151320 336870
rect 151268 336806 151320 336812
rect 151176 324420 151228 324426
rect 151176 324362 151228 324368
rect 151188 245614 151216 324362
rect 151280 269074 151308 336806
rect 152476 325650 152504 368562
rect 152568 365702 152596 390526
rect 155236 386374 155264 487766
rect 157260 451926 157288 496839
rect 163504 496120 163556 496126
rect 163504 496062 163556 496068
rect 162124 489184 162176 489190
rect 162124 489126 162176 489132
rect 157248 451920 157300 451926
rect 157248 451862 157300 451868
rect 162136 396030 162164 489126
rect 162124 396024 162176 396030
rect 162124 395966 162176 395972
rect 162216 394800 162268 394806
rect 162216 394742 162268 394748
rect 160744 393440 160796 393446
rect 160744 393382 160796 393388
rect 159364 392012 159416 392018
rect 159364 391954 159416 391960
rect 157984 387864 158036 387870
rect 157984 387806 158036 387812
rect 155224 386368 155276 386374
rect 155224 386310 155276 386316
rect 155316 385144 155368 385150
rect 155316 385086 155368 385092
rect 152556 365696 152608 365702
rect 152556 365638 152608 365644
rect 152740 363044 152792 363050
rect 152740 362986 152792 362992
rect 152648 338156 152700 338162
rect 152648 338098 152700 338104
rect 152556 328568 152608 328574
rect 152556 328510 152608 328516
rect 152464 325644 152516 325650
rect 152464 325586 152516 325592
rect 152464 313404 152516 313410
rect 152464 313346 152516 313352
rect 151268 269068 151320 269074
rect 151268 269010 151320 269016
rect 151176 245608 151228 245614
rect 151176 245550 151228 245556
rect 152476 224942 152504 313346
rect 152568 253910 152596 328510
rect 152660 271862 152688 338098
rect 152752 314634 152780 362986
rect 155328 354686 155356 385086
rect 156696 385076 156748 385082
rect 156696 385018 156748 385024
rect 156604 374060 156656 374066
rect 156604 374002 156656 374008
rect 155316 354680 155368 354686
rect 155316 354622 155368 354628
rect 155500 353388 155552 353394
rect 155500 353330 155552 353336
rect 155408 345160 155460 345166
rect 155408 345102 155460 345108
rect 153844 343732 153896 343738
rect 153844 343674 153896 343680
rect 152740 314628 152792 314634
rect 152740 314570 152792 314576
rect 153856 281518 153884 343674
rect 155316 321632 155368 321638
rect 155316 321574 155368 321580
rect 155224 316056 155276 316062
rect 155224 315998 155276 316004
rect 153844 281512 153896 281518
rect 153844 281454 153896 281460
rect 152648 271856 152700 271862
rect 152648 271798 152700 271804
rect 152556 253904 152608 253910
rect 152556 253846 152608 253852
rect 155236 230450 155264 315998
rect 155328 241466 155356 321574
rect 155420 282878 155448 345102
rect 155512 298110 155540 353330
rect 156616 335238 156644 374002
rect 156708 357338 156736 385018
rect 157996 361486 158024 387806
rect 159376 369850 159404 391954
rect 160756 371210 160784 393382
rect 162228 373998 162256 394742
rect 162216 373992 162268 373998
rect 162216 373934 162268 373940
rect 160744 371204 160796 371210
rect 160744 371146 160796 371152
rect 162124 369980 162176 369986
rect 162124 369922 162176 369928
rect 159364 369844 159416 369850
rect 159364 369786 159416 369792
rect 160744 367192 160796 367198
rect 160744 367134 160796 367140
rect 159364 362976 159416 362982
rect 159364 362918 159416 362924
rect 157984 361480 158036 361486
rect 157984 361422 158036 361428
rect 158260 360256 158312 360262
rect 158260 360198 158312 360204
rect 156696 357332 156748 357338
rect 156696 357274 156748 357280
rect 158168 356108 158220 356114
rect 158168 356050 158220 356056
rect 156788 354748 156840 354754
rect 156788 354690 156840 354696
rect 156604 335232 156656 335238
rect 156604 335174 156656 335180
rect 156696 323060 156748 323066
rect 156696 323002 156748 323008
rect 156604 318912 156656 318918
rect 156604 318854 156656 318860
rect 155500 298104 155552 298110
rect 155500 298046 155552 298052
rect 155408 282872 155460 282878
rect 155408 282814 155460 282820
rect 155316 241460 155368 241466
rect 155316 241402 155368 241408
rect 156616 235958 156644 318854
rect 156708 244254 156736 323002
rect 156800 300830 156828 354690
rect 158076 325780 158128 325786
rect 158076 325722 158128 325728
rect 157984 313336 158036 313342
rect 157984 313278 158036 313284
rect 156788 300824 156840 300830
rect 156788 300766 156840 300772
rect 156696 244248 156748 244254
rect 156696 244190 156748 244196
rect 156604 235952 156656 235958
rect 156604 235894 156656 235900
rect 155224 230444 155276 230450
rect 155224 230386 155276 230392
rect 157996 226302 158024 313278
rect 158088 247042 158116 325722
rect 158180 304978 158208 356050
rect 158272 309126 158300 360198
rect 159376 317422 159404 362918
rect 159548 342304 159600 342310
rect 159548 342246 159600 342252
rect 159456 329928 159508 329934
rect 159456 329870 159508 329876
rect 159364 317416 159416 317422
rect 159364 317358 159416 317364
rect 159364 310616 159416 310622
rect 159364 310558 159416 310564
rect 158260 309120 158312 309126
rect 158260 309062 158312 309068
rect 158168 304972 158220 304978
rect 158168 304914 158220 304920
rect 158076 247036 158128 247042
rect 158076 246978 158128 246984
rect 157984 226296 158036 226302
rect 157984 226238 158036 226244
rect 152464 224936 152516 224942
rect 152464 224878 152516 224884
rect 159376 220794 159404 310558
rect 159468 256698 159496 329870
rect 159560 277370 159588 342246
rect 160756 322930 160784 367134
rect 160928 341012 160980 341018
rect 160928 340954 160980 340960
rect 160836 325848 160888 325854
rect 160836 325790 160888 325796
rect 160744 322924 160796 322930
rect 160744 322866 160796 322872
rect 160744 307828 160796 307834
rect 160744 307770 160796 307776
rect 159548 277364 159600 277370
rect 159548 277306 159600 277312
rect 159456 256692 159508 256698
rect 159456 256634 159508 256640
rect 159364 220788 159416 220794
rect 159364 220730 159416 220736
rect 160756 215218 160784 307770
rect 160848 249762 160876 325790
rect 160940 276010 160968 340954
rect 162136 327078 162164 369922
rect 162308 346520 162360 346526
rect 162308 346462 162360 346468
rect 162124 327072 162176 327078
rect 162124 327014 162176 327020
rect 162216 320272 162268 320278
rect 162216 320214 162268 320220
rect 162124 302252 162176 302258
rect 162124 302194 162176 302200
rect 160928 276004 160980 276010
rect 160928 275946 160980 275952
rect 160836 249756 160888 249762
rect 160836 249698 160888 249704
rect 160744 215212 160796 215218
rect 160744 215154 160796 215160
rect 162136 205630 162164 302194
rect 162228 238746 162256 320214
rect 162320 285666 162348 346462
rect 162308 285660 162360 285666
rect 162308 285602 162360 285608
rect 162216 238740 162268 238746
rect 162216 238682 162268 238688
rect 162124 205624 162176 205630
rect 162124 205566 162176 205572
rect 163516 198422 163544 496062
rect 175924 493332 175976 493338
rect 175924 493274 175976 493280
rect 166264 491972 166316 491978
rect 166264 491914 166316 491920
rect 164884 406428 164936 406434
rect 164884 406370 164936 406376
rect 163688 365764 163740 365770
rect 163688 365706 163740 365712
rect 163596 334008 163648 334014
rect 163596 333950 163648 333956
rect 163608 264858 163636 333950
rect 163700 320142 163728 365706
rect 163688 320136 163740 320142
rect 163688 320078 163740 320084
rect 163596 264852 163648 264858
rect 163596 264794 163648 264800
rect 163504 198416 163556 198422
rect 163504 198358 163556 198364
rect 164896 198014 164924 406370
rect 165068 389836 165120 389842
rect 165068 389778 165120 389784
rect 164976 371272 165028 371278
rect 164976 371214 165028 371220
rect 164988 331158 165016 371214
rect 165080 366994 165108 389778
rect 166276 389162 166304 491914
rect 170404 490612 170456 490618
rect 170404 490554 170456 490560
rect 169760 421116 169812 421122
rect 169760 421058 169812 421064
rect 166264 389156 166316 389162
rect 166264 389098 166316 389104
rect 166264 376780 166316 376786
rect 166264 376722 166316 376728
rect 165068 366988 165120 366994
rect 165068 366930 165120 366936
rect 165160 358896 165212 358902
rect 165160 358838 165212 358844
rect 164976 331152 165028 331158
rect 164976 331094 165028 331100
rect 165068 329860 165120 329866
rect 165068 329802 165120 329808
rect 164976 311908 165028 311914
rect 164976 311850 165028 311856
rect 164988 222154 165016 311850
rect 165080 255202 165108 329802
rect 165172 309058 165200 358838
rect 166276 340882 166304 376722
rect 169116 364472 169168 364478
rect 169116 364414 169168 364420
rect 166448 357536 166500 357542
rect 166448 357478 166500 357484
rect 166264 340876 166316 340882
rect 166264 340818 166316 340824
rect 166356 339516 166408 339522
rect 166356 339458 166408 339464
rect 166264 327208 166316 327214
rect 166264 327150 166316 327156
rect 165160 309052 165212 309058
rect 165160 308994 165212 309000
rect 165068 255196 165120 255202
rect 165068 255138 165120 255144
rect 166276 251190 166304 327150
rect 166368 273154 166396 339458
rect 166460 306338 166488 357478
rect 169024 324352 169076 324358
rect 169024 324294 169076 324300
rect 166448 306332 166500 306338
rect 166448 306274 166500 306280
rect 166356 273148 166408 273154
rect 166356 273090 166408 273096
rect 166264 251184 166316 251190
rect 166264 251126 166316 251132
rect 169036 246974 169064 324294
rect 169128 318782 169156 364414
rect 169116 318776 169168 318782
rect 169116 318718 169168 318724
rect 169024 246968 169076 246974
rect 169024 246910 169076 246916
rect 164976 222148 165028 222154
rect 164976 222090 165028 222096
rect 164884 198008 164936 198014
rect 164884 197950 164936 197956
rect 151084 197260 151136 197266
rect 151084 197202 151136 197208
rect 131764 197124 131816 197130
rect 131764 197066 131816 197072
rect 130476 197056 130528 197062
rect 130476 196998 130528 197004
rect 130384 196988 130436 196994
rect 130384 196930 130436 196936
rect 168286 195392 168342 195401
rect 168286 195327 168342 195336
rect 167366 195256 167422 195265
rect 167366 195191 167422 195200
rect 166908 139596 166960 139602
rect 166908 139538 166960 139544
rect 165528 139528 165580 139534
rect 165528 139470 165580 139476
rect 165540 96626 165568 139470
rect 166920 117881 166948 139538
rect 167380 136649 167408 195191
rect 168102 145616 168158 145625
rect 168102 145551 168158 145560
rect 167552 140276 167604 140282
rect 167552 140218 167604 140224
rect 167460 140140 167512 140146
rect 167460 140082 167512 140088
rect 167366 136640 167422 136649
rect 167366 136575 167422 136584
rect 166906 117872 166962 117881
rect 166906 117807 166962 117816
rect 165528 96620 165580 96626
rect 165528 96562 165580 96568
rect 167000 96620 167052 96626
rect 167000 96562 167052 96568
rect 167012 96529 167040 96562
rect 166998 96520 167054 96529
rect 166998 96455 167054 96464
rect 167472 80209 167500 140082
rect 167564 136134 167592 140218
rect 167828 140072 167880 140078
rect 167828 140014 167880 140020
rect 167734 139632 167790 139641
rect 167734 139567 167790 139576
rect 167644 139460 167696 139466
rect 167644 139402 167696 139408
rect 167552 136128 167604 136134
rect 167552 136070 167604 136076
rect 167552 135992 167604 135998
rect 167552 135934 167604 135940
rect 167564 134094 167592 135934
rect 167552 134088 167604 134094
rect 167552 134030 167604 134036
rect 167656 111353 167684 139402
rect 167642 111344 167698 111353
rect 167642 111279 167698 111288
rect 167748 106457 167776 139567
rect 167840 134230 167868 140014
rect 168012 139936 168064 139942
rect 168012 139878 168064 139884
rect 167920 139868 167972 139874
rect 167920 139810 167972 139816
rect 167828 134224 167880 134230
rect 167828 134166 167880 134172
rect 167828 134088 167880 134094
rect 167828 134030 167880 134036
rect 167734 106448 167790 106457
rect 167734 106383 167790 106392
rect 167840 98297 167868 134030
rect 167826 98288 167882 98297
rect 167826 98223 167882 98232
rect 167932 90001 167960 139810
rect 168024 136218 168052 139878
rect 168116 139505 168144 145551
rect 168196 141092 168248 141098
rect 168196 141034 168248 141040
rect 168102 139496 168158 139505
rect 168102 139431 168158 139440
rect 168024 136190 168144 136218
rect 168012 136128 168064 136134
rect 168012 136070 168064 136076
rect 167918 89992 167974 90001
rect 167918 89927 167974 89936
rect 168024 88369 168052 136070
rect 168010 88360 168066 88369
rect 168010 88295 168066 88304
rect 168116 83473 168144 136190
rect 168208 134337 168236 141034
rect 168300 139913 168328 195327
rect 168932 151088 168984 151094
rect 168932 151030 168984 151036
rect 168840 148368 168892 148374
rect 168840 148310 168892 148316
rect 168380 140208 168432 140214
rect 168380 140150 168432 140156
rect 168286 139904 168342 139913
rect 168286 139839 168342 139848
rect 168288 139664 168340 139670
rect 168288 139606 168340 139612
rect 168194 134328 168250 134337
rect 168194 134263 168250 134272
rect 168196 134224 168248 134230
rect 168196 134166 168248 134172
rect 168208 86737 168236 134166
rect 168300 114617 168328 139606
rect 168392 135998 168420 140150
rect 168380 135992 168432 135998
rect 168380 135934 168432 135940
rect 168852 126177 168880 148310
rect 168838 126168 168894 126177
rect 168838 126103 168894 126112
rect 168944 124545 168972 151030
rect 169208 145580 169260 145586
rect 169208 145522 169260 145528
rect 169116 139732 169168 139738
rect 169116 139674 169168 139680
rect 168930 124536 168986 124545
rect 168930 124471 168986 124480
rect 169128 116249 169156 139674
rect 169220 119649 169248 145522
rect 169668 140956 169720 140962
rect 169668 140898 169720 140904
rect 169576 140888 169628 140894
rect 169576 140830 169628 140836
rect 169300 140004 169352 140010
rect 169300 139946 169352 139952
rect 169206 119640 169262 119649
rect 169206 119575 169262 119584
rect 169114 116240 169170 116249
rect 169114 116175 169170 116184
rect 168286 114608 168342 114617
rect 168286 114543 168342 114552
rect 169312 112985 169340 139946
rect 169392 139800 169444 139806
rect 169392 139742 169444 139748
rect 169298 112976 169354 112985
rect 169298 112911 169354 112920
rect 169404 109721 169432 139742
rect 169482 139632 169538 139641
rect 169482 139567 169538 139576
rect 169390 109712 169446 109721
rect 169390 109647 169446 109656
rect 169496 108089 169524 139567
rect 169482 108080 169538 108089
rect 169482 108015 169538 108024
rect 169588 101561 169616 140830
rect 169574 101552 169630 101561
rect 169574 101487 169630 101496
rect 169680 99929 169708 140898
rect 169772 131073 169800 421058
rect 170416 389094 170444 490554
rect 173164 414044 173216 414050
rect 173164 413986 173216 413992
rect 171048 409896 171100 409902
rect 171048 409838 171100 409844
rect 170404 389088 170456 389094
rect 170404 389030 170456 389036
rect 170404 372632 170456 372638
rect 170404 372574 170456 372580
rect 170416 332586 170444 372574
rect 170588 345092 170640 345098
rect 170588 345034 170640 345040
rect 170404 332580 170456 332586
rect 170404 332522 170456 332528
rect 170496 331288 170548 331294
rect 170496 331230 170548 331236
rect 170404 313948 170456 313954
rect 170404 313890 170456 313896
rect 170416 227730 170444 313890
rect 170508 258058 170536 331230
rect 170600 282810 170628 345034
rect 170588 282804 170640 282810
rect 170588 282746 170640 282752
rect 170496 258052 170548 258058
rect 170496 257994 170548 258000
rect 170404 227724 170456 227730
rect 170404 227666 170456 227672
rect 169852 188352 169904 188358
rect 169852 188294 169904 188300
rect 169864 139233 169892 188294
rect 170220 152516 170272 152522
rect 170220 152458 170272 152464
rect 170128 141024 170180 141030
rect 170128 140966 170180 140972
rect 170036 140820 170088 140826
rect 170036 140762 170088 140768
rect 169944 140344 169996 140350
rect 169944 140286 169996 140292
rect 169850 139224 169906 139233
rect 169850 139159 169906 139168
rect 169758 131064 169814 131073
rect 169758 130999 169814 131008
rect 169666 99920 169722 99929
rect 169666 99855 169722 99864
rect 169956 95169 169984 140286
rect 170048 103329 170076 140762
rect 170140 104961 170168 140966
rect 170232 133249 170260 152458
rect 170310 139768 170366 139777
rect 170310 139703 170366 139712
rect 170324 135697 170352 139703
rect 170310 135688 170366 135697
rect 170310 135623 170366 135632
rect 170218 133240 170274 133249
rect 170218 133175 170274 133184
rect 170126 104952 170182 104961
rect 170126 104887 170182 104896
rect 170034 103320 170090 103329
rect 170034 103255 170090 103264
rect 169942 95160 169998 95169
rect 169942 95095 169998 95104
rect 168194 86728 168250 86737
rect 168194 86663 168250 86672
rect 168102 83464 168158 83473
rect 168102 83399 168158 83408
rect 168102 81832 168158 81841
rect 168102 81767 168158 81776
rect 167458 80200 167514 80209
rect 167458 80135 167514 80144
rect 168010 75304 168066 75313
rect 168010 75239 168066 75248
rect 167274 73536 167330 73545
rect 167274 73471 167330 73480
rect 165528 65000 165580 65006
rect 165528 64942 165580 64948
rect 165540 31754 165568 64942
rect 167182 44024 167238 44033
rect 167182 43959 167238 43968
rect 165528 31748 165580 31754
rect 165528 31690 165580 31696
rect 167196 29986 167224 43959
rect 167184 29980 167236 29986
rect 167184 29922 167236 29928
rect 78678 28928 78734 28937
rect 167288 28898 167316 73471
rect 167642 71904 167698 71913
rect 167642 71839 167698 71848
rect 167656 70394 167684 71839
rect 167656 70366 167868 70394
rect 167734 68640 167790 68649
rect 167734 68575 167790 68584
rect 167366 53952 167422 53961
rect 167366 53887 167422 53896
rect 78678 28863 78734 28872
rect 167276 28892 167328 28898
rect 167276 28834 167328 28840
rect 28908 28348 28960 28354
rect 28908 28290 28960 28296
rect 167380 28218 167408 53887
rect 167550 48920 167606 48929
rect 167550 48855 167606 48864
rect 167458 47288 167514 47297
rect 167458 47223 167514 47232
rect 167368 28212 167420 28218
rect 167368 28154 167420 28160
rect 167472 28150 167500 47223
rect 167564 29646 167592 48855
rect 167748 41750 167776 68575
rect 167840 42090 167868 70366
rect 167918 70272 167974 70281
rect 167918 70207 167974 70216
rect 167828 42084 167880 42090
rect 167828 42026 167880 42032
rect 167826 41848 167882 41857
rect 167826 41783 167882 41792
rect 167736 41744 167788 41750
rect 167736 41686 167788 41692
rect 167840 29850 167868 41783
rect 167932 37262 167960 70207
rect 168024 40050 168052 75239
rect 168116 44198 168144 81767
rect 168194 76936 168250 76945
rect 168194 76871 168250 76880
rect 168104 44192 168156 44198
rect 168104 44134 168156 44140
rect 168208 40746 168236 76871
rect 169758 67008 169814 67017
rect 169758 66943 169814 66952
rect 168286 65376 168342 65385
rect 168286 65311 168342 65320
rect 168300 65006 168328 65311
rect 168288 65000 168340 65006
rect 168288 64942 168340 64948
rect 169666 62112 169722 62121
rect 169666 62047 169722 62056
rect 169482 58848 169538 58857
rect 169482 58783 169538 58792
rect 169390 52184 169446 52193
rect 169390 52119 169446 52128
rect 169024 44192 169076 44198
rect 169024 44134 169076 44140
rect 168286 41440 168342 41449
rect 168286 41375 168342 41384
rect 168116 40718 168236 40746
rect 168012 40044 168064 40050
rect 168012 39986 168064 39992
rect 168010 39128 168066 39137
rect 168010 39063 168066 39072
rect 167920 37256 167972 37262
rect 167920 37198 167972 37204
rect 168024 30054 168052 39063
rect 168116 33318 168144 40718
rect 168300 39953 168328 41375
rect 168286 39944 168342 39953
rect 168286 39879 168342 39888
rect 168286 37496 168342 37505
rect 168286 37431 168342 37440
rect 168300 35894 168328 37431
rect 168932 37256 168984 37262
rect 168932 37198 168984 37204
rect 168944 35894 168972 37198
rect 168208 35866 168328 35894
rect 168852 35866 168972 35894
rect 168104 33312 168156 33318
rect 168104 33254 168156 33260
rect 168012 30048 168064 30054
rect 168012 29990 168064 29996
rect 168208 29918 168236 35866
rect 168286 35320 168342 35329
rect 168286 35255 168342 35264
rect 168196 29912 168248 29918
rect 168196 29854 168248 29860
rect 167828 29844 167880 29850
rect 167828 29786 167880 29792
rect 168300 29714 168328 35255
rect 168288 29708 168340 29714
rect 168288 29650 168340 29656
rect 167552 29640 167604 29646
rect 167552 29582 167604 29588
rect 168852 28762 168880 35866
rect 168932 33516 168984 33522
rect 168932 33458 168984 33464
rect 168840 28756 168892 28762
rect 168840 28698 168892 28704
rect 167460 28144 167512 28150
rect 167460 28086 167512 28092
rect 168944 27946 168972 33458
rect 169036 30122 169064 44134
rect 169208 42084 169260 42090
rect 169208 42026 169260 42032
rect 169116 41744 169168 41750
rect 169116 41686 169168 41692
rect 169024 30116 169076 30122
rect 169024 30058 169076 30064
rect 169128 28966 169156 41686
rect 169116 28960 169168 28966
rect 169116 28902 169168 28908
rect 169220 28490 169248 42026
rect 169300 40044 169352 40050
rect 169300 39986 169352 39992
rect 169312 28558 169340 39986
rect 169404 31686 169432 52119
rect 169392 31680 169444 31686
rect 169392 31622 169444 31628
rect 169496 31618 169524 58783
rect 169574 55584 169630 55593
rect 169574 55519 169630 55528
rect 169588 33522 169616 55519
rect 169576 33516 169628 33522
rect 169576 33458 169628 33464
rect 169680 33402 169708 62047
rect 169588 33374 169708 33402
rect 169484 31612 169536 31618
rect 169484 31554 169536 31560
rect 169588 28830 169616 33374
rect 169668 33312 169720 33318
rect 169668 33254 169720 33260
rect 169680 30326 169708 33254
rect 169668 30320 169720 30326
rect 169668 30262 169720 30268
rect 169576 28824 169628 28830
rect 169576 28766 169628 28772
rect 169300 28552 169352 28558
rect 169300 28494 169352 28500
rect 169208 28484 169260 28490
rect 169208 28426 169260 28432
rect 169772 28422 169800 66943
rect 169850 50552 169906 50561
rect 169850 50487 169906 50496
rect 169864 30190 169892 50487
rect 169942 45792 169998 45801
rect 169942 45727 169998 45736
rect 169956 30258 169984 45727
rect 170586 33688 170642 33697
rect 170586 33623 170642 33632
rect 170494 32056 170550 32065
rect 170494 31991 170550 32000
rect 170402 31104 170458 31113
rect 170402 31039 170458 31048
rect 169944 30252 169996 30258
rect 169944 30194 169996 30200
rect 169852 30184 169904 30190
rect 169852 30126 169904 30132
rect 170416 29782 170444 31039
rect 170404 29776 170456 29782
rect 170508 29753 170536 31991
rect 170600 30297 170628 33623
rect 170586 30288 170642 30297
rect 170586 30223 170642 30232
rect 170404 29718 170456 29724
rect 170494 29744 170550 29753
rect 170494 29679 170550 29688
rect 169760 28416 169812 28422
rect 169760 28358 169812 28364
rect 171060 28082 171088 409838
rect 173176 141098 173204 413986
rect 174544 394732 174596 394738
rect 174544 394674 174596 394680
rect 173348 379568 173400 379574
rect 173348 379510 173400 379516
rect 173256 362228 173308 362234
rect 173256 362170 173308 362176
rect 173268 321570 173296 362170
rect 173360 345030 173388 379510
rect 174556 372570 174584 394674
rect 174544 372564 174596 372570
rect 174544 372506 174596 372512
rect 174544 368552 174596 368558
rect 174544 368494 174596 368500
rect 173348 345024 173400 345030
rect 173348 344966 173400 344972
rect 173440 343664 173492 343670
rect 173440 343606 173492 343612
rect 173256 321564 173308 321570
rect 173256 321506 173308 321512
rect 173256 318844 173308 318850
rect 173256 318786 173308 318792
rect 173268 234598 173296 318786
rect 173452 280158 173480 343606
rect 174556 327010 174584 368494
rect 174728 349172 174780 349178
rect 174728 349114 174780 349120
rect 174636 328500 174688 328506
rect 174636 328442 174688 328448
rect 174544 327004 174596 327010
rect 174544 326946 174596 326952
rect 174544 317484 174596 317490
rect 174544 317426 174596 317432
rect 173440 280152 173492 280158
rect 173440 280094 173492 280100
rect 173348 279472 173400 279478
rect 173348 279414 173400 279420
rect 173256 234592 173308 234598
rect 173256 234534 173308 234540
rect 173360 202774 173388 279414
rect 174556 233170 174584 317426
rect 174648 252550 174676 328442
rect 174740 291106 174768 349114
rect 174728 291100 174780 291106
rect 174728 291042 174780 291048
rect 174636 252544 174688 252550
rect 174636 252486 174688 252492
rect 174544 233164 174596 233170
rect 174544 233106 174596 233112
rect 173348 202768 173400 202774
rect 173348 202710 173400 202716
rect 175936 198218 175964 493274
rect 176016 486532 176068 486538
rect 176016 486474 176068 486480
rect 176028 391950 176056 486474
rect 176016 391944 176068 391950
rect 176016 391886 176068 391892
rect 176200 382288 176252 382294
rect 176200 382230 176252 382236
rect 176016 367124 176068 367130
rect 176016 367066 176068 367072
rect 176028 322862 176056 367066
rect 176108 350600 176160 350606
rect 176108 350542 176160 350548
rect 176016 322856 176068 322862
rect 176016 322798 176068 322804
rect 176016 320204 176068 320210
rect 176016 320146 176068 320152
rect 176028 237386 176056 320146
rect 176120 292534 176148 350542
rect 176212 350538 176240 382230
rect 176200 350532 176252 350538
rect 176200 350474 176252 350480
rect 176108 292528 176160 292534
rect 176108 292470 176160 292476
rect 176200 291848 176252 291854
rect 176200 291790 176252 291796
rect 176016 237380 176068 237386
rect 176016 237322 176068 237328
rect 176212 237318 176240 291790
rect 176200 237312 176252 237318
rect 176200 237254 176252 237260
rect 177316 198286 177344 498850
rect 189816 497140 189868 497146
rect 189816 497082 189868 497088
rect 189724 497072 189776 497078
rect 189724 497014 189776 497020
rect 185584 497004 185636 497010
rect 185584 496946 185636 496952
rect 184204 496188 184256 496194
rect 184204 496130 184256 496136
rect 177396 493400 177448 493406
rect 177396 493342 177448 493348
rect 177408 393310 177436 493342
rect 182824 480956 182876 480962
rect 182824 480898 182876 480904
rect 181444 478168 181496 478174
rect 181444 478110 181496 478116
rect 178684 416084 178736 416090
rect 178684 416026 178736 416032
rect 177396 393304 177448 393310
rect 177396 393246 177448 393252
rect 177488 389224 177540 389230
rect 177488 389166 177540 389172
rect 177396 369912 177448 369918
rect 177396 369854 177448 369860
rect 177408 328438 177436 369854
rect 177500 362914 177528 389166
rect 177488 362908 177540 362914
rect 177488 362850 177540 362856
rect 177580 358828 177632 358834
rect 177580 358770 177632 358776
rect 177396 328432 177448 328438
rect 177396 328374 177448 328380
rect 177488 322992 177540 322998
rect 177488 322934 177540 322940
rect 177396 306400 177448 306406
rect 177396 306342 177448 306348
rect 177408 212498 177436 306342
rect 177500 241398 177528 322934
rect 177592 307766 177620 358770
rect 177580 307760 177632 307766
rect 177580 307702 177632 307708
rect 177488 241392 177540 241398
rect 177488 241334 177540 241340
rect 177396 212492 177448 212498
rect 177396 212434 177448 212440
rect 177304 198280 177356 198286
rect 177304 198222 177356 198228
rect 175924 198212 175976 198218
rect 175924 198154 175976 198160
rect 178696 198082 178724 416026
rect 180064 413296 180116 413302
rect 180064 413238 180116 413244
rect 178868 378208 178920 378214
rect 178868 378150 178920 378156
rect 178776 361616 178828 361622
rect 178776 361558 178828 361564
rect 178788 313206 178816 361558
rect 178880 343534 178908 378150
rect 178868 343528 178920 343534
rect 178868 343470 178920 343476
rect 178868 340944 178920 340950
rect 178868 340886 178920 340892
rect 178776 313200 178828 313206
rect 178776 313142 178828 313148
rect 178776 305176 178828 305182
rect 178776 305118 178828 305124
rect 178788 211070 178816 305118
rect 178880 277302 178908 340886
rect 178868 277296 178920 277302
rect 178868 277238 178920 277244
rect 178776 211064 178828 211070
rect 178776 211006 178828 211012
rect 180076 198529 180104 413238
rect 180156 380996 180208 381002
rect 180156 380938 180208 380944
rect 180168 347750 180196 380938
rect 180156 347744 180208 347750
rect 180156 347686 180208 347692
rect 180248 346452 180300 346458
rect 180248 346394 180300 346400
rect 180156 314696 180208 314702
rect 180156 314638 180208 314644
rect 180168 229022 180196 314638
rect 180260 286958 180288 346394
rect 180340 340196 180392 340202
rect 180340 340138 180392 340144
rect 180352 310486 180380 340138
rect 180340 310480 180392 310486
rect 180340 310422 180392 310428
rect 180248 286952 180300 286958
rect 180248 286894 180300 286900
rect 180156 229016 180208 229022
rect 180156 228958 180208 228964
rect 181456 198665 181484 478110
rect 181536 393372 181588 393378
rect 181536 393314 181588 393320
rect 181548 371142 181576 393314
rect 181628 375420 181680 375426
rect 181628 375362 181680 375368
rect 181536 371136 181588 371142
rect 181536 371078 181588 371084
rect 181536 364404 181588 364410
rect 181536 364346 181588 364352
rect 181548 317354 181576 364346
rect 181640 339386 181668 375362
rect 181628 339380 181680 339386
rect 181628 339322 181680 339328
rect 181628 336796 181680 336802
rect 181628 336738 181680 336744
rect 181536 317348 181588 317354
rect 181536 317290 181588 317296
rect 181536 303680 181588 303686
rect 181536 303622 181588 303628
rect 181548 206922 181576 303622
rect 181640 269006 181668 336738
rect 181628 269000 181680 269006
rect 181628 268942 181680 268948
rect 181536 206916 181588 206922
rect 181536 206858 181588 206864
rect 182836 198694 182864 480898
rect 183008 396092 183060 396098
rect 183008 396034 183060 396040
rect 182916 383716 182968 383722
rect 182916 383658 182968 383664
rect 182928 353190 182956 383658
rect 183020 375290 183048 396034
rect 183008 375284 183060 375290
rect 183008 375226 183060 375232
rect 183100 357468 183152 357474
rect 183100 357410 183152 357416
rect 182916 353184 182968 353190
rect 182916 353126 182968 353132
rect 183008 332648 183060 332654
rect 183008 332590 183060 332596
rect 182916 310548 182968 310554
rect 182916 310490 182968 310496
rect 182928 220726 182956 310490
rect 183020 259350 183048 332590
rect 183112 304910 183140 357410
rect 183100 304904 183152 304910
rect 183100 304846 183152 304852
rect 183008 259344 183060 259350
rect 183008 259286 183060 259292
rect 182916 220720 182968 220726
rect 182916 220662 182968 220668
rect 182824 198688 182876 198694
rect 181442 198656 181498 198665
rect 182824 198630 182876 198636
rect 184216 198626 184244 496130
rect 184296 400920 184348 400926
rect 184296 400862 184348 400868
rect 181442 198591 181498 198600
rect 184204 198620 184256 198626
rect 184204 198562 184256 198568
rect 180062 198520 180118 198529
rect 180062 198455 180118 198464
rect 184308 198354 184336 400862
rect 184480 386436 184532 386442
rect 184480 386378 184532 386384
rect 184388 380928 184440 380934
rect 184388 380870 184440 380876
rect 184400 349042 184428 380870
rect 184492 358766 184520 386378
rect 184480 358760 184532 358766
rect 184480 358702 184532 358708
rect 184572 353320 184624 353326
rect 184572 353262 184624 353268
rect 184388 349036 184440 349042
rect 184388 348978 184440 348984
rect 184480 327140 184532 327146
rect 184480 327082 184532 327088
rect 184388 309800 184440 309806
rect 184388 309742 184440 309748
rect 184400 224874 184428 309742
rect 184492 251122 184520 327082
rect 184584 299402 184612 353262
rect 184572 299396 184624 299402
rect 184572 299338 184624 299344
rect 184480 251116 184532 251122
rect 184480 251058 184532 251064
rect 184388 224868 184440 224874
rect 184388 224810 184440 224816
rect 185596 198966 185624 496946
rect 188344 496936 188396 496942
rect 188344 496878 188396 496884
rect 185676 424380 185728 424386
rect 185676 424322 185728 424328
rect 185584 198960 185636 198966
rect 185584 198902 185636 198908
rect 184296 198348 184348 198354
rect 184296 198290 184348 198296
rect 185688 198150 185716 424322
rect 186228 422408 186280 422414
rect 186228 422350 186280 422356
rect 185676 198144 185728 198150
rect 185676 198086 185728 198092
rect 178684 198076 178736 198082
rect 178684 198018 178736 198024
rect 186240 197810 186268 422350
rect 186964 421524 187016 421530
rect 186964 421466 187016 421472
rect 186320 419484 186372 419490
rect 186320 419426 186372 419432
rect 186332 418441 186360 419426
rect 186318 418432 186374 418441
rect 186318 418367 186374 418376
rect 186318 415304 186374 415313
rect 186318 415239 186374 415248
rect 186332 414050 186360 415239
rect 186320 414044 186372 414050
rect 186320 413986 186372 413992
rect 186976 413846 187004 421466
rect 187516 420300 187568 420306
rect 187516 420242 187568 420248
rect 187056 420164 187108 420170
rect 187056 420106 187108 420112
rect 186964 413840 187016 413846
rect 186964 413782 187016 413788
rect 186870 413128 186926 413137
rect 186870 413063 186926 413072
rect 186320 412616 186372 412622
rect 186320 412558 186372 412564
rect 186332 412185 186360 412558
rect 186318 412176 186374 412185
rect 186318 412111 186374 412120
rect 186412 411256 186464 411262
rect 186412 411198 186464 411204
rect 186318 411088 186374 411097
rect 186318 411023 186374 411032
rect 186332 409902 186360 411023
rect 186424 410009 186452 411198
rect 186410 410000 186466 410009
rect 186410 409935 186466 409944
rect 186320 409896 186372 409902
rect 186320 409838 186372 409844
rect 186320 407108 186372 407114
rect 186320 407050 186372 407056
rect 186332 406881 186360 407050
rect 186318 406872 186374 406881
rect 186318 406807 186374 406816
rect 186320 404320 186372 404326
rect 186320 404262 186372 404268
rect 186332 403753 186360 404262
rect 186318 403744 186374 403753
rect 186318 403679 186374 403688
rect 186320 401600 186372 401606
rect 186318 401568 186320 401577
rect 186372 401568 186374 401577
rect 186318 401503 186374 401512
rect 186320 396024 186372 396030
rect 186320 395966 186372 395972
rect 186332 395321 186360 395966
rect 186318 395312 186374 395321
rect 186318 395247 186374 395256
rect 186320 393304 186372 393310
rect 186320 393246 186372 393252
rect 186332 393145 186360 393246
rect 186318 393136 186374 393145
rect 186318 393071 186374 393080
rect 186320 391944 186372 391950
rect 186320 391886 186372 391892
rect 186332 391105 186360 391886
rect 186318 391096 186374 391105
rect 186318 391031 186374 391040
rect 186412 389156 186464 389162
rect 186412 389098 186464 389104
rect 186320 389088 186372 389094
rect 186320 389030 186372 389036
rect 186332 388929 186360 389030
rect 186318 388920 186374 388929
rect 186318 388855 186374 388864
rect 186424 387977 186452 389098
rect 186410 387968 186466 387977
rect 186410 387903 186466 387912
rect 186320 386368 186372 386374
rect 186320 386310 186372 386316
rect 186332 385801 186360 386310
rect 186318 385792 186374 385801
rect 186318 385727 186374 385736
rect 186412 380860 186464 380866
rect 186412 380802 186464 380808
rect 186424 379545 186452 380802
rect 186410 379536 186466 379545
rect 186320 379500 186372 379506
rect 186410 379471 186466 379480
rect 186320 379442 186372 379448
rect 186332 378457 186360 379442
rect 186318 378448 186374 378457
rect 186318 378383 186374 378392
rect 186320 378140 186372 378146
rect 186320 378082 186372 378088
rect 186332 377369 186360 378082
rect 186318 377360 186374 377369
rect 186318 377295 186374 377304
rect 186320 376712 186372 376718
rect 186320 376654 186372 376660
rect 186332 376281 186360 376654
rect 186318 376272 186374 376281
rect 186318 376207 186374 376216
rect 186320 375352 186372 375358
rect 186320 375294 186372 375300
rect 186410 375320 186466 375329
rect 186332 374241 186360 375294
rect 186410 375255 186412 375264
rect 186464 375255 186466 375264
rect 186412 375226 186464 375232
rect 186318 374232 186374 374241
rect 186318 374167 186374 374176
rect 186320 373992 186372 373998
rect 186320 373934 186372 373940
rect 186332 373153 186360 373934
rect 186318 373144 186374 373153
rect 186318 373079 186374 373088
rect 186320 372564 186372 372570
rect 186320 372506 186372 372512
rect 186332 372065 186360 372506
rect 186318 372056 186374 372065
rect 186318 371991 186374 372000
rect 186320 371204 186372 371210
rect 186320 371146 186372 371152
rect 186332 371113 186360 371146
rect 186412 371136 186464 371142
rect 186318 371104 186374 371113
rect 186412 371078 186464 371084
rect 186318 371039 186374 371048
rect 186424 370025 186452 371078
rect 186410 370016 186466 370025
rect 186410 369951 186466 369960
rect 186320 369844 186372 369850
rect 186320 369786 186372 369792
rect 186332 368937 186360 369786
rect 186318 368928 186374 368937
rect 186318 368863 186374 368872
rect 186320 368484 186372 368490
rect 186320 368426 186372 368432
rect 186332 367849 186360 368426
rect 186318 367840 186374 367849
rect 186318 367775 186374 367784
rect 186412 367056 186464 367062
rect 186412 366998 186464 367004
rect 186320 366988 186372 366994
rect 186320 366930 186372 366936
rect 186332 366897 186360 366930
rect 186318 366888 186374 366897
rect 186318 366823 186374 366832
rect 186424 365809 186452 366998
rect 186410 365800 186466 365809
rect 186410 365735 186466 365744
rect 186320 365696 186372 365702
rect 186320 365638 186372 365644
rect 186332 364721 186360 365638
rect 186318 364712 186374 364721
rect 186318 364647 186374 364656
rect 186320 364336 186372 364342
rect 186320 364278 186372 364284
rect 186332 363633 186360 364278
rect 186318 363624 186374 363633
rect 186318 363559 186374 363568
rect 186320 362908 186372 362914
rect 186320 362850 186372 362856
rect 186332 362681 186360 362850
rect 186318 362672 186374 362681
rect 186318 362607 186374 362616
rect 186318 361584 186374 361593
rect 186318 361519 186320 361528
rect 186372 361519 186374 361528
rect 186320 361490 186372 361496
rect 186412 361480 186464 361486
rect 186412 361422 186464 361428
rect 186424 360505 186452 361422
rect 186410 360496 186466 360505
rect 186410 360431 186466 360440
rect 186320 360188 186372 360194
rect 186320 360130 186372 360136
rect 186332 359417 186360 360130
rect 186318 359408 186374 359417
rect 186318 359343 186374 359352
rect 186320 357400 186372 357406
rect 186318 357368 186320 357377
rect 186372 357368 186374 357377
rect 186318 357303 186374 357312
rect 186412 357332 186464 357338
rect 186412 357274 186464 357280
rect 186424 356289 186452 357274
rect 186410 356280 186466 356289
rect 186410 356215 186466 356224
rect 186320 356040 186372 356046
rect 186320 355982 186372 355988
rect 186332 355337 186360 355982
rect 186318 355328 186374 355337
rect 186318 355263 186374 355272
rect 186320 354680 186372 354686
rect 186320 354622 186372 354628
rect 186332 354249 186360 354622
rect 186318 354240 186374 354249
rect 186318 354175 186374 354184
rect 186320 353252 186372 353258
rect 186320 353194 186372 353200
rect 186332 352073 186360 353194
rect 186412 353184 186464 353190
rect 186410 353152 186412 353161
rect 186464 353152 186466 353161
rect 186410 353087 186466 353096
rect 186318 352064 186374 352073
rect 186318 351999 186374 352008
rect 186320 351892 186372 351898
rect 186320 351834 186372 351840
rect 186332 351121 186360 351834
rect 186318 351112 186374 351121
rect 186318 351047 186374 351056
rect 186320 350532 186372 350538
rect 186320 350474 186372 350480
rect 186332 350033 186360 350474
rect 186318 350024 186374 350033
rect 186318 349959 186374 349968
rect 186320 349104 186372 349110
rect 186320 349046 186372 349052
rect 186332 347857 186360 349046
rect 186412 349036 186464 349042
rect 186412 348978 186464 348984
rect 186424 348945 186452 348978
rect 186410 348936 186466 348945
rect 186410 348871 186466 348880
rect 186318 347848 186374 347857
rect 186318 347783 186374 347792
rect 186320 347744 186372 347750
rect 186320 347686 186372 347692
rect 186332 346905 186360 347686
rect 186318 346896 186374 346905
rect 186318 346831 186374 346840
rect 186320 346384 186372 346390
rect 186320 346326 186372 346332
rect 186332 345817 186360 346326
rect 186318 345808 186374 345817
rect 186318 345743 186374 345752
rect 186320 345024 186372 345030
rect 186320 344966 186372 344972
rect 186332 344729 186360 344966
rect 186318 344720 186374 344729
rect 186318 344655 186374 344664
rect 186318 343632 186374 343641
rect 186318 343567 186320 343576
rect 186372 343567 186374 343576
rect 186320 343538 186372 343544
rect 186412 343528 186464 343534
rect 186412 343470 186464 343476
rect 186424 342689 186452 343470
rect 186410 342680 186466 342689
rect 186410 342615 186466 342624
rect 186320 342236 186372 342242
rect 186320 342178 186372 342184
rect 186332 341601 186360 342178
rect 186318 341592 186374 341601
rect 186318 341527 186374 341536
rect 186320 340876 186372 340882
rect 186320 340818 186372 340824
rect 186332 340513 186360 340818
rect 186318 340504 186374 340513
rect 186318 340439 186374 340448
rect 186320 339448 186372 339454
rect 186318 339416 186320 339425
rect 186372 339416 186374 339425
rect 186318 339351 186374 339360
rect 186412 339380 186464 339386
rect 186412 339322 186464 339328
rect 186424 338473 186452 339322
rect 186410 338464 186466 338473
rect 186410 338399 186466 338408
rect 186320 338088 186372 338094
rect 186320 338030 186372 338036
rect 186332 337385 186360 338030
rect 186318 337376 186374 337385
rect 186318 337311 186374 337320
rect 186320 336728 186372 336734
rect 186320 336670 186372 336676
rect 186332 336297 186360 336670
rect 186318 336288 186374 336297
rect 186318 336223 186374 336232
rect 186320 335300 186372 335306
rect 186320 335242 186372 335248
rect 186332 335209 186360 335242
rect 186412 335232 186464 335238
rect 186318 335200 186374 335209
rect 186412 335174 186464 335180
rect 186318 335135 186374 335144
rect 186424 334257 186452 335174
rect 186410 334248 186466 334257
rect 186410 334183 186466 334192
rect 186320 333940 186372 333946
rect 186320 333882 186372 333888
rect 186332 333169 186360 333882
rect 186318 333160 186374 333169
rect 186318 333095 186374 333104
rect 186320 332580 186372 332586
rect 186320 332522 186372 332528
rect 186332 332081 186360 332522
rect 186318 332072 186374 332081
rect 186318 332007 186374 332016
rect 186412 331220 186464 331226
rect 186412 331162 186464 331168
rect 186320 331152 186372 331158
rect 186320 331094 186372 331100
rect 186332 330993 186360 331094
rect 186318 330984 186374 330993
rect 186318 330919 186374 330928
rect 186424 330041 186452 331162
rect 186410 330032 186466 330041
rect 186410 329967 186466 329976
rect 186320 329792 186372 329798
rect 186320 329734 186372 329740
rect 186332 328953 186360 329734
rect 186318 328944 186374 328953
rect 186318 328879 186374 328888
rect 186320 328432 186372 328438
rect 186320 328374 186372 328380
rect 186332 327865 186360 328374
rect 186318 327856 186374 327865
rect 186318 327791 186374 327800
rect 186320 327072 186372 327078
rect 186320 327014 186372 327020
rect 186332 326777 186360 327014
rect 186412 327004 186464 327010
rect 186412 326946 186464 326952
rect 186318 326768 186374 326777
rect 186318 326703 186374 326712
rect 186424 325825 186452 326946
rect 186410 325816 186466 325825
rect 186410 325751 186466 325760
rect 186320 325644 186372 325650
rect 186320 325586 186372 325592
rect 186332 324737 186360 325586
rect 186318 324728 186374 324737
rect 186318 324663 186374 324672
rect 186320 324284 186372 324290
rect 186320 324226 186372 324232
rect 186332 323649 186360 324226
rect 186318 323640 186374 323649
rect 186318 323575 186374 323584
rect 186320 322924 186372 322930
rect 186320 322866 186372 322872
rect 186332 322697 186360 322866
rect 186412 322856 186464 322862
rect 186412 322798 186464 322804
rect 186318 322688 186374 322697
rect 186318 322623 186374 322632
rect 186424 321609 186452 322798
rect 186410 321600 186466 321609
rect 186320 321564 186372 321570
rect 186410 321535 186466 321544
rect 186320 321506 186372 321512
rect 186332 320521 186360 321506
rect 186318 320512 186374 320521
rect 186318 320447 186374 320456
rect 186320 320136 186372 320142
rect 186320 320078 186372 320084
rect 186332 319433 186360 320078
rect 186318 319424 186374 319433
rect 186318 319359 186374 319368
rect 186320 318776 186372 318782
rect 186320 318718 186372 318724
rect 186332 318481 186360 318718
rect 186318 318472 186374 318481
rect 186318 318407 186374 318416
rect 186320 317416 186372 317422
rect 186320 317358 186372 317364
rect 186410 317384 186466 317393
rect 186332 316305 186360 317358
rect 186410 317319 186412 317328
rect 186464 317319 186466 317328
rect 186412 317290 186464 317296
rect 186318 316296 186374 316305
rect 186318 316231 186374 316240
rect 186320 315988 186372 315994
rect 186320 315930 186372 315936
rect 186332 315217 186360 315930
rect 186318 315208 186374 315217
rect 186318 315143 186374 315152
rect 186320 314628 186372 314634
rect 186320 314570 186372 314576
rect 186332 314265 186360 314570
rect 186318 314256 186374 314265
rect 186318 314191 186374 314200
rect 186412 313268 186464 313274
rect 186412 313210 186464 313216
rect 186320 313200 186372 313206
rect 186318 313168 186320 313177
rect 186372 313168 186374 313177
rect 186318 313103 186374 313112
rect 186424 312089 186452 313210
rect 186410 312080 186466 312089
rect 186410 312015 186466 312024
rect 186320 311840 186372 311846
rect 186320 311782 186372 311788
rect 186332 311001 186360 311782
rect 186318 310992 186374 311001
rect 186318 310927 186374 310936
rect 186320 310480 186372 310486
rect 186320 310422 186372 310428
rect 186332 310049 186360 310422
rect 186318 310040 186374 310049
rect 186318 309975 186374 309984
rect 186320 309120 186372 309126
rect 186320 309062 186372 309068
rect 186332 308961 186360 309062
rect 186412 309052 186464 309058
rect 186412 308994 186464 309000
rect 186318 308952 186374 308961
rect 186318 308887 186374 308896
rect 186424 307873 186452 308994
rect 186410 307864 186466 307873
rect 186410 307799 186466 307808
rect 186320 307760 186372 307766
rect 186320 307702 186372 307708
rect 186332 306785 186360 307702
rect 186318 306776 186374 306785
rect 186318 306711 186374 306720
rect 186320 306332 186372 306338
rect 186320 306274 186372 306280
rect 186332 305833 186360 306274
rect 186318 305824 186374 305833
rect 186318 305759 186374 305768
rect 186412 304972 186464 304978
rect 186412 304914 186464 304920
rect 186424 303657 186452 304914
rect 186688 304904 186740 304910
rect 186688 304846 186740 304852
rect 186700 304745 186728 304846
rect 186686 304736 186742 304745
rect 186686 304671 186742 304680
rect 186410 303648 186466 303657
rect 186320 303612 186372 303618
rect 186410 303583 186466 303592
rect 186320 303554 186372 303560
rect 186332 302569 186360 303554
rect 186318 302560 186374 302569
rect 186318 302495 186374 302504
rect 186320 302184 186372 302190
rect 186320 302126 186372 302132
rect 186332 301617 186360 302126
rect 186318 301608 186374 301617
rect 186318 301543 186374 301552
rect 186320 300824 186372 300830
rect 186320 300766 186372 300772
rect 186332 300529 186360 300766
rect 186318 300520 186374 300529
rect 186318 300455 186374 300464
rect 186320 299464 186372 299470
rect 186318 299432 186320 299441
rect 186372 299432 186374 299441
rect 186318 299367 186374 299376
rect 186412 299396 186464 299402
rect 186412 299338 186464 299344
rect 186424 298353 186452 299338
rect 186410 298344 186466 298353
rect 186410 298279 186466 298288
rect 186320 298104 186372 298110
rect 186320 298046 186372 298052
rect 186332 297401 186360 298046
rect 186318 297392 186374 297401
rect 186318 297327 186374 297336
rect 186320 296676 186372 296682
rect 186320 296618 186372 296624
rect 186332 296313 186360 296618
rect 186318 296304 186374 296313
rect 186318 296239 186374 296248
rect 186320 295316 186372 295322
rect 186320 295258 186372 295264
rect 186332 295225 186360 295258
rect 186412 295248 186464 295254
rect 186318 295216 186374 295225
rect 186412 295190 186464 295196
rect 186318 295151 186374 295160
rect 186424 294273 186452 295190
rect 186410 294264 186466 294273
rect 186410 294199 186466 294208
rect 186320 293956 186372 293962
rect 186320 293898 186372 293904
rect 186332 293185 186360 293898
rect 186318 293176 186374 293185
rect 186318 293111 186374 293120
rect 186320 292528 186372 292534
rect 186320 292470 186372 292476
rect 186332 292097 186360 292470
rect 186318 292088 186374 292097
rect 186318 292023 186374 292032
rect 186412 291168 186464 291174
rect 186412 291110 186464 291116
rect 186320 291100 186372 291106
rect 186320 291042 186372 291048
rect 186332 291009 186360 291042
rect 186318 291000 186374 291009
rect 186318 290935 186374 290944
rect 186424 290057 186452 291110
rect 186410 290048 186466 290057
rect 186410 289983 186466 289992
rect 186320 289808 186372 289814
rect 186320 289750 186372 289756
rect 186332 288969 186360 289750
rect 186318 288960 186374 288969
rect 186318 288895 186374 288904
rect 186320 288380 186372 288386
rect 186320 288322 186372 288328
rect 186332 287881 186360 288322
rect 186318 287872 186374 287881
rect 186318 287807 186374 287816
rect 186320 287020 186372 287026
rect 186320 286962 186372 286968
rect 186332 286793 186360 286962
rect 186412 286952 186464 286958
rect 186412 286894 186464 286900
rect 186318 286784 186374 286793
rect 186318 286719 186374 286728
rect 186424 285841 186452 286894
rect 186410 285832 186466 285841
rect 186410 285767 186466 285776
rect 186320 285660 186372 285666
rect 186320 285602 186372 285608
rect 186332 284753 186360 285602
rect 186318 284744 186374 284753
rect 186318 284679 186374 284688
rect 186320 284300 186372 284306
rect 186320 284242 186372 284248
rect 186332 283665 186360 284242
rect 186318 283656 186374 283665
rect 186318 283591 186374 283600
rect 186320 282872 186372 282878
rect 186320 282814 186372 282820
rect 186332 282577 186360 282814
rect 186412 282804 186464 282810
rect 186412 282746 186464 282752
rect 186318 282568 186374 282577
rect 186318 282503 186374 282512
rect 186424 281625 186452 282746
rect 186410 281616 186466 281625
rect 186410 281551 186466 281560
rect 186320 281512 186372 281518
rect 186320 281454 186372 281460
rect 186332 280537 186360 281454
rect 186318 280528 186374 280537
rect 186318 280463 186374 280472
rect 186320 280152 186372 280158
rect 186320 280094 186372 280100
rect 186332 279449 186360 280094
rect 186318 279440 186374 279449
rect 186318 279375 186374 279384
rect 186320 278724 186372 278730
rect 186320 278666 186372 278672
rect 186332 278361 186360 278666
rect 186318 278352 186374 278361
rect 186318 278287 186374 278296
rect 186318 277400 186374 277409
rect 186318 277335 186320 277344
rect 186372 277335 186374 277344
rect 186320 277306 186372 277312
rect 186412 277296 186464 277302
rect 186412 277238 186464 277244
rect 186424 276321 186452 277238
rect 186410 276312 186466 276321
rect 186410 276247 186466 276256
rect 186320 276004 186372 276010
rect 186320 275946 186372 275952
rect 186332 275233 186360 275946
rect 186318 275224 186374 275233
rect 186318 275159 186374 275168
rect 186320 274644 186372 274650
rect 186320 274586 186372 274592
rect 186332 274145 186360 274586
rect 186318 274136 186374 274145
rect 186318 274071 186374 274080
rect 186320 273216 186372 273222
rect 186318 273184 186320 273193
rect 186372 273184 186374 273193
rect 186318 273119 186374 273128
rect 186412 273148 186464 273154
rect 186412 273090 186464 273096
rect 186424 272105 186452 273090
rect 186410 272096 186466 272105
rect 186410 272031 186466 272040
rect 186320 271856 186372 271862
rect 186320 271798 186372 271804
rect 186332 271017 186360 271798
rect 186318 271008 186374 271017
rect 186318 270943 186374 270952
rect 186320 270496 186372 270502
rect 186320 270438 186372 270444
rect 186332 269929 186360 270438
rect 186318 269920 186374 269929
rect 186318 269855 186374 269864
rect 186320 269068 186372 269074
rect 186320 269010 186372 269016
rect 186332 267889 186360 269010
rect 186412 269000 186464 269006
rect 186410 268968 186412 268977
rect 186464 268968 186466 268977
rect 186410 268903 186466 268912
rect 186318 267880 186374 267889
rect 186318 267815 186374 267824
rect 186320 267708 186372 267714
rect 186320 267650 186372 267656
rect 186332 266801 186360 267650
rect 186318 266792 186374 266801
rect 186318 266727 186374 266736
rect 186320 266348 186372 266354
rect 186320 266290 186372 266296
rect 186332 265713 186360 266290
rect 186318 265704 186374 265713
rect 186318 265639 186374 265648
rect 186320 264920 186372 264926
rect 186320 264862 186372 264868
rect 186332 264761 186360 264862
rect 186412 264852 186464 264858
rect 186412 264794 186464 264800
rect 186318 264752 186374 264761
rect 186318 264687 186374 264696
rect 186424 263673 186452 264794
rect 186410 263664 186466 263673
rect 186410 263599 186466 263608
rect 186320 263560 186372 263566
rect 186320 263502 186372 263508
rect 186332 262585 186360 263502
rect 186318 262576 186374 262585
rect 186318 262511 186374 262520
rect 186320 262200 186372 262206
rect 186320 262142 186372 262148
rect 186332 261633 186360 262142
rect 186318 261624 186374 261633
rect 186318 261559 186374 261568
rect 186320 260840 186372 260846
rect 186320 260782 186372 260788
rect 186332 260545 186360 260782
rect 186318 260536 186374 260545
rect 186318 260471 186374 260480
rect 186410 259448 186466 259457
rect 186320 259412 186372 259418
rect 186410 259383 186466 259392
rect 186320 259354 186372 259360
rect 186332 258369 186360 259354
rect 186424 259350 186452 259383
rect 186412 259344 186464 259350
rect 186412 259286 186464 259292
rect 186318 258360 186374 258369
rect 186318 258295 186374 258304
rect 186320 258052 186372 258058
rect 186320 257994 186372 258000
rect 186332 257417 186360 257994
rect 186318 257408 186374 257417
rect 186318 257343 186374 257352
rect 186320 256692 186372 256698
rect 186320 256634 186372 256640
rect 186332 256329 186360 256634
rect 186318 256320 186374 256329
rect 186318 256255 186374 256264
rect 186320 255264 186372 255270
rect 186318 255232 186320 255241
rect 186372 255232 186374 255241
rect 186318 255167 186374 255176
rect 186412 255196 186464 255202
rect 186412 255138 186464 255144
rect 186424 254153 186452 255138
rect 186410 254144 186466 254153
rect 186410 254079 186466 254088
rect 186320 253904 186372 253910
rect 186320 253846 186372 253852
rect 186332 253201 186360 253846
rect 186318 253192 186374 253201
rect 186318 253127 186374 253136
rect 186320 252544 186372 252550
rect 186320 252486 186372 252492
rect 186332 252113 186360 252486
rect 186318 252104 186374 252113
rect 186318 252039 186374 252048
rect 186320 251184 186372 251190
rect 186320 251126 186372 251132
rect 186332 251025 186360 251126
rect 186412 251116 186464 251122
rect 186412 251058 186464 251064
rect 186318 251016 186374 251025
rect 186318 250951 186374 250960
rect 186424 249937 186452 251058
rect 186410 249928 186466 249937
rect 186410 249863 186466 249872
rect 186320 249756 186372 249762
rect 186320 249698 186372 249704
rect 186332 248985 186360 249698
rect 186318 248976 186374 248985
rect 186318 248911 186374 248920
rect 186320 248396 186372 248402
rect 186320 248338 186372 248344
rect 186332 247897 186360 248338
rect 186318 247888 186374 247897
rect 186318 247823 186374 247832
rect 186320 247036 186372 247042
rect 186320 246978 186372 246984
rect 186332 246809 186360 246978
rect 186412 246968 186464 246974
rect 186412 246910 186464 246916
rect 186318 246800 186374 246809
rect 186318 246735 186374 246744
rect 186424 245721 186452 246910
rect 186410 245712 186466 245721
rect 186410 245647 186466 245656
rect 186320 245608 186372 245614
rect 186320 245550 186372 245556
rect 186332 244769 186360 245550
rect 186318 244760 186374 244769
rect 186318 244695 186374 244704
rect 186320 244248 186372 244254
rect 186320 244190 186372 244196
rect 186332 243681 186360 244190
rect 186318 243672 186374 243681
rect 186318 243607 186374 243616
rect 186320 242888 186372 242894
rect 186320 242830 186372 242836
rect 186332 242593 186360 242830
rect 186318 242584 186374 242593
rect 186318 242519 186374 242528
rect 186318 241496 186374 241505
rect 186318 241431 186374 241440
rect 186412 241460 186464 241466
rect 186332 241398 186360 241431
rect 186412 241402 186464 241408
rect 186320 241392 186372 241398
rect 186320 241334 186372 241340
rect 186424 240553 186452 241402
rect 186410 240544 186466 240553
rect 186410 240479 186466 240488
rect 186320 240100 186372 240106
rect 186320 240042 186372 240048
rect 186332 239465 186360 240042
rect 186318 239456 186374 239465
rect 186318 239391 186374 239400
rect 186320 238740 186372 238746
rect 186320 238682 186372 238688
rect 186332 238377 186360 238682
rect 186318 238368 186374 238377
rect 186318 238303 186374 238312
rect 186320 237380 186372 237386
rect 186320 237322 186372 237328
rect 186332 237289 186360 237322
rect 186412 237312 186464 237318
rect 186318 237280 186374 237289
rect 186412 237254 186464 237260
rect 186318 237215 186374 237224
rect 186424 236337 186452 237254
rect 186410 236328 186466 236337
rect 186410 236263 186466 236272
rect 186320 235952 186372 235958
rect 186320 235894 186372 235900
rect 186332 235249 186360 235894
rect 186318 235240 186374 235249
rect 186318 235175 186374 235184
rect 186320 234592 186372 234598
rect 186320 234534 186372 234540
rect 186332 234161 186360 234534
rect 186318 234152 186374 234161
rect 186318 234087 186374 234096
rect 186320 233232 186372 233238
rect 186320 233174 186372 233180
rect 186332 233073 186360 233174
rect 186412 233164 186464 233170
rect 186412 233106 186464 233112
rect 186318 233064 186374 233073
rect 186318 232999 186374 233008
rect 186424 232121 186452 233106
rect 186410 232112 186466 232121
rect 186410 232047 186466 232056
rect 186320 231804 186372 231810
rect 186320 231746 186372 231752
rect 186332 231033 186360 231746
rect 186318 231024 186374 231033
rect 186318 230959 186374 230968
rect 186320 230444 186372 230450
rect 186320 230386 186372 230392
rect 186332 229945 186360 230386
rect 186318 229936 186374 229945
rect 186318 229871 186374 229880
rect 186320 229084 186372 229090
rect 186320 229026 186372 229032
rect 186332 228993 186360 229026
rect 186412 229016 186464 229022
rect 186318 228984 186374 228993
rect 186412 228958 186464 228964
rect 186318 228919 186374 228928
rect 186424 227905 186452 228958
rect 186410 227896 186466 227905
rect 186410 227831 186466 227840
rect 186320 227724 186372 227730
rect 186320 227666 186372 227672
rect 186332 226817 186360 227666
rect 186318 226808 186374 226817
rect 186318 226743 186374 226752
rect 186320 226296 186372 226302
rect 186320 226238 186372 226244
rect 186332 225729 186360 226238
rect 186318 225720 186374 225729
rect 186318 225655 186374 225664
rect 186320 224936 186372 224942
rect 186320 224878 186372 224884
rect 186332 224777 186360 224878
rect 186412 224868 186464 224874
rect 186412 224810 186464 224816
rect 186318 224768 186374 224777
rect 186318 224703 186374 224712
rect 186424 223689 186452 224810
rect 186410 223680 186466 223689
rect 186410 223615 186466 223624
rect 186320 223576 186372 223582
rect 186320 223518 186372 223524
rect 186332 222601 186360 223518
rect 186318 222592 186374 222601
rect 186318 222527 186374 222536
rect 186320 222148 186372 222154
rect 186320 222090 186372 222096
rect 186332 221513 186360 222090
rect 186318 221504 186374 221513
rect 186318 221439 186374 221448
rect 186412 220788 186464 220794
rect 186412 220730 186464 220736
rect 186424 219473 186452 220730
rect 186504 220720 186556 220726
rect 186504 220662 186556 220668
rect 186516 220561 186544 220662
rect 186502 220552 186558 220561
rect 186502 220487 186558 220496
rect 186410 219464 186466 219473
rect 186320 219428 186372 219434
rect 186410 219399 186466 219408
rect 186320 219370 186372 219376
rect 186332 218385 186360 219370
rect 186318 218376 186374 218385
rect 186318 218311 186374 218320
rect 186320 218000 186372 218006
rect 186320 217942 186372 217948
rect 186332 217297 186360 217942
rect 186318 217288 186374 217297
rect 186318 217223 186374 217232
rect 186320 216640 186372 216646
rect 186320 216582 186372 216588
rect 186332 216345 186360 216582
rect 186318 216336 186374 216345
rect 186318 216271 186374 216280
rect 186412 215280 186464 215286
rect 186318 215248 186374 215257
rect 186412 215222 186464 215228
rect 186318 215183 186320 215192
rect 186372 215183 186374 215192
rect 186320 215154 186372 215160
rect 186424 214169 186452 215222
rect 186410 214160 186466 214169
rect 186410 214095 186466 214104
rect 186320 213920 186372 213926
rect 186320 213862 186372 213868
rect 186332 213081 186360 213862
rect 186318 213072 186374 213081
rect 186318 213007 186374 213016
rect 186320 212492 186372 212498
rect 186320 212434 186372 212440
rect 186332 212129 186360 212434
rect 186318 212120 186374 212129
rect 186318 212055 186374 212064
rect 186320 211132 186372 211138
rect 186320 211074 186372 211080
rect 186332 211041 186360 211074
rect 186412 211064 186464 211070
rect 186318 211032 186374 211041
rect 186412 211006 186464 211012
rect 186318 210967 186374 210976
rect 186424 209953 186452 211006
rect 186410 209944 186466 209953
rect 186410 209879 186466 209888
rect 186320 209772 186372 209778
rect 186320 209714 186372 209720
rect 186332 208865 186360 209714
rect 186318 208856 186374 208865
rect 186318 208791 186374 208800
rect 186320 208344 186372 208350
rect 186320 208286 186372 208292
rect 186332 207913 186360 208286
rect 186318 207904 186374 207913
rect 186318 207839 186374 207848
rect 186320 206984 186372 206990
rect 186320 206926 186372 206932
rect 186332 205737 186360 206926
rect 186412 206916 186464 206922
rect 186412 206858 186464 206864
rect 186424 206825 186452 206858
rect 186410 206816 186466 206825
rect 186410 206751 186466 206760
rect 186318 205728 186374 205737
rect 186318 205663 186374 205672
rect 186320 205624 186372 205630
rect 186320 205566 186372 205572
rect 186332 204649 186360 205566
rect 186318 204640 186374 204649
rect 186318 204575 186374 204584
rect 186320 204264 186372 204270
rect 186320 204206 186372 204212
rect 186332 203697 186360 204206
rect 186318 203688 186374 203697
rect 186318 203623 186374 203632
rect 186412 202836 186464 202842
rect 186412 202778 186464 202784
rect 186320 202768 186372 202774
rect 186320 202710 186372 202716
rect 186332 202609 186360 202710
rect 186318 202600 186374 202609
rect 186318 202535 186374 202544
rect 186424 201521 186452 202778
rect 186410 201512 186466 201521
rect 186320 201476 186372 201482
rect 186410 201447 186466 201456
rect 186320 201418 186372 201424
rect 186332 200569 186360 201418
rect 186318 200560 186374 200569
rect 186318 200495 186374 200504
rect 186228 197804 186280 197810
rect 186228 197746 186280 197752
rect 186884 180130 186912 413063
rect 187068 402665 187096 420106
rect 187332 420028 187384 420034
rect 187332 419970 187384 419976
rect 187148 419960 187200 419966
rect 187148 419902 187200 419908
rect 187054 402656 187110 402665
rect 187054 402591 187110 402600
rect 187160 394233 187188 419902
rect 187240 419892 187292 419898
rect 187240 419834 187292 419840
rect 187252 413930 187280 419834
rect 187344 414066 187372 419970
rect 187424 419552 187476 419558
rect 187424 419494 187476 419500
rect 187436 414186 187464 419494
rect 187528 414225 187556 420242
rect 187606 416392 187662 416401
rect 187606 416327 187662 416336
rect 187514 414216 187570 414225
rect 187424 414180 187476 414186
rect 187514 414151 187570 414160
rect 187424 414122 187476 414128
rect 187344 414038 187556 414066
rect 187424 413976 187476 413982
rect 187252 413902 187372 413930
rect 187424 413918 187476 413924
rect 187240 413840 187292 413846
rect 187240 413782 187292 413788
rect 187146 394224 187202 394233
rect 187146 394159 187202 394168
rect 187252 390017 187280 413782
rect 187344 396273 187372 413902
rect 187330 396264 187386 396273
rect 187330 396199 187386 396208
rect 187238 390008 187294 390017
rect 187238 389943 187294 389952
rect 187330 386880 187386 386889
rect 187330 386815 187386 386824
rect 187238 381576 187294 381585
rect 187238 381511 187294 381520
rect 187146 380488 187202 380497
rect 187146 380423 187202 380432
rect 187160 191146 187188 380423
rect 187148 191140 187200 191146
rect 187148 191082 187200 191088
rect 187252 186998 187280 381511
rect 187240 186992 187292 186998
rect 187240 186934 187292 186940
rect 186872 180124 186924 180130
rect 186872 180066 186924 180072
rect 187344 155242 187372 386815
rect 187436 384713 187464 413918
rect 187528 407969 187556 414038
rect 187514 407960 187570 407969
rect 187514 407895 187570 407904
rect 187514 400480 187570 400489
rect 187514 400415 187570 400424
rect 187422 384704 187478 384713
rect 187422 384639 187478 384648
rect 187424 358760 187476 358766
rect 187424 358702 187476 358708
rect 187436 358465 187464 358702
rect 187422 358456 187478 358465
rect 187422 358391 187478 358400
rect 187528 184210 187556 400415
rect 187516 184204 187568 184210
rect 187516 184146 187568 184152
rect 187620 177342 187648 416327
rect 188356 199102 188384 496878
rect 188896 422340 188948 422346
rect 188896 422282 188948 422288
rect 188436 409148 188488 409154
rect 188436 409090 188488 409096
rect 188344 199096 188396 199102
rect 188344 199038 188396 199044
rect 188448 198558 188476 409090
rect 188528 407788 188580 407794
rect 188528 407730 188580 407736
rect 188436 198552 188488 198558
rect 188436 198494 188488 198500
rect 188540 198490 188568 407730
rect 188802 405784 188858 405793
rect 188802 405719 188858 405728
rect 188710 404696 188766 404705
rect 188710 404631 188766 404640
rect 188528 198484 188580 198490
rect 188528 198426 188580 198432
rect 188724 191214 188752 404631
rect 188712 191208 188764 191214
rect 188712 191150 188764 191156
rect 188816 182850 188844 405719
rect 188908 197878 188936 422282
rect 189356 419688 189408 419694
rect 189356 419630 189408 419636
rect 189080 419620 189132 419626
rect 189080 419562 189132 419568
rect 188986 397352 189042 397361
rect 188986 397287 189042 397296
rect 188896 197872 188948 197878
rect 188896 197814 188948 197820
rect 188804 182844 188856 182850
rect 188804 182786 188856 182792
rect 187608 177336 187660 177342
rect 187608 177278 187660 177284
rect 187332 155236 187384 155242
rect 187332 155178 187384 155184
rect 189000 149734 189028 397287
rect 189092 392057 189120 419562
rect 189170 408912 189226 408921
rect 189170 408847 189226 408856
rect 189078 392048 189134 392057
rect 189078 391983 189134 391992
rect 189078 382664 189134 382673
rect 189078 382599 189134 382608
rect 188988 149728 189040 149734
rect 188988 149670 189040 149676
rect 189092 144226 189120 382599
rect 189184 189786 189212 408847
rect 189262 399528 189318 399537
rect 189262 399463 189318 399472
rect 189276 192506 189304 399463
rect 189368 398449 189396 419630
rect 189354 398440 189410 398449
rect 189354 398375 189410 398384
rect 189736 199170 189764 497014
rect 189724 199164 189776 199170
rect 189724 199106 189776 199112
rect 189828 199034 189856 497082
rect 190368 420232 190420 420238
rect 190368 420174 190420 420180
rect 190380 417897 190408 420174
rect 190472 419914 190500 507826
rect 191852 441614 191880 509254
rect 193220 496120 193272 496126
rect 193220 496062 193272 496068
rect 193232 441614 193260 496062
rect 195980 491972 196032 491978
rect 195980 491914 196032 491920
rect 195992 441614 196020 491914
rect 204904 490612 204956 490618
rect 204904 490554 204956 490560
rect 198740 486532 198792 486538
rect 198740 486474 198792 486480
rect 198752 441614 198780 486474
rect 191852 441586 192064 441614
rect 193232 441586 193904 441614
rect 195992 441586 196112 441614
rect 198752 441586 199056 441614
rect 190736 420096 190788 420102
rect 190734 420064 190736 420073
rect 190788 420064 190790 420073
rect 190734 419999 190790 420008
rect 192036 419914 192064 441586
rect 193876 419914 193904 441586
rect 196084 419914 196112 441586
rect 198004 425740 198056 425746
rect 198004 425682 198056 425688
rect 198016 423434 198044 425682
rect 198004 423428 198056 423434
rect 198004 423370 198056 423376
rect 198016 419914 198044 423370
rect 190472 419886 190854 419914
rect 192036 419886 192510 419914
rect 193876 419886 194258 419914
rect 196006 419886 196112 419914
rect 197754 419886 198044 419914
rect 199028 419914 199056 441586
rect 200856 428596 200908 428602
rect 200856 428538 200908 428544
rect 200868 419914 200896 428538
rect 203248 424380 203300 424386
rect 203248 424322 203300 424328
rect 203260 419914 203288 424322
rect 204916 423502 204944 490554
rect 205640 480956 205692 480962
rect 205640 480898 205692 480904
rect 205652 441614 205680 480898
rect 207032 441614 207060 527138
rect 209780 493332 209832 493338
rect 209780 493274 209832 493280
rect 205652 441586 206048 441614
rect 207032 441586 207888 441614
rect 204904 423496 204956 423502
rect 204904 423438 204956 423444
rect 204916 419914 204944 423438
rect 199028 419886 199502 419914
rect 200868 419886 201250 419914
rect 202998 419886 203288 419914
rect 204746 419886 204944 419914
rect 206020 419914 206048 441586
rect 207860 419914 207888 441586
rect 209792 419914 209820 493274
rect 211804 487824 211856 487830
rect 211804 487766 211856 487772
rect 211816 423570 211844 487766
rect 212540 471300 212592 471306
rect 212540 471242 212592 471248
rect 212552 441614 212580 471242
rect 213932 441614 213960 529926
rect 216680 489184 216732 489190
rect 216680 489126 216732 489132
rect 212552 441586 213040 441614
rect 213932 441586 214880 441614
rect 211804 423564 211856 423570
rect 211804 423506 211856 423512
rect 211816 419914 211844 423506
rect 206020 419886 206494 419914
rect 207860 419886 208242 419914
rect 209792 419886 209990 419914
rect 211738 419886 211844 419914
rect 213012 419914 213040 441586
rect 214852 419914 214880 441586
rect 216692 419914 216720 489126
rect 219440 450628 219492 450634
rect 219440 450570 219492 450576
rect 219452 441614 219480 450570
rect 222212 441614 222240 529994
rect 224960 453348 225012 453354
rect 224960 453290 225012 453296
rect 224972 441614 225000 453290
rect 226352 441614 226380 532714
rect 230480 467152 230532 467158
rect 230480 467094 230532 467100
rect 219452 441586 220032 441614
rect 222212 441586 222332 441614
rect 224972 441586 225368 441614
rect 226352 441586 227024 441614
rect 218612 426148 218664 426154
rect 218612 426090 218664 426096
rect 218624 423638 218652 426090
rect 218612 423632 218664 423638
rect 218612 423574 218664 423580
rect 218624 419914 218652 423574
rect 220004 419914 220032 441586
rect 222304 419914 222332 441586
rect 223580 425808 223632 425814
rect 223580 425750 223632 425756
rect 213012 419886 213486 419914
rect 214852 419886 215234 419914
rect 216692 419886 216982 419914
rect 218624 419886 218730 419914
rect 220004 419886 220478 419914
rect 222226 419886 222332 419914
rect 223592 419914 223620 425750
rect 225340 419914 225368 441586
rect 226996 419914 227024 441586
rect 229100 425876 229152 425882
rect 229100 425818 229152 425824
rect 229112 419914 229140 425818
rect 230492 419914 230520 467094
rect 231872 441614 231900 532782
rect 236000 454708 236052 454714
rect 236000 454650 236052 454656
rect 231872 441586 232360 441614
rect 232332 419914 232360 441586
rect 233976 425944 234028 425950
rect 233976 425886 234028 425892
rect 233988 419914 234016 425886
rect 236012 419914 236040 454650
rect 237392 441614 237420 535434
rect 237392 441586 237512 441614
rect 237484 419914 237512 441586
rect 239312 426012 239364 426018
rect 239312 425954 239364 425960
rect 239324 419914 239352 425954
rect 241336 423156 241388 423162
rect 241336 423098 241388 423104
rect 241348 419914 241376 423098
rect 242912 419914 242940 536794
rect 396630 535936 396686 535945
rect 396630 535871 396686 535880
rect 396644 535498 396672 535871
rect 396632 535492 396684 535498
rect 396632 535434 396684 535440
rect 396722 533760 396778 533769
rect 396722 533695 396778 533704
rect 396736 532846 396764 533695
rect 396724 532840 396776 532846
rect 396630 532808 396686 532817
rect 396724 532782 396776 532788
rect 396630 532743 396632 532752
rect 396684 532743 396686 532752
rect 396632 532714 396684 532720
rect 396722 531040 396778 531049
rect 396722 530975 396778 530984
rect 396736 530058 396764 530975
rect 396724 530052 396776 530058
rect 396724 529994 396776 530000
rect 396632 529984 396684 529990
rect 396630 529952 396632 529961
rect 396684 529952 396686 529961
rect 396630 529887 396686 529896
rect 396630 528184 396686 528193
rect 396630 528119 396686 528128
rect 396644 527202 396672 528119
rect 396632 527196 396684 527202
rect 396632 527138 396684 527144
rect 396354 509960 396410 509969
rect 396354 509895 396410 509904
rect 396368 509318 396396 509895
rect 396356 509312 396408 509318
rect 396356 509254 396408 509260
rect 397366 508328 397422 508337
rect 397366 508263 397422 508272
rect 396630 508056 396686 508065
rect 396630 507991 396686 508000
rect 396644 507890 396672 507991
rect 396632 507884 396684 507890
rect 396632 507826 396684 507832
rect 338120 498840 338172 498846
rect 338120 498782 338172 498788
rect 284944 496936 284996 496942
rect 284944 496878 284996 496884
rect 255320 494828 255372 494834
rect 255320 494770 255372 494776
rect 252560 485172 252612 485178
rect 252560 485114 252612 485120
rect 245660 457496 245712 457502
rect 245660 457438 245712 457444
rect 245672 441614 245700 457438
rect 252572 441614 252600 485114
rect 245672 441586 246344 441614
rect 252572 441586 253336 441614
rect 244464 426080 244516 426086
rect 244464 426022 244516 426028
rect 244476 419914 244504 426022
rect 246316 419914 246344 441586
rect 251456 430024 251508 430030
rect 251456 429966 251508 429972
rect 248512 426216 248564 426222
rect 248512 426158 248564 426164
rect 248524 419914 248552 426158
rect 250536 423224 250588 423230
rect 250536 423166 250588 423172
rect 250548 419914 250576 423166
rect 223592 419886 223974 419914
rect 225340 419886 225722 419914
rect 226996 419886 227470 419914
rect 229112 419886 229218 419914
rect 230492 419886 230966 419914
rect 232332 419886 232714 419914
rect 233988 419886 234462 419914
rect 236012 419886 236210 419914
rect 237484 419886 237958 419914
rect 239324 419886 239706 419914
rect 241348 419886 241454 419914
rect 242912 419886 243202 419914
rect 244476 419886 244950 419914
rect 246316 419886 246698 419914
rect 248446 419886 248552 419914
rect 250194 419886 250576 419914
rect 251468 419914 251496 429966
rect 253308 419914 253336 441586
rect 255332 419914 255360 494770
rect 263600 483676 263652 483682
rect 263600 483618 263652 483624
rect 263612 441614 263640 483618
rect 281540 482384 281592 482390
rect 281540 482326 281592 482332
rect 273260 478168 273312 478174
rect 273260 478110 273312 478116
rect 273272 441614 273300 478110
rect 281552 441614 281580 482326
rect 284956 450634 284984 496878
rect 331220 482316 331272 482322
rect 331220 482258 331272 482264
rect 302240 479596 302292 479602
rect 302240 479538 302292 479544
rect 288440 476876 288492 476882
rect 288440 476818 288492 476824
rect 284944 450628 284996 450634
rect 284944 450570 284996 450576
rect 263612 441586 263824 441614
rect 273272 441586 274128 441614
rect 281552 441586 281672 441614
rect 262220 434104 262272 434110
rect 262220 434046 262272 434052
rect 258448 431384 258500 431390
rect 258448 431326 258500 431332
rect 256792 426284 256844 426290
rect 256792 426226 256844 426232
rect 256804 419914 256832 426226
rect 258460 419914 258488 431326
rect 260288 427168 260340 427174
rect 260288 427110 260340 427116
rect 260300 419914 260328 427110
rect 262232 419914 262260 434046
rect 263796 419914 263824 441586
rect 269120 435464 269172 435470
rect 269120 435406 269172 435412
rect 265440 432744 265492 432750
rect 265440 432686 265492 432692
rect 265452 419914 265480 432686
rect 267096 427236 267148 427242
rect 267096 427178 267148 427184
rect 267108 419914 267136 427178
rect 269132 419914 269160 435406
rect 270592 427304 270644 427310
rect 270592 427246 270644 427252
rect 270604 419914 270632 427246
rect 273168 424448 273220 424454
rect 273168 424390 273220 424396
rect 273180 419914 273208 424390
rect 251468 419886 251942 419914
rect 253308 419886 253690 419914
rect 255332 419886 255438 419914
rect 256804 419886 257186 419914
rect 258460 419886 258934 419914
rect 260300 419886 260682 419914
rect 262232 419886 262430 419914
rect 263796 419886 264178 419914
rect 265452 419886 265834 419914
rect 267108 419886 267582 419914
rect 269132 419886 269330 419914
rect 270604 419886 271078 419914
rect 272826 419886 273208 419914
rect 274100 419914 274128 441586
rect 277584 427372 277636 427378
rect 277584 427314 277636 427320
rect 276664 424584 276716 424590
rect 276664 424526 276716 424532
rect 276676 419914 276704 424526
rect 274100 419886 274574 419914
rect 276322 419886 276704 419914
rect 277596 419914 277624 427314
rect 279976 424516 280028 424522
rect 279976 424458 280028 424464
rect 279988 419914 280016 424458
rect 281644 419914 281672 441586
rect 284576 427440 284628 427446
rect 284576 427382 284628 427388
rect 283656 424720 283708 424726
rect 283656 424662 283708 424668
rect 283668 419914 283696 424662
rect 277596 419886 278070 419914
rect 279818 419886 280016 419914
rect 281566 419886 281672 419914
rect 283314 419886 283696 419914
rect 284588 419914 284616 427382
rect 286968 424652 287020 424658
rect 286968 424594 287020 424600
rect 286980 419914 287008 424594
rect 284588 419886 285062 419914
rect 286810 419886 287008 419914
rect 288452 419914 288480 476818
rect 298100 475380 298152 475386
rect 298100 475322 298152 475328
rect 291200 472728 291252 472734
rect 291200 472670 291252 472676
rect 291212 441614 291240 472670
rect 295340 446480 295392 446486
rect 295340 446422 295392 446428
rect 291212 441586 291608 441614
rect 290648 424856 290700 424862
rect 290648 424798 290700 424804
rect 290660 419914 290688 424798
rect 288452 419886 288558 419914
rect 290306 419886 290688 419914
rect 291580 419914 291608 441586
rect 293868 424788 293920 424794
rect 293868 424730 293920 424736
rect 293880 419914 293908 424730
rect 291580 419886 292054 419914
rect 293802 419886 293908 419914
rect 295352 419914 295380 446422
rect 298112 441614 298140 475322
rect 298112 441586 298600 441614
rect 297640 424924 297692 424930
rect 297640 424866 297692 424872
rect 297652 419914 297680 424866
rect 295352 419886 295550 419914
rect 297298 419886 297680 419914
rect 298572 419914 298600 441586
rect 300676 424992 300728 424998
rect 300676 424934 300728 424940
rect 300688 419914 300716 424934
rect 302252 419914 302280 479538
rect 305000 474088 305052 474094
rect 305000 474030 305052 474036
rect 305012 441614 305040 474030
rect 309140 469872 309192 469878
rect 309140 469814 309192 469820
rect 305012 441586 305592 441614
rect 303896 436892 303948 436898
rect 303896 436834 303948 436840
rect 303908 419914 303936 436834
rect 305564 419914 305592 441586
rect 307852 438252 307904 438258
rect 307852 438194 307904 438200
rect 307864 419914 307892 438194
rect 298572 419886 299046 419914
rect 300688 419886 300794 419914
rect 302252 419886 302542 419914
rect 303908 419886 304290 419914
rect 305564 419886 306038 419914
rect 307786 419886 307892 419914
rect 309152 419914 309180 469814
rect 316040 465724 316092 465730
rect 316040 465666 316092 465672
rect 311900 447908 311952 447914
rect 311900 447850 311952 447856
rect 311912 441614 311940 447850
rect 311912 441586 312584 441614
rect 310888 440972 310940 440978
rect 310888 440914 310940 440920
rect 310900 419914 310928 440914
rect 312556 419914 312584 441586
rect 314660 439612 314712 439618
rect 314660 439554 314712 439560
rect 314672 419914 314700 439554
rect 316052 419914 316080 465666
rect 325700 451988 325752 451994
rect 325700 451930 325752 451936
rect 322940 450628 322992 450634
rect 322940 450570 322992 450576
rect 318800 449268 318852 449274
rect 318800 449210 318852 449216
rect 317420 442332 317472 442338
rect 317420 442274 317472 442280
rect 317432 441614 317460 442274
rect 318812 441614 318840 449210
rect 321560 443760 321612 443766
rect 321560 443702 321612 443708
rect 317432 441586 317920 441614
rect 318812 441586 319576 441614
rect 317892 419914 317920 441586
rect 319548 419914 319576 441586
rect 321572 419914 321600 443702
rect 322952 441614 322980 450570
rect 324320 445120 324372 445126
rect 324320 445062 324372 445068
rect 324332 441614 324360 445062
rect 325712 441614 325740 451930
rect 331232 441614 331260 482258
rect 338132 441614 338160 498782
rect 359464 496868 359516 496874
rect 359464 496810 359516 496816
rect 340880 494760 340932 494766
rect 340880 494702 340932 494708
rect 340892 441614 340920 494702
rect 342904 474020 342956 474026
rect 342904 473962 342956 473968
rect 322952 441586 323072 441614
rect 324332 441586 324912 441614
rect 325712 441586 326568 441614
rect 331232 441586 331904 441614
rect 338132 441586 338712 441614
rect 340892 441586 341012 441614
rect 323044 419914 323072 441586
rect 324884 419914 324912 441586
rect 326540 419914 326568 441586
rect 330116 423020 330168 423026
rect 330116 422962 330168 422968
rect 329104 421048 329156 421054
rect 329104 420990 329156 420996
rect 329116 419914 329144 420990
rect 309152 419886 309534 419914
rect 310900 419886 311282 419914
rect 312556 419886 313030 419914
rect 314672 419886 314778 419914
rect 316052 419886 316526 419914
rect 317892 419886 318274 419914
rect 319548 419886 320022 419914
rect 321572 419886 321770 419914
rect 323044 419886 323518 419914
rect 324884 419886 325266 419914
rect 326540 419886 327014 419914
rect 328762 419886 329144 419914
rect 330128 419914 330156 422962
rect 331876 419914 331904 441586
rect 335360 434036 335412 434042
rect 335360 433978 335412 433984
rect 334256 422544 334308 422550
rect 334256 422486 334308 422492
rect 334268 419914 334296 422486
rect 330128 419886 330510 419914
rect 331876 419886 332258 419914
rect 334006 419886 334296 419914
rect 335372 419914 335400 433978
rect 338684 419914 338712 441586
rect 340984 419914 341012 441586
rect 342916 423638 342944 473962
rect 356060 472660 356112 472666
rect 356060 472602 356112 472608
rect 356072 441614 356100 472602
rect 356072 441586 356192 441614
rect 342904 423632 342956 423638
rect 342904 423574 342956 423580
rect 344100 423632 344152 423638
rect 344100 423574 344152 423580
rect 335372 419886 335754 419914
rect 338684 419886 339158 419914
rect 340906 419886 341012 419914
rect 344112 419914 344140 423574
rect 351092 422544 351144 422550
rect 351092 422486 351144 422492
rect 347780 422408 347832 422414
rect 347780 422350 347832 422356
rect 346308 421252 346360 421258
rect 346308 421194 346360 421200
rect 346320 419914 346348 421194
rect 344112 419886 344402 419914
rect 346150 419886 346348 419914
rect 347792 419914 347820 422350
rect 349896 421184 349948 421190
rect 349896 421126 349948 421132
rect 349908 419914 349936 421126
rect 351104 420209 351132 422486
rect 351736 422476 351788 422482
rect 351736 422418 351788 422424
rect 351090 420200 351146 420209
rect 351090 420135 351146 420144
rect 351748 419914 351776 422418
rect 353208 422408 353260 422414
rect 353208 422350 353260 422356
rect 353220 419914 353248 422350
rect 355232 421320 355284 421326
rect 355232 421262 355284 421268
rect 355244 419914 355272 421262
rect 347792 419886 347898 419914
rect 349646 419886 349936 419914
rect 351394 419886 351776 419914
rect 353142 419886 353248 419914
rect 354890 419886 355272 419914
rect 356164 419914 356192 441586
rect 357992 440904 358044 440910
rect 357992 440846 358044 440852
rect 358004 419914 358032 440846
rect 359372 427100 359424 427106
rect 359372 427042 359424 427048
rect 359384 422294 359412 427042
rect 359476 423026 359504 496810
rect 383660 485104 383712 485110
rect 383660 485046 383712 485052
rect 378140 445052 378192 445058
rect 378140 444994 378192 445000
rect 378152 441614 378180 444994
rect 383672 441614 383700 485046
rect 389180 479528 389232 479534
rect 389180 479470 389232 479476
rect 389192 441614 389220 479470
rect 378152 441586 379008 441614
rect 383672 441586 384160 441614
rect 389192 441586 389496 441614
rect 363880 423292 363932 423298
rect 363880 423234 363932 423240
rect 359464 423020 359516 423026
rect 359464 422962 359516 422968
rect 362224 422544 362276 422550
rect 362224 422486 362276 422492
rect 360108 422476 360160 422482
rect 360108 422418 360160 422424
rect 359384 422266 359688 422294
rect 359660 419914 359688 422266
rect 360120 421598 360148 422418
rect 360108 421592 360160 421598
rect 360108 421534 360160 421540
rect 362236 419914 362264 422486
rect 363892 419914 363920 423234
rect 365628 422884 365680 422890
rect 365628 422826 365680 422832
rect 365640 419914 365668 422826
rect 374368 422680 374420 422686
rect 374368 422622 374420 422628
rect 370870 422376 370926 422385
rect 368572 422340 368624 422346
rect 370870 422311 370926 422320
rect 368572 422282 368624 422288
rect 367376 420368 367428 420374
rect 367376 420310 367428 420316
rect 367388 419914 367416 420310
rect 356164 419886 356638 419914
rect 358004 419886 358386 419914
rect 359660 419886 360134 419914
rect 361882 419886 362264 419914
rect 363630 419886 363920 419914
rect 365378 419886 365668 419914
rect 367126 419886 367416 419914
rect 368584 419914 368612 422282
rect 370884 419914 370912 422311
rect 374380 419914 374408 422622
rect 377864 422476 377916 422482
rect 377864 422418 377916 422424
rect 376208 421388 376260 421394
rect 376208 421330 376260 421336
rect 376220 419914 376248 421330
rect 377876 419914 377904 422418
rect 368584 419886 368874 419914
rect 370622 419886 370912 419914
rect 374118 419886 374408 419914
rect 375866 419886 376248 419914
rect 377614 419886 377904 419914
rect 378980 419914 379008 441586
rect 382556 422952 382608 422958
rect 382556 422894 382608 422900
rect 380898 421016 380954 421025
rect 380898 420951 380954 420960
rect 380912 419914 380940 420951
rect 382568 419914 382596 422894
rect 384132 419914 384160 441586
rect 386236 422748 386288 422754
rect 386236 422690 386288 422696
rect 386248 419914 386276 422690
rect 388352 421456 388404 421462
rect 388352 421398 388404 421404
rect 388364 419914 388392 421398
rect 378980 419886 379362 419914
rect 380912 419886 381110 419914
rect 382568 419886 382858 419914
rect 384132 419886 384606 419914
rect 386248 419886 386354 419914
rect 388102 419886 388392 419914
rect 389468 419914 389496 441586
rect 394700 438184 394752 438190
rect 394700 438126 394752 438132
rect 391204 421116 391256 421122
rect 391204 421058 391256 421064
rect 393688 421116 393740 421122
rect 393688 421058 393740 421064
rect 391216 419914 391244 421058
rect 393700 419914 393728 421058
rect 389468 419886 389850 419914
rect 391216 419886 391598 419914
rect 393346 419886 393728 419914
rect 394712 419914 394740 438126
rect 397380 428670 397408 508263
rect 419630 498128 419686 498137
rect 419630 498063 419686 498072
rect 433522 498128 433578 498137
rect 433522 498063 433578 498072
rect 440238 498128 440294 498137
rect 440238 498063 440294 498072
rect 454682 498128 454738 498137
rect 454682 498063 454738 498072
rect 455786 498128 455842 498137
rect 462318 498128 462374 498137
rect 455786 498063 455842 498072
rect 457444 498092 457496 498098
rect 410524 497072 410576 497078
rect 410524 497014 410576 497020
rect 409880 486464 409932 486470
rect 409880 486406 409932 486412
rect 407764 476808 407816 476814
rect 407764 476750 407816 476756
rect 397368 428664 397420 428670
rect 397368 428606 397420 428612
rect 407776 423638 407804 476750
rect 409236 450560 409288 450566
rect 409236 450502 409288 450508
rect 407764 423632 407816 423638
rect 407764 423574 407816 423580
rect 408684 423632 408736 423638
rect 408684 423574 408736 423580
rect 396540 423088 396592 423094
rect 396540 423030 396592 423036
rect 396552 419914 396580 423030
rect 403532 423020 403584 423026
rect 403532 422962 403584 422968
rect 398748 422816 398800 422822
rect 398748 422758 398800 422764
rect 398760 419914 398788 422758
rect 400678 421016 400734 421025
rect 400678 420951 400734 420960
rect 402336 420980 402388 420986
rect 400692 419914 400720 420951
rect 402336 420922 402388 420928
rect 402348 419914 402376 420922
rect 394712 419886 395094 419914
rect 396552 419886 396842 419914
rect 398590 419886 398788 419914
rect 400338 419886 400720 419914
rect 402086 419886 402376 419914
rect 403544 419914 403572 422962
rect 405648 422612 405700 422618
rect 405648 422554 405700 422560
rect 405660 419914 405688 422554
rect 407672 422272 407724 422278
rect 407672 422214 407724 422220
rect 407684 419914 407712 422214
rect 403544 419886 403834 419914
rect 405582 419886 405688 419914
rect 407330 419886 407712 419914
rect 408696 419914 408724 423574
rect 409248 422294 409276 450502
rect 409420 436824 409472 436830
rect 409420 436766 409472 436772
rect 409248 422266 409368 422294
rect 408696 419886 409078 419914
rect 372528 419824 372580 419830
rect 372370 419772 372528 419778
rect 372370 419766 372580 419772
rect 372370 419750 372568 419766
rect 190366 417888 190422 417897
rect 190366 417823 190422 417832
rect 409340 413137 409368 422266
rect 409326 413128 409382 413137
rect 409326 413063 409382 413072
rect 409326 410272 409382 410281
rect 409248 410230 409326 410258
rect 189908 405000 189960 405006
rect 189908 404942 189960 404948
rect 189816 199028 189868 199034
rect 189816 198970 189868 198976
rect 189920 197946 189948 404942
rect 190000 401668 190052 401674
rect 190000 401610 190052 401616
rect 190012 198762 190040 401610
rect 191852 200110 191958 200138
rect 195624 200110 195914 200138
rect 198752 200110 199870 200138
rect 203918 200110 204208 200138
rect 207874 200110 208256 200138
rect 190000 198756 190052 198762
rect 190000 198698 190052 198704
rect 189908 197940 189960 197946
rect 189908 197882 189960 197888
rect 189264 192500 189316 192506
rect 189264 192442 189316 192448
rect 189172 189780 189224 189786
rect 189172 189722 189224 189728
rect 189080 144220 189132 144226
rect 189080 144162 189132 144168
rect 188344 142928 188396 142934
rect 188344 142870 188396 142876
rect 176200 142860 176252 142866
rect 176200 142802 176252 142808
rect 176212 142254 176240 142802
rect 176200 142248 176252 142254
rect 176200 142190 176252 142196
rect 173164 141092 173216 141098
rect 173164 141034 173216 141040
rect 176212 139890 176240 142190
rect 188356 142186 188384 142870
rect 191852 142866 191880 200110
rect 195624 199646 195652 200110
rect 194600 199640 194652 199646
rect 194600 199582 194652 199588
rect 195612 199640 195664 199646
rect 195612 199582 195664 199588
rect 194612 198762 194640 199582
rect 194600 198756 194652 198762
rect 194600 198698 194652 198704
rect 194612 143546 194640 198698
rect 194600 143540 194652 143546
rect 194600 143482 194652 143488
rect 195060 143540 195112 143546
rect 195060 143482 195112 143488
rect 192576 143472 192628 143478
rect 192576 143414 192628 143420
rect 192588 142866 192616 143414
rect 195072 142934 195100 143482
rect 195060 142928 195112 142934
rect 195060 142870 195112 142876
rect 191840 142860 191892 142866
rect 191840 142802 191892 142808
rect 192576 142860 192628 142866
rect 192576 142802 192628 142808
rect 188344 142180 188396 142186
rect 188344 142122 188396 142128
rect 188356 139890 188384 142122
rect 198752 141438 198780 200110
rect 200120 197804 200172 197810
rect 200120 197746 200172 197752
rect 198740 141432 198792 141438
rect 198740 141374 198792 141380
rect 176134 139862 176240 139890
rect 188278 139862 188384 139890
rect 200132 139890 200160 197746
rect 204180 193866 204208 200110
rect 208228 198762 208256 200110
rect 211172 200110 211922 200138
rect 215312 200110 215878 200138
rect 219544 200110 219926 200138
rect 223882 200110 224264 200138
rect 208216 198756 208268 198762
rect 208216 198698 208268 198704
rect 204168 193860 204220 193866
rect 204168 193802 204220 193808
rect 211172 146946 211200 200110
rect 212540 197872 212592 197878
rect 212540 197814 212592 197820
rect 211160 146940 211212 146946
rect 211160 146882 211212 146888
rect 212552 139890 212580 197814
rect 215312 145586 215340 200110
rect 219544 198014 219572 200110
rect 224236 198014 224264 200110
rect 227732 200110 227930 200138
rect 235552 200110 235934 200138
rect 239600 200110 239890 200138
rect 243648 200110 243938 200138
rect 247512 200110 247894 200138
rect 251942 200110 252232 200138
rect 219532 198008 219584 198014
rect 219532 197950 219584 197956
rect 224224 198008 224276 198014
rect 224224 197950 224276 197956
rect 227732 197946 227760 200110
rect 235552 198082 235580 200110
rect 239600 199170 239628 200110
rect 239588 199164 239640 199170
rect 239588 199106 239640 199112
rect 243648 198218 243676 200110
rect 243636 198212 243688 198218
rect 243636 198154 243688 198160
rect 247512 198150 247540 200110
rect 247500 198144 247552 198150
rect 247500 198086 247552 198092
rect 235540 198076 235592 198082
rect 235540 198018 235592 198024
rect 252204 197985 252232 200110
rect 255608 200110 255898 200138
rect 259656 200110 259946 200138
rect 263902 200110 264192 200138
rect 255608 198286 255636 200110
rect 259656 199102 259684 200110
rect 261852 199436 261904 199442
rect 261852 199378 261904 199384
rect 259644 199096 259696 199102
rect 259644 199038 259696 199044
rect 255596 198280 255648 198286
rect 255596 198222 255648 198228
rect 261864 198014 261892 199378
rect 264164 198014 264192 200110
rect 267752 200110 267858 200138
rect 271906 200110 272012 200138
rect 267752 198422 267780 200110
rect 271984 198966 272012 200110
rect 274652 200110 275862 200138
rect 279528 200110 279910 200138
rect 282932 200110 283866 200138
rect 287072 200110 287914 200138
rect 291870 200110 292160 200138
rect 295918 200110 296208 200138
rect 271972 198960 272024 198966
rect 271972 198902 272024 198908
rect 267740 198416 267792 198422
rect 267740 198358 267792 198364
rect 261852 198008 261904 198014
rect 252190 197976 252246 197985
rect 227720 197940 227772 197946
rect 261852 197950 261904 197956
rect 264152 198008 264204 198014
rect 264152 197950 264204 197956
rect 252190 197911 252246 197920
rect 227720 197882 227772 197888
rect 260838 192536 260894 192545
rect 224960 192500 225012 192506
rect 260838 192471 260894 192480
rect 224960 192442 225012 192448
rect 224972 151814 225000 192442
rect 236000 191208 236052 191214
rect 236000 191150 236052 191156
rect 236012 151814 236040 191150
rect 248420 189780 248472 189786
rect 248420 189722 248472 189728
rect 248432 151814 248460 189722
rect 260852 151814 260880 192471
rect 274652 178702 274680 200110
rect 279528 198354 279556 200110
rect 279516 198348 279568 198354
rect 279516 198290 279568 198296
rect 280252 198008 280304 198014
rect 280252 197950 280304 197956
rect 274640 178696 274692 178702
rect 274640 178638 274692 178644
rect 224972 151786 225092 151814
rect 236012 151786 236776 151814
rect 248432 151786 249104 151814
rect 260852 151786 261248 151814
rect 215300 145580 215352 145586
rect 215300 145522 215352 145528
rect 225064 139890 225092 151786
rect 200132 139862 200514 139890
rect 212552 139862 212750 139890
rect 224986 139862 225092 139890
rect 236748 139890 236776 151786
rect 249076 139890 249104 151786
rect 261220 139890 261248 151786
rect 280160 146940 280212 146946
rect 280160 146882 280212 146888
rect 274272 142860 274324 142866
rect 274272 142802 274324 142808
rect 274284 139890 274312 142802
rect 236748 139862 237222 139890
rect 249076 139862 249458 139890
rect 261220 139862 261694 139890
rect 273930 139862 274312 139890
rect 279424 49020 279476 49026
rect 279424 48962 279476 48968
rect 278964 37324 279016 37330
rect 278964 37266 279016 37272
rect 174294 30110 174584 30138
rect 182758 30110 183048 30138
rect 191222 30110 191512 30138
rect 199686 30110 199884 30138
rect 208150 30110 208348 30138
rect 171048 28076 171100 28082
rect 171048 28018 171100 28024
rect 174556 28014 174584 30110
rect 183020 29034 183048 30110
rect 183008 29028 183060 29034
rect 183008 28970 183060 28976
rect 191484 28801 191512 30110
rect 191470 28792 191526 28801
rect 191470 28727 191526 28736
rect 199856 28665 199884 30110
rect 208320 29170 208348 30110
rect 216508 30110 216614 30138
rect 224972 30110 225078 30138
rect 233542 30110 233832 30138
rect 242006 30110 242296 30138
rect 250470 30110 250760 30138
rect 258934 30110 259224 30138
rect 208308 29164 208360 29170
rect 208308 29106 208360 29112
rect 216508 29102 216536 30110
rect 216496 29096 216548 29102
rect 216496 29038 216548 29044
rect 199842 28656 199898 28665
rect 199842 28591 199898 28600
rect 224972 28354 225000 30110
rect 233804 28529 233832 30110
rect 233790 28520 233846 28529
rect 233790 28455 233846 28464
rect 242268 28393 242296 30110
rect 242254 28384 242310 28393
rect 224960 28348 225012 28354
rect 250732 28354 250760 30110
rect 242254 28319 242310 28328
rect 250720 28348 250772 28354
rect 224960 28290 225012 28296
rect 250720 28290 250772 28296
rect 259196 28286 259224 30110
rect 267016 30110 267398 30138
rect 275862 30110 275968 30138
rect 259184 28280 259236 28286
rect 259184 28222 259236 28228
rect 267016 28082 267044 30110
rect 275940 28082 275968 30110
rect 278976 29918 279004 37266
rect 279332 32428 279384 32434
rect 279332 32370 279384 32376
rect 278964 29912 279016 29918
rect 278964 29854 279016 29860
rect 279344 29753 279372 32370
rect 279330 29744 279386 29753
rect 279330 29679 279386 29688
rect 279436 29646 279464 48962
rect 279516 41472 279568 41478
rect 279516 41414 279568 41420
rect 279528 29850 279556 41414
rect 280172 37233 280200 146882
rect 280264 92449 280292 197950
rect 282184 192500 282236 192506
rect 282184 192442 282236 192448
rect 281540 149728 281592 149734
rect 281540 149670 281592 149676
rect 281552 133657 281580 149670
rect 281538 133648 281594 133657
rect 281538 133583 281594 133592
rect 280250 92440 280306 92449
rect 280250 92375 280306 92384
rect 282196 78577 282224 192442
rect 282368 189780 282420 189786
rect 282368 189722 282420 189728
rect 282276 149728 282328 149734
rect 282276 149670 282328 149676
rect 282182 78568 282238 78577
rect 282182 78503 282238 78512
rect 282288 64705 282316 149670
rect 282380 106185 282408 189722
rect 282932 151094 282960 200110
rect 284944 193860 284996 193866
rect 284944 193802 284996 193808
rect 282920 151088 282972 151094
rect 282920 151030 282972 151036
rect 282460 146940 282512 146946
rect 282460 146882 282512 146888
rect 282472 119921 282500 146882
rect 282458 119912 282514 119921
rect 282458 119847 282514 119856
rect 282366 106176 282422 106185
rect 282366 106111 282422 106120
rect 282274 64696 282330 64705
rect 282274 64631 282330 64640
rect 280804 57248 280856 57254
rect 280804 57190 280856 57196
rect 280158 37224 280214 37233
rect 280158 37159 280214 37168
rect 279976 34536 280028 34542
rect 279976 34478 280028 34484
rect 279516 29844 279568 29850
rect 279516 29786 279568 29792
rect 279988 29714 280016 34478
rect 280068 31068 280120 31074
rect 280068 31010 280120 31016
rect 280080 29782 280108 31010
rect 280816 30025 280844 57190
rect 282184 54528 282236 54534
rect 282184 54470 282236 54476
rect 280896 43444 280948 43450
rect 280896 43386 280948 43392
rect 280802 30016 280858 30025
rect 280908 29986 280936 43386
rect 280988 40724 281040 40730
rect 280988 40666 281040 40672
rect 280802 29951 280858 29960
rect 280896 29980 280948 29986
rect 280896 29922 280948 29928
rect 281000 29889 281028 40666
rect 281080 39364 281132 39370
rect 281080 39306 281132 39312
rect 281092 30054 281120 39306
rect 281172 36576 281224 36582
rect 281172 36518 281224 36524
rect 281080 30048 281132 30054
rect 281080 29990 281132 29996
rect 280986 29880 281042 29889
rect 280986 29815 281042 29824
rect 280068 29776 280120 29782
rect 280068 29718 280120 29724
rect 279976 29708 280028 29714
rect 279976 29650 280028 29656
rect 279424 29640 279476 29646
rect 279424 29582 279476 29588
rect 281184 28354 281212 36518
rect 281172 28348 281224 28354
rect 281172 28290 281224 28296
rect 282196 28218 282224 54470
rect 282828 51060 282880 51066
rect 282828 51002 282880 51008
rect 282840 50833 282868 51002
rect 282826 50824 282882 50833
rect 282826 50759 282882 50768
rect 282276 47592 282328 47598
rect 282276 47534 282328 47540
rect 282184 28212 282236 28218
rect 282184 28154 282236 28160
rect 282288 28150 282316 47534
rect 282276 28144 282328 28150
rect 282276 28086 282328 28092
rect 267004 28076 267056 28082
rect 267004 28018 267056 28024
rect 275928 28076 275980 28082
rect 275928 28018 275980 28024
rect 174544 28008 174596 28014
rect 174544 27950 174596 27956
rect 168932 27940 168984 27946
rect 168932 27882 168984 27888
rect 284956 6866 284984 193802
rect 286324 186992 286376 186998
rect 286324 186934 286376 186940
rect 286336 120086 286364 186934
rect 287072 125594 287100 200110
rect 292132 198121 292160 200110
rect 296180 198966 296208 200110
rect 299492 200110 299874 200138
rect 303632 200110 303922 200138
rect 307772 200110 307878 200138
rect 311926 200110 312032 200138
rect 296168 198960 296220 198966
rect 296168 198902 296220 198908
rect 292118 198112 292174 198121
rect 292118 198047 292174 198056
rect 289084 165640 289136 165646
rect 289084 165582 289136 165588
rect 287060 125588 287112 125594
rect 287060 125530 287112 125536
rect 286324 120080 286376 120086
rect 286324 120022 286376 120028
rect 289096 29170 289124 165582
rect 299492 148374 299520 200110
rect 303632 196994 303660 200110
rect 303620 196988 303672 196994
rect 303620 196930 303672 196936
rect 305644 177336 305696 177342
rect 305644 177278 305696 177284
rect 299480 148368 299532 148374
rect 299480 148310 299532 148316
rect 305656 135250 305684 177278
rect 305644 135244 305696 135250
rect 305644 135186 305696 135192
rect 289084 29164 289136 29170
rect 289084 29106 289136 29112
rect 307772 28354 307800 200110
rect 312004 198898 312032 200110
rect 315592 200110 315882 200138
rect 319640 200110 319930 200138
rect 323504 200110 323886 200138
rect 327552 200110 327934 200138
rect 331600 200110 331890 200138
rect 335372 200110 335938 200138
rect 339512 200110 339894 200138
rect 343850 200110 344232 200138
rect 311992 198892 312044 198898
rect 311992 198834 312044 198840
rect 315592 197062 315620 200110
rect 319640 198830 319668 200110
rect 319628 198824 319680 198830
rect 319628 198766 319680 198772
rect 323504 198490 323532 200110
rect 327552 199034 327580 200110
rect 327540 199028 327592 199034
rect 327540 198970 327592 198976
rect 323492 198484 323544 198490
rect 323492 198426 323544 198432
rect 323584 198076 323636 198082
rect 323584 198018 323636 198024
rect 319444 198008 319496 198014
rect 319444 197950 319496 197956
rect 315580 197056 315632 197062
rect 315580 196998 315632 197004
rect 309784 180124 309836 180130
rect 309784 180066 309836 180072
rect 309796 133890 309824 180066
rect 309784 133884 309836 133890
rect 309784 133826 309836 133832
rect 307760 28348 307812 28354
rect 307760 28290 307812 28296
rect 319456 28082 319484 197950
rect 323596 142866 323624 198018
rect 331600 197130 331628 200110
rect 331588 197124 331640 197130
rect 331588 197066 331640 197072
rect 323584 142860 323636 142866
rect 323584 142802 323636 142808
rect 335372 36582 335400 200110
rect 339512 198558 339540 200110
rect 344204 198830 344232 200110
rect 347792 200110 347898 200138
rect 351472 200110 351854 200138
rect 355520 200110 355902 200138
rect 359858 200110 360148 200138
rect 363906 200110 364288 200138
rect 367862 200110 368152 200138
rect 344192 198824 344244 198830
rect 344192 198766 344244 198772
rect 339500 198552 339552 198558
rect 339500 198494 339552 198500
rect 347792 129742 347820 200110
rect 351472 198626 351500 200110
rect 351460 198620 351512 198626
rect 351460 198562 351512 198568
rect 355520 197198 355548 200110
rect 360120 198393 360148 200110
rect 364260 198558 364288 200110
rect 368124 198626 368152 200110
rect 371252 200110 371910 200138
rect 375576 200110 375866 200138
rect 379624 200110 379914 200138
rect 383672 200110 383870 200138
rect 387812 200110 387918 200138
rect 391584 200110 391874 200138
rect 395632 200110 395922 200138
rect 399878 200110 400168 200138
rect 368112 198620 368164 198626
rect 368112 198562 368164 198568
rect 364248 198552 364300 198558
rect 364248 198494 364300 198500
rect 360106 198384 360162 198393
rect 360106 198319 360162 198328
rect 355508 197192 355560 197198
rect 355508 197134 355560 197140
rect 349804 178696 349856 178702
rect 349804 178638 349856 178644
rect 347780 129736 347832 129742
rect 347780 129678 347832 129684
rect 349816 124166 349844 178638
rect 371252 152522 371280 200110
rect 375576 197266 375604 200110
rect 379624 198694 379652 200110
rect 379612 198688 379664 198694
rect 379612 198630 379664 198636
rect 383672 197334 383700 200110
rect 387812 198529 387840 200110
rect 387798 198520 387854 198529
rect 387798 198455 387854 198464
rect 391584 198014 391612 200110
rect 393228 199504 393280 199510
rect 393228 199446 393280 199452
rect 391572 198008 391624 198014
rect 391572 197950 391624 197956
rect 383660 197328 383712 197334
rect 383660 197270 383712 197276
rect 375564 197260 375616 197266
rect 375564 197202 375616 197208
rect 392676 195696 392728 195702
rect 392676 195638 392728 195644
rect 392584 195628 392636 195634
rect 392584 195570 392636 195576
rect 389824 192568 389876 192574
rect 389824 192510 389876 192516
rect 387340 181076 387392 181082
rect 387340 181018 387392 181024
rect 387352 175234 387380 181018
rect 384304 175228 384356 175234
rect 384304 175170 384356 175176
rect 387340 175228 387392 175234
rect 387340 175170 387392 175176
rect 384316 168434 384344 175170
rect 382280 168428 382332 168434
rect 382280 168370 382332 168376
rect 384304 168428 384356 168434
rect 384304 168370 384356 168376
rect 382292 164830 382320 168370
rect 381544 164824 381596 164830
rect 381544 164766 381596 164772
rect 382280 164824 382332 164830
rect 382280 164766 382332 164772
rect 381556 154358 381584 164766
rect 379520 154352 379572 154358
rect 379520 154294 379572 154300
rect 381544 154352 381596 154358
rect 381544 154294 381596 154300
rect 371240 152516 371292 152522
rect 371240 152458 371292 152464
rect 379532 146334 379560 154294
rect 379520 146328 379572 146334
rect 379520 146270 379572 146276
rect 377312 146260 377364 146266
rect 377312 146202 377364 146208
rect 377324 142866 377352 146202
rect 376024 142860 376076 142866
rect 376024 142802 376076 142808
rect 377312 142860 377364 142866
rect 377312 142802 377364 142808
rect 376036 126682 376064 142802
rect 375012 126676 375064 126682
rect 375012 126618 375064 126624
rect 376024 126676 376076 126682
rect 376024 126618 376076 126624
rect 375024 124234 375052 126618
rect 372620 124228 372672 124234
rect 372620 124170 372672 124176
rect 375012 124228 375064 124234
rect 375012 124170 375064 124176
rect 349804 124160 349856 124166
rect 349804 124102 349856 124108
rect 372632 123146 372660 124170
rect 371884 123140 371936 123146
rect 371884 123082 371936 123088
rect 372620 123140 372672 123146
rect 372620 123082 372672 123088
rect 371896 98054 371924 123082
rect 371884 98048 371936 98054
rect 371884 97990 371936 97996
rect 367744 97980 367796 97986
rect 367744 97922 367796 97928
rect 367756 91118 367784 97922
rect 364984 91112 365036 91118
rect 364984 91054 365036 91060
rect 367744 91112 367796 91118
rect 367744 91054 367796 91060
rect 364996 84046 365024 91054
rect 360200 84040 360252 84046
rect 360200 83982 360252 83988
rect 364984 84040 365036 84046
rect 364984 83982 365036 83988
rect 360212 81462 360240 83982
rect 356704 81456 356756 81462
rect 356704 81398 356756 81404
rect 360200 81456 360252 81462
rect 360200 81398 360252 81404
rect 356716 68338 356744 81398
rect 355324 68332 355376 68338
rect 355324 68274 355376 68280
rect 356704 68332 356756 68338
rect 356704 68274 356756 68280
rect 355336 56642 355364 68274
rect 355324 56636 355376 56642
rect 355324 56578 355376 56584
rect 351920 56568 351972 56574
rect 351920 56510 351972 56516
rect 351932 53854 351960 56510
rect 347504 53848 347556 53854
rect 347504 53790 347556 53796
rect 351920 53848 351972 53854
rect 351920 53790 351972 53796
rect 347516 51066 347544 53790
rect 347504 51060 347556 51066
rect 347504 51002 347556 51008
rect 335360 36576 335412 36582
rect 335360 36518 335412 36524
rect 389836 28286 389864 192510
rect 390560 182912 390612 182918
rect 390560 182854 390612 182860
rect 390572 181082 390600 182854
rect 390560 181076 390612 181082
rect 390560 181018 390612 181024
rect 392596 140049 392624 195570
rect 392688 140282 392716 195638
rect 393136 195560 393188 195566
rect 393136 195502 393188 195508
rect 392952 195424 393004 195430
rect 392952 195366 393004 195372
rect 392768 192704 392820 192710
rect 392768 192646 392820 192652
rect 392676 140276 392728 140282
rect 392676 140218 392728 140224
rect 392582 140040 392638 140049
rect 392582 139975 392638 139984
rect 392596 92478 392624 139975
rect 392584 92472 392636 92478
rect 392584 92414 392636 92420
rect 392688 89690 392716 140218
rect 392780 139913 392808 192646
rect 392766 139904 392822 139913
rect 392766 139839 392822 139848
rect 392780 123486 392808 139839
rect 392768 123480 392820 123486
rect 392768 123422 392820 123428
rect 392676 89684 392728 89690
rect 392676 89626 392728 89632
rect 392964 82142 392992 195366
rect 393044 195356 393096 195362
rect 393044 195298 393096 195304
rect 392584 82136 392636 82142
rect 392584 82078 392636 82084
rect 392952 82136 393004 82142
rect 392952 82078 393004 82084
rect 391940 31544 391992 31550
rect 391940 31486 391992 31492
rect 391952 31074 391980 31486
rect 391940 31068 391992 31074
rect 391940 31010 391992 31016
rect 392596 30122 392624 82078
rect 393056 66910 393084 195298
rect 392676 66904 392728 66910
rect 392676 66846 392728 66852
rect 393044 66904 393096 66910
rect 393044 66846 393096 66852
rect 392584 30116 392636 30122
rect 392584 30058 392636 30064
rect 392688 28422 392716 66846
rect 393148 59265 393176 195502
rect 393134 59256 393190 59265
rect 393134 59191 393190 59200
rect 393240 31550 393268 199446
rect 395436 198144 395488 198150
rect 395436 198086 395488 198092
rect 394424 195832 394476 195838
rect 394424 195774 394476 195780
rect 394332 195492 394384 195498
rect 394332 195434 394384 195440
rect 393964 192636 394016 192642
rect 393964 192578 394016 192584
rect 393976 142154 394004 192578
rect 393884 142126 394004 142154
rect 393780 141024 393832 141030
rect 393780 140966 393832 140972
rect 393792 104854 393820 140966
rect 393884 140962 393912 142126
rect 394148 141704 394200 141710
rect 394148 141646 394200 141652
rect 393872 140956 393924 140962
rect 393872 140898 393924 140904
rect 393884 128382 393912 140898
rect 394160 140894 394188 141646
rect 394240 141568 394292 141574
rect 394240 141510 394292 141516
rect 394252 141030 394280 141510
rect 394240 141024 394292 141030
rect 394240 140966 394292 140972
rect 394148 140888 394200 140894
rect 394148 140830 394200 140836
rect 394160 140298 394188 140830
rect 394240 140616 394292 140622
rect 394240 140558 394292 140564
rect 394068 140270 394188 140298
rect 393872 128376 393924 128382
rect 393872 128318 393924 128324
rect 393780 104848 393832 104854
rect 393780 104790 393832 104796
rect 394068 102134 394096 140270
rect 394148 140208 394200 140214
rect 394148 140150 394200 140156
rect 394056 102128 394108 102134
rect 394056 102070 394108 102076
rect 394160 99346 394188 140150
rect 394148 99340 394200 99346
rect 394148 99282 394200 99288
rect 394252 95198 394280 140558
rect 394240 95192 394292 95198
rect 394240 95134 394292 95140
rect 394344 78606 394372 195434
rect 394332 78600 394384 78606
rect 394332 78542 394384 78548
rect 394344 64874 394372 78542
rect 393976 64846 394372 64874
rect 393228 31544 393280 31550
rect 393228 31486 393280 31492
rect 393976 30161 394004 64846
rect 394436 63481 394464 195774
rect 395250 195528 395306 195537
rect 395250 195463 395306 195472
rect 394608 192908 394660 192914
rect 394608 192850 394660 192856
rect 394516 192772 394568 192778
rect 394516 192714 394568 192720
rect 394422 63472 394478 63481
rect 394422 63407 394478 63416
rect 394528 40730 394556 192714
rect 394516 40724 394568 40730
rect 394516 40666 394568 40672
rect 394620 32434 394648 192850
rect 395160 139936 395212 139942
rect 395160 139878 395212 139884
rect 395172 106282 395200 139878
rect 395264 139777 395292 195463
rect 395344 184204 395396 184210
rect 395344 184146 395396 184152
rect 395250 139768 395306 139777
rect 395250 139703 395306 139712
rect 395160 106276 395212 106282
rect 395160 106218 395212 106224
rect 395264 85542 395292 139703
rect 395252 85536 395304 85542
rect 395252 85478 395304 85484
rect 394608 32428 394660 32434
rect 394608 32370 394660 32376
rect 393962 30152 394018 30161
rect 393962 30087 394018 30096
rect 395356 28694 395384 184146
rect 395448 140146 395476 198086
rect 395632 198082 395660 200110
rect 399576 199844 399628 199850
rect 399576 199786 399628 199792
rect 398380 199708 398432 199714
rect 398380 199650 398432 199656
rect 397368 198688 397420 198694
rect 397368 198630 397420 198636
rect 397276 198484 397328 198490
rect 397276 198426 397328 198432
rect 397184 198416 397236 198422
rect 397184 198358 397236 198364
rect 395804 198348 395856 198354
rect 395804 198290 395856 198296
rect 395712 198212 395764 198218
rect 395712 198154 395764 198160
rect 395620 198076 395672 198082
rect 395620 198018 395672 198024
rect 395528 198008 395580 198014
rect 395528 197950 395580 197956
rect 395436 140140 395488 140146
rect 395436 140082 395488 140088
rect 395448 97986 395476 140082
rect 395540 140078 395568 197950
rect 395620 197396 395672 197402
rect 395620 197338 395672 197344
rect 395528 140072 395580 140078
rect 395528 140014 395580 140020
rect 395436 97980 395488 97986
rect 395436 97922 395488 97928
rect 395540 86970 395568 140014
rect 395632 139942 395660 197338
rect 395620 139936 395672 139942
rect 395620 139878 395672 139884
rect 395620 118720 395672 118726
rect 395620 118662 395672 118668
rect 395632 91050 395660 118662
rect 395620 91044 395672 91050
rect 395620 90986 395672 90992
rect 395724 88330 395752 198154
rect 395816 197402 395844 198290
rect 395896 198280 395948 198286
rect 395896 198222 395948 198228
rect 395804 197396 395856 197402
rect 395804 197338 395856 197344
rect 395804 141500 395856 141506
rect 395804 141442 395856 141448
rect 395712 88324 395764 88330
rect 395712 88266 395764 88272
rect 395528 86964 395580 86970
rect 395528 86906 395580 86912
rect 395436 71868 395488 71874
rect 395436 71810 395488 71816
rect 395344 28688 395396 28694
rect 395344 28630 395396 28636
rect 395448 28490 395476 71810
rect 395816 28626 395844 141442
rect 395908 79694 395936 198222
rect 396724 198144 396776 198150
rect 396724 198086 396776 198092
rect 395988 195900 396040 195906
rect 395988 195842 396040 195848
rect 395896 79688 395948 79694
rect 395896 79630 395948 79636
rect 396000 57254 396028 195842
rect 396736 140078 396764 198086
rect 397000 195968 397052 195974
rect 397000 195910 397052 195916
rect 396908 195764 396960 195770
rect 396908 195706 396960 195712
rect 396080 140072 396132 140078
rect 396080 140014 396132 140020
rect 396724 140072 396776 140078
rect 396724 140014 396776 140020
rect 396092 139874 396120 140014
rect 396540 140004 396592 140010
rect 396540 139946 396592 139952
rect 396080 139868 396132 139874
rect 396080 139810 396132 139816
rect 396092 118726 396120 139810
rect 396080 118720 396132 118726
rect 396080 118662 396132 118668
rect 396552 113082 396580 139946
rect 396816 139936 396868 139942
rect 396816 139878 396868 139884
rect 396632 139596 396684 139602
rect 396632 139538 396684 139544
rect 396644 118658 396672 139538
rect 396828 139534 396856 139878
rect 396816 139528 396868 139534
rect 396816 139470 396868 139476
rect 396632 118652 396684 118658
rect 396632 118594 396684 118600
rect 396540 113076 396592 113082
rect 396540 113018 396592 113024
rect 396828 96529 396856 139470
rect 396814 96520 396870 96529
rect 396814 96455 396870 96464
rect 396920 75274 396948 195706
rect 396908 75268 396960 75274
rect 396908 75210 396960 75216
rect 396920 64874 396948 75210
rect 396736 64846 396948 64874
rect 395988 57248 396040 57254
rect 395988 57190 396040 57196
rect 395804 28620 395856 28626
rect 395804 28562 395856 28568
rect 396736 28558 396764 64846
rect 397012 54534 397040 195910
rect 397092 195220 397144 195226
rect 397092 195162 397144 195168
rect 397000 54528 397052 54534
rect 397000 54470 397052 54476
rect 397012 53961 397040 54470
rect 396998 53952 397054 53961
rect 396998 53887 397054 53896
rect 397104 49026 397132 195162
rect 397092 49020 397144 49026
rect 397092 48962 397144 48968
rect 397196 44033 397224 198358
rect 397182 44024 397238 44033
rect 397182 43959 397238 43968
rect 397196 43450 397224 43959
rect 397184 43444 397236 43450
rect 397184 43386 397236 43392
rect 397288 39370 397316 198426
rect 397276 39364 397328 39370
rect 397276 39306 397328 39312
rect 397380 34218 397408 198630
rect 397828 196852 397880 196858
rect 397828 196794 397880 196800
rect 397460 187740 397512 187746
rect 397460 187682 397512 187688
rect 397472 182918 397500 187682
rect 397460 182912 397512 182918
rect 397460 182854 397512 182860
rect 397840 135969 397868 196794
rect 397920 140752 397972 140758
rect 397920 140694 397972 140700
rect 397932 139505 397960 140694
rect 398196 140344 398248 140350
rect 398196 140286 398248 140292
rect 398012 140276 398064 140282
rect 398012 140218 398064 140224
rect 398024 139738 398052 140218
rect 398104 140140 398156 140146
rect 398104 140082 398156 140088
rect 398012 139732 398064 139738
rect 398012 139674 398064 139680
rect 397918 139496 397974 139505
rect 397918 139431 397974 139440
rect 398024 137442 398052 139674
rect 398116 139670 398144 140082
rect 398208 139806 398236 140286
rect 398288 140072 398340 140078
rect 398288 140014 398340 140020
rect 398196 139800 398248 139806
rect 398196 139742 398248 139748
rect 398104 139664 398156 139670
rect 398104 139606 398156 139612
rect 397932 137414 398052 137442
rect 397826 135960 397882 135969
rect 397826 135895 397882 135904
rect 397460 135244 397512 135250
rect 397460 135186 397512 135192
rect 397472 134337 397500 135186
rect 397458 134328 397514 134337
rect 397458 134263 397514 134272
rect 397460 133884 397512 133890
rect 397460 133826 397512 133832
rect 397472 132705 397500 133826
rect 397458 132696 397514 132705
rect 397458 132631 397514 132640
rect 397932 132494 397960 137414
rect 397840 132466 397960 132494
rect 397460 129736 397512 129742
rect 397460 129678 397512 129684
rect 397472 129441 397500 129678
rect 397458 129432 397514 129441
rect 397458 129367 397514 129376
rect 397460 125588 397512 125594
rect 397460 125530 397512 125536
rect 397472 124545 397500 125530
rect 397458 124536 397514 124545
rect 397458 124471 397514 124480
rect 397460 124160 397512 124166
rect 397460 124102 397512 124108
rect 397472 122913 397500 124102
rect 397458 122904 397514 122913
rect 397458 122839 397514 122848
rect 397460 120080 397512 120086
rect 397460 120022 397512 120028
rect 397472 119649 397500 120022
rect 397458 119640 397514 119649
rect 397458 119575 397514 119584
rect 397840 116249 397868 132466
rect 397920 123480 397972 123486
rect 397920 123422 397972 123428
rect 397826 116240 397882 116249
rect 397826 116175 397882 116184
rect 397932 113174 397960 123422
rect 398116 122834 398144 139606
rect 398024 122806 398144 122834
rect 398024 114617 398052 122806
rect 398104 118652 398156 118658
rect 398104 118594 398156 118600
rect 398116 117881 398144 118594
rect 398102 117872 398158 117881
rect 398102 117807 398158 117816
rect 398010 114608 398066 114617
rect 398010 114543 398066 114552
rect 397932 113146 398144 113174
rect 397552 113076 397604 113082
rect 397552 113018 397604 113024
rect 397564 112985 397592 113018
rect 397550 112976 397606 112985
rect 397550 112911 397606 112920
rect 397460 104848 397512 104854
rect 397458 104816 397460 104825
rect 397512 104816 397514 104825
rect 397458 104751 397514 104760
rect 397460 102128 397512 102134
rect 397460 102070 397512 102076
rect 397472 101561 397500 102070
rect 397458 101552 397514 101561
rect 397458 101487 397514 101496
rect 397460 99340 397512 99346
rect 397460 99282 397512 99288
rect 397472 98297 397500 99282
rect 397458 98288 397514 98297
rect 397458 98223 397514 98232
rect 397460 95192 397512 95198
rect 397460 95134 397512 95140
rect 397472 94897 397500 95134
rect 397458 94888 397514 94897
rect 397458 94823 397514 94832
rect 398116 93265 398144 113146
rect 398208 109721 398236 139742
rect 398194 109712 398250 109721
rect 398194 109647 398250 109656
rect 398196 97980 398248 97986
rect 398196 97922 398248 97928
rect 398102 93256 398158 93265
rect 398102 93191 398158 93200
rect 397460 92472 397512 92478
rect 397460 92414 397512 92420
rect 397472 91633 397500 92414
rect 397458 91624 397514 91633
rect 397458 91559 397514 91568
rect 397920 91044 397972 91050
rect 397920 90986 397972 90992
rect 397932 90001 397960 90986
rect 397918 89992 397974 90001
rect 397918 89927 397974 89936
rect 397460 89684 397512 89690
rect 397460 89626 397512 89632
rect 397472 88369 397500 89626
rect 397458 88360 397514 88369
rect 397458 88295 397514 88304
rect 397736 86964 397788 86970
rect 397736 86906 397788 86912
rect 397748 86737 397776 86906
rect 397734 86728 397790 86737
rect 397734 86663 397790 86672
rect 397552 85536 397604 85542
rect 397552 85478 397604 85484
rect 397564 85105 397592 85478
rect 397550 85096 397606 85105
rect 397550 85031 397606 85040
rect 397460 82136 397512 82142
rect 397460 82078 397512 82084
rect 397472 81841 397500 82078
rect 397458 81832 397514 81841
rect 397458 81767 397514 81776
rect 398208 80209 398236 97922
rect 398194 80200 398250 80209
rect 398194 80135 398250 80144
rect 398196 79688 398248 79694
rect 398196 79630 398248 79636
rect 397460 78600 397512 78606
rect 397458 78568 397460 78577
rect 397512 78568 397514 78577
rect 397458 78503 397514 78512
rect 398010 76936 398066 76945
rect 398010 76871 398066 76880
rect 398024 74534 398052 76871
rect 398102 75304 398158 75313
rect 398102 75239 398104 75248
rect 398156 75239 398158 75248
rect 398104 75210 398156 75216
rect 398024 74506 398144 74534
rect 397918 71904 397974 71913
rect 397918 71839 397920 71848
rect 397972 71839 397974 71848
rect 397920 71810 397972 71816
rect 397458 67008 397514 67017
rect 397458 66943 397514 66952
rect 397472 66910 397500 66943
rect 397460 66904 397512 66910
rect 397460 66846 397512 66852
rect 397458 60480 397514 60489
rect 397458 60415 397514 60424
rect 397472 59265 397500 60415
rect 397458 59256 397514 59265
rect 397458 59191 397514 59200
rect 397460 57248 397512 57254
rect 397458 57216 397460 57225
rect 397512 57216 397514 57225
rect 397458 57151 397514 57160
rect 398012 56228 398064 56234
rect 398012 56170 398064 56176
rect 397918 50552 397974 50561
rect 397918 50487 397974 50496
rect 397460 49020 397512 49026
rect 397460 48962 397512 48968
rect 397472 48929 397500 48962
rect 397458 48920 397514 48929
rect 397458 48855 397514 48864
rect 397460 47592 397512 47598
rect 397460 47534 397512 47540
rect 397472 47297 397500 47534
rect 397458 47288 397514 47297
rect 397458 47223 397514 47232
rect 397458 42392 397514 42401
rect 397458 42327 397514 42336
rect 397472 41478 397500 42327
rect 397460 41472 397512 41478
rect 397460 41414 397512 41420
rect 397458 40760 397514 40769
rect 397458 40695 397460 40704
rect 397512 40695 397514 40704
rect 397736 40724 397788 40730
rect 397460 40666 397512 40672
rect 397736 40666 397788 40672
rect 397460 39364 397512 39370
rect 397460 39306 397512 39312
rect 397472 39137 397500 39306
rect 397458 39128 397514 39137
rect 397458 39063 397514 39072
rect 397550 37496 397606 37505
rect 397550 37431 397606 37440
rect 397564 37330 397592 37431
rect 397552 37324 397604 37330
rect 397552 37266 397604 37272
rect 397458 34232 397514 34241
rect 397380 34190 397458 34218
rect 397380 33153 397408 34190
rect 397458 34167 397514 34176
rect 397366 33144 397422 33153
rect 397366 33079 397422 33088
rect 397458 32600 397514 32609
rect 397458 32535 397514 32544
rect 397472 32434 397500 32535
rect 397460 32428 397512 32434
rect 397460 32370 397512 32376
rect 397460 31544 397512 31550
rect 397460 31486 397512 31492
rect 397472 30977 397500 31486
rect 397458 30968 397514 30977
rect 397458 30903 397514 30912
rect 397748 30258 397776 40666
rect 397736 30252 397788 30258
rect 397736 30194 397788 30200
rect 397932 30190 397960 50487
rect 397920 30184 397972 30190
rect 397920 30126 397972 30132
rect 396724 28552 396776 28558
rect 396724 28494 396776 28500
rect 395436 28484 395488 28490
rect 395436 28426 395488 28432
rect 392676 28416 392728 28422
rect 392676 28358 392728 28364
rect 389824 28280 389876 28286
rect 389824 28222 389876 28228
rect 319444 28076 319496 28082
rect 319444 28018 319496 28024
rect 398024 27946 398052 56170
rect 398116 30326 398144 74506
rect 398208 73545 398236 79630
rect 398194 73536 398250 73545
rect 398194 73471 398250 73480
rect 398104 30320 398156 30326
rect 398104 30262 398156 30268
rect 398208 28898 398236 73471
rect 398300 71913 398328 140014
rect 398392 131073 398420 199650
rect 399208 199640 399260 199646
rect 399208 199582 399260 199588
rect 398930 199472 398986 199481
rect 398930 199407 398986 199416
rect 398748 196784 398800 196790
rect 398748 196726 398800 196732
rect 398472 144288 398524 144294
rect 398472 144230 398524 144236
rect 398378 131064 398434 131073
rect 398378 130999 398434 131008
rect 398380 128376 398432 128382
rect 398380 128318 398432 128324
rect 398392 99929 398420 128318
rect 398378 99920 398434 99929
rect 398378 99855 398434 99864
rect 398286 71904 398342 71913
rect 398286 71839 398342 71848
rect 398286 70272 398342 70281
rect 398286 70207 398342 70216
rect 398196 28892 398248 28898
rect 398196 28834 398248 28840
rect 398300 28762 398328 70207
rect 398378 68640 398434 68649
rect 398378 68575 398434 68584
rect 398392 28966 398420 68575
rect 398484 65385 398512 144230
rect 398564 142928 398616 142934
rect 398564 142870 398616 142876
rect 398470 65376 398526 65385
rect 398470 65311 398526 65320
rect 398484 31754 398512 65311
rect 398576 58857 398604 142870
rect 398656 141772 398708 141778
rect 398656 141714 398708 141720
rect 398562 58848 398618 58857
rect 398562 58783 398618 58792
rect 398472 31748 398524 31754
rect 398472 31690 398524 31696
rect 398576 31618 398604 58783
rect 398668 52193 398696 141714
rect 398654 52184 398710 52193
rect 398654 52119 398710 52128
rect 398668 31686 398696 52119
rect 398760 47297 398788 196726
rect 398840 139800 398892 139806
rect 398840 139742 398892 139748
rect 398852 139466 398880 139742
rect 398840 139460 398892 139466
rect 398840 139402 398892 139408
rect 398852 111353 398880 139402
rect 398838 111344 398894 111353
rect 398838 111279 398894 111288
rect 398840 88324 398892 88330
rect 398840 88266 398892 88272
rect 398852 76945 398880 88266
rect 398838 76936 398894 76945
rect 398838 76871 398894 76880
rect 398746 47288 398802 47297
rect 398746 47223 398802 47232
rect 398748 46912 398800 46918
rect 398748 46854 398800 46860
rect 398760 45665 398788 46854
rect 398746 45656 398802 45665
rect 398746 45591 398802 45600
rect 398760 40730 398788 45591
rect 398944 45554 398972 199407
rect 399116 196716 399168 196722
rect 399116 196658 399168 196664
rect 399024 196648 399076 196654
rect 399024 196590 399076 196596
rect 399036 46918 399064 196590
rect 399128 56234 399156 196658
rect 399220 68649 399248 199582
rect 399482 144120 399538 144129
rect 399482 144055 399538 144064
rect 399392 142860 399444 142866
rect 399392 142802 399444 142808
rect 399300 141636 399352 141642
rect 399300 141578 399352 141584
rect 399206 68640 399262 68649
rect 399206 68575 399262 68584
rect 399206 62112 399262 62121
rect 399206 62047 399262 62056
rect 399116 56228 399168 56234
rect 399116 56170 399168 56176
rect 399128 55593 399156 56170
rect 399114 55584 399170 55593
rect 399114 55519 399170 55528
rect 399024 46912 399076 46918
rect 399024 46854 399076 46860
rect 398852 45526 398972 45554
rect 398852 42401 398880 45526
rect 398838 42392 398894 42401
rect 398838 42327 398894 42336
rect 398748 40724 398800 40730
rect 398748 40666 398800 40672
rect 398656 31680 398708 31686
rect 398656 31622 398708 31628
rect 398564 31612 398616 31618
rect 398564 31554 398616 31560
rect 398380 28960 398432 28966
rect 398380 28902 398432 28908
rect 399220 28830 399248 62047
rect 399312 37505 399340 141578
rect 399404 50561 399432 142802
rect 399496 62121 399524 144055
rect 399588 127809 399616 199786
rect 399760 197872 399812 197878
rect 399760 197814 399812 197820
rect 399574 127800 399630 127809
rect 399574 127735 399630 127744
rect 399576 106276 399628 106282
rect 399576 106218 399628 106224
rect 399588 83473 399616 106218
rect 399574 83464 399630 83473
rect 399574 83399 399630 83408
rect 399482 62112 399538 62121
rect 399482 62047 399538 62056
rect 399390 50552 399446 50561
rect 399390 50487 399446 50496
rect 399298 37496 399354 37505
rect 399298 37431 399354 37440
rect 399772 35873 399800 197814
rect 400140 195294 400168 200110
rect 403544 200110 403926 200138
rect 407132 200110 407882 200138
rect 401048 200048 401100 200054
rect 401048 199990 401100 199996
rect 400956 199912 401008 199918
rect 400956 199854 401008 199860
rect 400864 197804 400916 197810
rect 400864 197746 400916 197752
rect 400128 195288 400180 195294
rect 400128 195230 400180 195236
rect 400680 191888 400732 191894
rect 400680 191830 400732 191836
rect 400692 187746 400720 191830
rect 400680 187740 400732 187746
rect 400680 187682 400732 187688
rect 400126 142760 400182 142769
rect 400126 142695 400182 142704
rect 400140 139806 400168 142695
rect 400220 140820 400272 140826
rect 400220 140762 400272 140768
rect 400128 139800 400180 139806
rect 400128 139742 400180 139748
rect 400232 103329 400260 140762
rect 400588 137896 400640 137902
rect 400588 137838 400640 137844
rect 400600 126721 400628 137838
rect 400586 126712 400642 126721
rect 400586 126647 400642 126656
rect 400588 121440 400640 121446
rect 400586 121408 400588 121417
rect 400640 121408 400642 121417
rect 400586 121343 400642 121352
rect 400218 103320 400274 103329
rect 400218 103255 400274 103264
rect 400876 74534 400904 197746
rect 400968 121446 400996 199854
rect 401060 137902 401088 199990
rect 403544 198665 403572 200110
rect 405004 199980 405056 199986
rect 405004 199922 405056 199928
rect 403530 198656 403586 198665
rect 403530 198591 403586 198600
rect 403624 197940 403676 197946
rect 403624 197882 403676 197888
rect 401232 192976 401284 192982
rect 401232 192918 401284 192924
rect 401140 192840 401192 192846
rect 401140 192782 401192 192788
rect 401152 139602 401180 192782
rect 401244 140826 401272 192918
rect 401232 140820 401284 140826
rect 401232 140762 401284 140768
rect 403636 140622 403664 197882
rect 404358 196072 404414 196081
rect 404358 196007 404414 196016
rect 403808 195152 403860 195158
rect 403808 195094 403860 195100
rect 403716 195084 403768 195090
rect 403716 195026 403768 195032
rect 403624 140616 403676 140622
rect 403624 140558 403676 140564
rect 403728 139942 403756 195026
rect 403820 140010 403848 195094
rect 404372 193338 404400 196007
rect 404280 193310 404400 193338
rect 404280 191894 404308 193310
rect 404268 191888 404320 191894
rect 404268 191830 404320 191836
rect 405016 141710 405044 199922
rect 406384 199572 406436 199578
rect 406384 199514 406436 199520
rect 406016 147008 406068 147014
rect 406016 146950 406068 146956
rect 406028 143478 406056 146950
rect 406016 143472 406068 143478
rect 406016 143414 406068 143420
rect 405004 141704 405056 141710
rect 405004 141646 405056 141652
rect 403808 140004 403860 140010
rect 403808 139946 403860 139952
rect 403716 139936 403768 139942
rect 403716 139878 403768 139884
rect 406028 139890 406056 143414
rect 406396 141574 406424 199514
rect 407132 188358 407160 200110
rect 407764 199776 407816 199782
rect 407764 199718 407816 199724
rect 407120 188352 407172 188358
rect 407120 188294 407172 188300
rect 406384 141568 406436 141574
rect 406384 141510 406436 141516
rect 407776 140214 407804 199718
rect 409248 196625 409276 410230
rect 409326 410207 409382 410216
rect 409326 404424 409382 404433
rect 409326 404359 409382 404368
rect 409340 196858 409368 404359
rect 409432 398857 409460 436766
rect 409418 398848 409474 398857
rect 409418 398783 409474 398792
rect 409892 355881 409920 486406
rect 410536 457502 410564 497014
rect 415398 496904 415454 496913
rect 415398 496839 415454 496848
rect 416778 496904 416834 496913
rect 416778 496839 416834 496848
rect 418158 496904 418214 496913
rect 418158 496839 418214 496848
rect 419538 496904 419594 496913
rect 419538 496839 419594 496848
rect 415412 496126 415440 496839
rect 415400 496120 415452 496126
rect 415400 496062 415452 496068
rect 410524 457496 410576 457502
rect 410524 457438 410576 457444
rect 410708 451920 410760 451926
rect 410708 451862 410760 451868
rect 410616 449200 410668 449206
rect 410616 449142 410668 449148
rect 410432 446412 410484 446418
rect 410432 446354 410484 446360
rect 410156 439544 410208 439550
rect 410156 439486 410208 439492
rect 409972 429888 410024 429894
rect 409972 429830 410024 429836
rect 409878 355872 409934 355881
rect 409878 355807 409934 355816
rect 409984 320929 410012 429830
rect 410064 428528 410116 428534
rect 410064 428470 410116 428476
rect 410076 333169 410104 428470
rect 410168 363497 410196 439486
rect 410248 431316 410300 431322
rect 410248 431258 410300 431264
rect 410260 369617 410288 431258
rect 410340 423292 410392 423298
rect 410340 423234 410392 423240
rect 410246 369608 410302 369617
rect 410246 369543 410302 369552
rect 410154 363488 410210 363497
rect 410154 363423 410210 363432
rect 410062 333160 410118 333169
rect 410062 333095 410118 333104
rect 409970 320920 410026 320929
rect 409970 320855 410026 320864
rect 409878 307728 409934 307737
rect 409878 307663 409934 307672
rect 409420 237380 409472 237386
rect 409420 237322 409472 237328
rect 409432 236201 409460 237322
rect 409418 236192 409474 236201
rect 409418 236127 409474 236136
rect 409328 196852 409380 196858
rect 409328 196794 409380 196800
rect 409234 196616 409290 196625
rect 409234 196551 409290 196560
rect 409432 142934 409460 236127
rect 409510 227896 409566 227905
rect 409510 227831 409566 227840
rect 409524 227798 409552 227831
rect 409512 227792 409564 227798
rect 409512 227734 409564 227740
rect 409420 142928 409472 142934
rect 409420 142870 409472 142876
rect 409524 141778 409552 227734
rect 409512 141772 409564 141778
rect 409512 141714 409564 141720
rect 409892 140282 409920 307663
rect 409972 306332 410024 306338
rect 409972 306274 410024 306280
rect 409984 305425 410012 306274
rect 409970 305416 410026 305425
rect 409970 305351 410026 305360
rect 409880 140276 409932 140282
rect 409880 140218 409932 140224
rect 407764 140208 407816 140214
rect 407764 140150 407816 140156
rect 409984 140146 410012 305351
rect 410154 299704 410210 299713
rect 410076 299662 410154 299690
rect 410076 140350 410104 299662
rect 410154 299639 410210 299648
rect 410156 296676 410208 296682
rect 410156 296618 410208 296624
rect 410168 295633 410196 296618
rect 410154 295624 410210 295633
rect 410154 295559 410210 295568
rect 410168 140758 410196 295559
rect 410246 252512 410302 252521
rect 410246 252447 410302 252456
rect 410156 140752 410208 140758
rect 410156 140694 410208 140700
rect 410064 140344 410116 140350
rect 410064 140286 410116 140292
rect 409972 140140 410024 140146
rect 409972 140082 410024 140088
rect 410260 140078 410288 252447
rect 410352 225049 410380 423234
rect 410444 394369 410472 446354
rect 410524 432676 410576 432682
rect 410524 432618 410576 432624
rect 410430 394360 410486 394369
rect 410430 394295 410486 394304
rect 410430 392320 410486 392329
rect 410430 392255 410486 392264
rect 410338 225040 410394 225049
rect 410338 224975 410394 224984
rect 410338 221640 410394 221649
rect 410338 221575 410394 221584
rect 410352 196790 410380 221575
rect 410444 199714 410472 392255
rect 410536 373833 410564 432618
rect 410628 400489 410656 449142
rect 410720 414905 410748 451862
rect 411996 447840 412048 447846
rect 411996 447782 412048 447788
rect 411904 443692 411956 443698
rect 411904 443634 411956 443640
rect 411812 442264 411864 442270
rect 411812 442206 411864 442212
rect 411720 436756 411772 436762
rect 411720 436698 411772 436704
rect 411260 435396 411312 435402
rect 411260 435338 411312 435344
rect 410706 414896 410762 414905
rect 410706 414831 410762 414840
rect 410614 400480 410670 400489
rect 410614 400415 410670 400424
rect 410522 373824 410578 373833
rect 410522 373759 410578 373768
rect 411272 371906 411300 435338
rect 411352 432608 411404 432614
rect 411352 432550 411404 432556
rect 411180 371878 411300 371906
rect 411180 371090 411208 371878
rect 411258 371784 411314 371793
rect 411258 371719 411314 371728
rect 411272 371278 411300 371719
rect 411260 371272 411312 371278
rect 411260 371214 411312 371220
rect 411180 371062 411300 371090
rect 411272 365537 411300 371062
rect 411258 365528 411314 365537
rect 411258 365463 411314 365472
rect 411258 359408 411314 359417
rect 411258 359343 411260 359352
rect 411312 359343 411314 359352
rect 411260 359314 411312 359320
rect 411364 357377 411392 432550
rect 411628 431248 411680 431254
rect 411628 431190 411680 431196
rect 411444 429956 411496 429962
rect 411444 429898 411496 429904
rect 411350 357368 411406 357377
rect 411350 357303 411406 357312
rect 411260 353184 411312 353190
rect 411258 353152 411260 353161
rect 411312 353152 411314 353161
rect 411258 353087 411314 353096
rect 410614 349072 410670 349081
rect 410614 349007 410670 349016
rect 410524 309120 410576 309126
rect 410524 309062 410576 309068
rect 410536 308009 410564 309062
rect 410522 308000 410578 308009
rect 410522 307935 410578 307944
rect 410524 300824 410576 300830
rect 410524 300766 410576 300772
rect 410536 299713 410564 300766
rect 410522 299704 410578 299713
rect 410522 299639 410578 299648
rect 410522 244216 410578 244225
rect 410522 244151 410578 244160
rect 410432 199708 410484 199714
rect 410432 199650 410484 199656
rect 410340 196784 410392 196790
rect 410340 196726 410392 196732
rect 410536 144294 410564 244151
rect 410628 193905 410656 349007
rect 411456 347041 411484 429898
rect 411536 428460 411588 428466
rect 411536 428402 411588 428408
rect 411442 347032 411498 347041
rect 411442 346967 411498 346976
rect 411258 344992 411314 345001
rect 411258 344927 411314 344936
rect 411272 343738 411300 344927
rect 411260 343732 411312 343738
rect 411260 343674 411312 343680
rect 411258 342952 411314 342961
rect 411258 342887 411314 342896
rect 411272 342310 411300 342887
rect 411260 342304 411312 342310
rect 411260 342246 411312 342252
rect 411442 340912 411498 340921
rect 411442 340847 411498 340856
rect 410706 338872 410762 338881
rect 410706 338807 410762 338816
rect 410720 194041 410748 338807
rect 411260 338088 411312 338094
rect 411260 338030 411312 338036
rect 411272 336841 411300 338030
rect 411258 336832 411314 336841
rect 411258 336767 411314 336776
rect 411258 330576 411314 330585
rect 411258 330511 411314 330520
rect 411272 329866 411300 330511
rect 411260 329860 411312 329866
rect 411260 329802 411312 329808
rect 411258 326496 411314 326505
rect 411258 326431 411314 326440
rect 411272 325718 411300 326431
rect 411260 325712 411312 325718
rect 411260 325654 411312 325660
rect 411258 324456 411314 324465
rect 411258 324391 411314 324400
rect 411272 324358 411300 324391
rect 411260 324352 411312 324358
rect 411260 324294 411312 324300
rect 411258 318200 411314 318209
rect 411258 318135 411314 318144
rect 411272 317490 411300 318135
rect 411260 317484 411312 317490
rect 411260 317426 411312 317432
rect 411258 316160 411314 316169
rect 411258 316095 411314 316104
rect 411272 316062 411300 316095
rect 411260 316056 411312 316062
rect 411260 315998 411312 316004
rect 411258 314120 411314 314129
rect 411258 314055 411314 314064
rect 411272 313342 411300 314055
rect 411260 313336 411312 313342
rect 411260 313278 411312 313284
rect 411258 312080 411314 312089
rect 411258 312015 411314 312024
rect 411272 311914 411300 312015
rect 411260 311908 411312 311914
rect 411260 311850 411312 311856
rect 411258 310040 411314 310049
rect 411258 309975 411314 309984
rect 411272 309194 411300 309975
rect 411260 309188 411312 309194
rect 411260 309130 411312 309136
rect 411258 303920 411314 303929
rect 411258 303855 411314 303864
rect 411272 303686 411300 303855
rect 411260 303680 411312 303686
rect 411260 303622 411312 303628
rect 411260 297968 411312 297974
rect 411260 297910 411312 297916
rect 411272 297673 411300 297910
rect 411258 297664 411314 297673
rect 411258 297599 411314 297608
rect 411258 293584 411314 293593
rect 411258 293519 411314 293528
rect 411272 292602 411300 293519
rect 411260 292596 411312 292602
rect 411260 292538 411312 292544
rect 411258 291544 411314 291553
rect 411258 291479 411314 291488
rect 411272 291242 411300 291479
rect 411260 291236 411312 291242
rect 411260 291178 411312 291184
rect 411258 289504 411314 289513
rect 411258 289439 411314 289448
rect 411272 288454 411300 289439
rect 411260 288448 411312 288454
rect 411260 288390 411312 288396
rect 411258 287464 411314 287473
rect 411258 287399 411314 287408
rect 411272 287094 411300 287399
rect 411260 287088 411312 287094
rect 411260 287030 411312 287036
rect 411258 285288 411314 285297
rect 411258 285223 411314 285232
rect 411272 284374 411300 285223
rect 411260 284368 411312 284374
rect 411260 284310 411312 284316
rect 411258 283248 411314 283257
rect 411258 283183 411314 283192
rect 411272 282946 411300 283183
rect 411260 282940 411312 282946
rect 411260 282882 411312 282888
rect 411258 281208 411314 281217
rect 411258 281143 411314 281152
rect 411272 280226 411300 281143
rect 411260 280220 411312 280226
rect 411260 280162 411312 280168
rect 411260 279472 411312 279478
rect 411260 279414 411312 279420
rect 411272 279177 411300 279414
rect 411258 279168 411314 279177
rect 411258 279103 411314 279112
rect 411258 277128 411314 277137
rect 411258 277063 411314 277072
rect 411272 276894 411300 277063
rect 411260 276888 411312 276894
rect 411260 276830 411312 276836
rect 411258 275088 411314 275097
rect 411258 275023 411314 275032
rect 411272 274718 411300 275023
rect 411260 274712 411312 274718
rect 411260 274654 411312 274660
rect 411260 273216 411312 273222
rect 411260 273158 411312 273164
rect 411272 273057 411300 273158
rect 411258 273048 411314 273057
rect 411258 272983 411314 272992
rect 411258 271008 411314 271017
rect 411258 270943 411314 270952
rect 411272 270570 411300 270943
rect 411260 270564 411312 270570
rect 411260 270506 411312 270512
rect 411258 268968 411314 268977
rect 411258 268903 411314 268912
rect 411272 267782 411300 268903
rect 411260 267776 411312 267782
rect 411260 267718 411312 267724
rect 411260 267028 411312 267034
rect 411260 266970 411312 266976
rect 411272 266801 411300 266970
rect 411258 266792 411314 266801
rect 411258 266727 411314 266736
rect 411258 264752 411314 264761
rect 411258 264687 411314 264696
rect 411272 263634 411300 264687
rect 411260 263628 411312 263634
rect 411260 263570 411312 263576
rect 411260 262880 411312 262886
rect 411260 262822 411312 262828
rect 411272 262721 411300 262822
rect 411258 262712 411314 262721
rect 411258 262647 411314 262656
rect 411258 260672 411314 260681
rect 411258 260607 411314 260616
rect 411272 259486 411300 260607
rect 411260 259480 411312 259486
rect 411260 259422 411312 259428
rect 411260 258732 411312 258738
rect 411260 258674 411312 258680
rect 411272 258641 411300 258674
rect 411258 258632 411314 258641
rect 411258 258567 411314 258576
rect 411258 256592 411314 256601
rect 411258 256527 411314 256536
rect 411272 255338 411300 256527
rect 411260 255332 411312 255338
rect 411260 255274 411312 255280
rect 411260 254584 411312 254590
rect 411258 254552 411260 254561
rect 411312 254552 411314 254561
rect 411258 254487 411314 254496
rect 410800 252544 410852 252550
rect 410798 252512 410800 252521
rect 410852 252512 410854 252521
rect 410798 252447 410854 252456
rect 411260 250504 411312 250510
rect 411260 250446 411312 250452
rect 411272 250345 411300 250446
rect 411258 250336 411314 250345
rect 411258 250271 411314 250280
rect 411258 246256 411314 246265
rect 411258 246191 411314 246200
rect 411272 245682 411300 246191
rect 411260 245676 411312 245682
rect 411260 245618 411312 245624
rect 410800 244248 410852 244254
rect 410798 244216 410800 244225
rect 410852 244216 410854 244225
rect 410798 244151 410854 244160
rect 411258 242176 411314 242185
rect 411258 242111 411314 242120
rect 411272 241874 411300 242111
rect 411260 241868 411312 241874
rect 411260 241810 411312 241816
rect 411258 240136 411314 240145
rect 411258 240071 411260 240080
rect 411312 240071 411314 240080
rect 411260 240042 411312 240048
rect 411258 238096 411314 238105
rect 411258 238031 411314 238040
rect 411272 237454 411300 238031
rect 411260 237448 411312 237454
rect 411260 237390 411312 237396
rect 411258 233880 411314 233889
rect 411258 233815 411314 233824
rect 411272 233306 411300 233815
rect 411260 233300 411312 233306
rect 411260 233242 411312 233248
rect 411350 231840 411406 231849
rect 411350 231775 411406 231784
rect 411364 231130 411392 231775
rect 411352 231124 411404 231130
rect 411352 231066 411404 231072
rect 411258 229800 411314 229809
rect 411258 229735 411314 229744
rect 411272 229158 411300 229735
rect 411260 229152 411312 229158
rect 411260 229094 411312 229100
rect 411258 223680 411314 223689
rect 411258 223615 411260 223624
rect 411312 223615 411314 223624
rect 411260 223586 411312 223592
rect 410800 222148 410852 222154
rect 410800 222090 410852 222096
rect 410812 221649 410840 222090
rect 410798 221640 410854 221649
rect 410798 221575 410854 221584
rect 411258 217424 411314 217433
rect 411258 217359 411314 217368
rect 411272 217326 411300 217359
rect 411260 217320 411312 217326
rect 411260 217262 411312 217268
rect 411260 213376 411312 213382
rect 411258 213344 411260 213353
rect 411312 213344 411314 213353
rect 411258 213279 411314 213288
rect 411260 211812 411312 211818
rect 411260 211754 411312 211760
rect 411272 211313 411300 211754
rect 411258 211304 411314 211313
rect 411258 211239 411314 211248
rect 411352 207664 411404 207670
rect 411352 207606 411404 207612
rect 411364 207233 411392 207606
rect 411350 207224 411406 207233
rect 411350 207159 411406 207168
rect 411258 205184 411314 205193
rect 411258 205119 411314 205128
rect 411272 204338 411300 205119
rect 411260 204332 411312 204338
rect 411260 204274 411312 204280
rect 411258 203144 411314 203153
rect 411258 203079 411260 203088
rect 411312 203079 411314 203088
rect 411260 203050 411312 203056
rect 411258 201104 411314 201113
rect 411258 201039 411314 201048
rect 411272 200802 411300 201039
rect 411260 200796 411312 200802
rect 411260 200738 411312 200744
rect 411272 199510 411300 200738
rect 411260 199504 411312 199510
rect 411260 199446 411312 199452
rect 411364 197878 411392 207159
rect 411456 199918 411484 340847
rect 411548 322425 411576 428402
rect 411640 351121 411668 431190
rect 411732 382106 411760 436698
rect 411824 386073 411852 442206
rect 411916 388249 411944 443634
rect 412008 396409 412036 447782
rect 416792 428602 416820 496839
rect 416780 428596 416832 428602
rect 416780 428538 416832 428544
rect 418172 425746 418200 496839
rect 419552 487830 419580 496839
rect 419644 490618 419672 498063
rect 432142 497176 432198 497185
rect 432142 497111 432198 497120
rect 432156 497078 432184 497111
rect 432144 497072 432196 497078
rect 426438 497040 426494 497049
rect 426438 496975 426494 496984
rect 427910 497040 427966 497049
rect 427910 496975 427966 496984
rect 430578 497040 430634 497049
rect 432144 497014 432196 497020
rect 433430 497040 433486 497049
rect 430578 496975 430634 496984
rect 432604 497004 432656 497010
rect 426452 496942 426480 496975
rect 426440 496936 426492 496942
rect 420918 496904 420974 496913
rect 420918 496839 420974 496848
rect 422298 496904 422354 496913
rect 422298 496839 422354 496848
rect 423678 496904 423734 496913
rect 425058 496904 425114 496913
rect 423678 496839 423734 496848
rect 424324 496868 424376 496874
rect 419632 490612 419684 490618
rect 419632 490554 419684 490560
rect 419540 487824 419592 487830
rect 419540 487766 419592 487772
rect 420932 426154 420960 496839
rect 422312 486538 422340 496839
rect 422300 486532 422352 486538
rect 422300 486474 422352 486480
rect 423692 480962 423720 496839
rect 427084 496936 427136 496942
rect 426440 496878 426492 496884
rect 426530 496904 426586 496913
rect 425058 496839 425114 496848
rect 427084 496878 427136 496884
rect 427818 496904 427874 496913
rect 426530 496839 426532 496848
rect 424324 496810 424376 496816
rect 423680 480956 423732 480962
rect 423680 480898 423732 480904
rect 424336 453354 424364 496810
rect 425072 471306 425100 496839
rect 426584 496839 426586 496848
rect 426532 496810 426584 496816
rect 425060 471300 425112 471306
rect 425060 471242 425112 471248
rect 424324 453348 424376 453354
rect 424324 453290 424376 453296
rect 420920 426148 420972 426154
rect 420920 426090 420972 426096
rect 418160 425740 418212 425746
rect 418160 425682 418212 425688
rect 427096 423162 427124 496878
rect 427818 496839 427874 496848
rect 427832 467158 427860 496839
rect 427924 491978 427952 496975
rect 430592 496942 430620 496975
rect 433430 496975 433486 496984
rect 432604 496946 432656 496952
rect 430580 496936 430632 496942
rect 429198 496904 429254 496913
rect 428464 496868 428516 496874
rect 430580 496878 430632 496884
rect 430670 496904 430726 496913
rect 429198 496839 429254 496848
rect 430670 496839 430726 496848
rect 428464 496810 428516 496816
rect 427912 491972 427964 491978
rect 427912 491914 427964 491920
rect 427820 467152 427872 467158
rect 427820 467094 427872 467100
rect 428476 423230 428504 496810
rect 429212 454714 429240 496839
rect 429200 454708 429252 454714
rect 429200 454650 429252 454656
rect 430684 424386 430712 496839
rect 432616 450634 432644 496946
rect 433338 496904 433394 496913
rect 433338 496839 433340 496848
rect 433392 496839 433394 496848
rect 433340 496810 433392 496816
rect 433444 493338 433472 496975
rect 433432 493332 433484 493338
rect 433432 493274 433484 493280
rect 433536 485178 433564 498063
rect 434718 497040 434774 497049
rect 434718 496975 434774 496984
rect 437478 497040 437534 497049
rect 437478 496975 437534 496984
rect 433524 485172 433576 485178
rect 433524 485114 433576 485120
rect 432604 450628 432656 450634
rect 432604 450570 432656 450576
rect 434732 426290 434760 496975
rect 434810 496904 434866 496913
rect 434810 496839 434866 496848
rect 436098 496904 436154 496913
rect 436098 496839 436154 496848
rect 434824 489190 434852 496839
rect 434812 489184 434864 489190
rect 434812 489126 434864 489132
rect 436112 427174 436140 496839
rect 436100 427168 436152 427174
rect 436100 427110 436152 427116
rect 434720 426284 434772 426290
rect 434720 426226 434772 426232
rect 437492 425814 437520 496975
rect 437570 496904 437626 496913
rect 437570 496839 437626 496848
rect 438858 496904 438914 496913
rect 438858 496839 438914 496848
rect 437584 483682 437612 496839
rect 437572 483676 437624 483682
rect 437572 483618 437624 483624
rect 438872 427242 438900 496839
rect 438860 427236 438912 427242
rect 438860 427178 438912 427184
rect 440252 425882 440280 498063
rect 441618 497040 441674 497049
rect 441618 496975 441674 496984
rect 443090 497040 443146 497049
rect 443090 496975 443146 496984
rect 445850 497040 445906 497049
rect 445850 496975 445906 496984
rect 447138 497040 447194 497049
rect 447138 496975 447194 496984
rect 448610 497040 448666 497049
rect 448610 496975 448666 496984
rect 449990 497040 450046 497049
rect 449990 496975 450046 496984
rect 452658 497040 452714 497049
rect 452658 496975 452714 496984
rect 440330 496904 440386 496913
rect 440330 496839 440386 496848
rect 440344 427310 440372 496839
rect 441632 427378 441660 496975
rect 441710 496904 441766 496913
rect 441710 496839 441766 496848
rect 442998 496904 443054 496913
rect 442998 496839 443054 496848
rect 441724 478174 441752 496839
rect 441712 478168 441764 478174
rect 441712 478110 441764 478116
rect 441620 427372 441672 427378
rect 441620 427314 441672 427320
rect 440332 427304 440384 427310
rect 440332 427246 440384 427252
rect 443012 425950 443040 496839
rect 443104 482390 443132 496975
rect 444378 496904 444434 496913
rect 444378 496839 444434 496848
rect 443092 482384 443144 482390
rect 443092 482326 443144 482332
rect 444392 427446 444420 496839
rect 445864 476882 445892 496975
rect 445942 496904 445998 496913
rect 445942 496839 445998 496848
rect 445852 476876 445904 476882
rect 445852 476818 445904 476824
rect 445760 428664 445812 428670
rect 445760 428606 445812 428612
rect 444380 427440 444432 427446
rect 444380 427382 444432 427388
rect 443000 425944 443052 425950
rect 443000 425886 443052 425892
rect 440240 425876 440292 425882
rect 440240 425818 440292 425824
rect 437480 425808 437532 425814
rect 437480 425750 437532 425756
rect 430672 424380 430724 424386
rect 430672 424322 430724 424328
rect 428464 423224 428516 423230
rect 428464 423166 428516 423172
rect 427084 423156 427136 423162
rect 427084 423098 427136 423104
rect 419540 422884 419592 422890
rect 419540 422826 419592 422832
rect 412732 422816 412784 422822
rect 412732 422758 412784 422764
rect 412640 422748 412692 422754
rect 412640 422690 412692 422696
rect 412086 418976 412142 418985
rect 412086 418911 412088 418920
rect 412140 418911 412142 418920
rect 412088 418882 412140 418888
rect 412652 418810 412680 422690
rect 412640 418804 412692 418810
rect 412640 418746 412692 418752
rect 412744 417450 412772 422758
rect 416136 422680 416188 422686
rect 416136 422622 416188 422628
rect 416044 422544 416096 422550
rect 416044 422486 416096 422492
rect 413284 421320 413336 421326
rect 413284 421262 413336 421268
rect 412732 417444 412784 417450
rect 412732 417386 412784 417392
rect 412086 416936 412142 416945
rect 412086 416871 412088 416880
rect 412140 416871 412142 416880
rect 412088 416842 412140 416848
rect 411994 396400 412050 396409
rect 411994 396335 412050 396344
rect 413296 393310 413324 421262
rect 413560 421252 413612 421258
rect 413560 421194 413612 421200
rect 413376 420300 413428 420306
rect 413376 420242 413428 420248
rect 413388 404326 413416 420242
rect 413468 420232 413520 420238
rect 413468 420174 413520 420180
rect 413480 407114 413508 420174
rect 413572 412010 413600 421194
rect 414756 420980 414808 420986
rect 414756 420922 414808 420928
rect 414664 420164 414716 420170
rect 414664 420106 414716 420112
rect 413836 418940 413888 418946
rect 413836 418882 413888 418888
rect 413652 416900 413704 416906
rect 413652 416842 413704 416848
rect 413560 412004 413612 412010
rect 413560 411946 413612 411952
rect 413664 409834 413692 416842
rect 413652 409828 413704 409834
rect 413652 409770 413704 409776
rect 413468 407108 413520 407114
rect 413468 407050 413520 407056
rect 413376 404320 413428 404326
rect 413376 404262 413428 404268
rect 413468 400240 413520 400246
rect 413468 400182 413520 400188
rect 413284 393304 413336 393310
rect 413284 393246 413336 393252
rect 413376 391264 413428 391270
rect 413376 391206 413428 391212
rect 411996 390312 412048 390318
rect 411994 390280 411996 390289
rect 412048 390280 412050 390289
rect 411994 390215 412050 390224
rect 411902 388240 411958 388249
rect 411902 388175 411958 388184
rect 411810 386064 411866 386073
rect 411810 385999 411866 386008
rect 411810 384024 411866 384033
rect 411810 383959 411866 383968
rect 411824 383722 411852 383959
rect 411812 383716 411864 383722
rect 411812 383658 411864 383664
rect 411732 382078 411852 382106
rect 411718 381984 411774 381993
rect 411718 381919 411774 381928
rect 411732 380934 411760 381919
rect 411720 380928 411772 380934
rect 411720 380870 411772 380876
rect 411824 375873 411852 382078
rect 412178 379944 412234 379953
rect 412178 379879 412234 379888
rect 411810 375864 411866 375873
rect 411810 375799 411866 375808
rect 411626 351112 411682 351121
rect 411626 351047 411682 351056
rect 411534 322416 411590 322425
rect 411534 322351 411590 322360
rect 411536 302184 411588 302190
rect 411536 302126 411588 302132
rect 411548 301753 411576 302126
rect 411534 301744 411590 301753
rect 411534 301679 411590 301688
rect 411628 250504 411680 250510
rect 411628 250446 411680 250452
rect 411640 248414 411668 250446
rect 411640 248386 411760 248414
rect 411534 225720 411590 225729
rect 411534 225655 411590 225664
rect 411548 225622 411576 225655
rect 411536 225616 411588 225622
rect 411536 225558 411588 225564
rect 411444 199912 411496 199918
rect 411444 199854 411496 199860
rect 411352 197872 411404 197878
rect 411352 197814 411404 197820
rect 410706 194032 410762 194041
rect 410706 193967 410762 193976
rect 410614 193896 410670 193905
rect 410614 193831 410670 193840
rect 410524 144288 410576 144294
rect 410524 144230 410576 144236
rect 411548 142866 411576 225558
rect 411626 209264 411682 209273
rect 411626 209199 411682 209208
rect 411640 209098 411668 209199
rect 411628 209092 411680 209098
rect 411628 209034 411680 209040
rect 411536 142860 411588 142866
rect 411536 142802 411588 142808
rect 411640 141642 411668 209034
rect 411732 197810 411760 248386
rect 411810 248296 411866 248305
rect 411810 248231 411866 248240
rect 411824 247722 411852 248231
rect 411812 247716 411864 247722
rect 411812 247658 411864 247664
rect 411824 199646 411852 247658
rect 412088 231124 412140 231130
rect 412088 231066 412140 231072
rect 412100 229094 412128 231066
rect 411916 229066 412128 229094
rect 411812 199640 411864 199646
rect 411812 199582 411864 199588
rect 411720 197804 411772 197810
rect 411720 197746 411772 197752
rect 411916 196722 411944 229066
rect 411996 220108 412048 220114
rect 411996 220050 412048 220056
rect 412008 219609 412036 220050
rect 411994 219600 412050 219609
rect 411994 219535 412050 219544
rect 411904 196716 411956 196722
rect 411904 196658 411956 196664
rect 412008 196654 412036 219535
rect 412088 216640 412140 216646
rect 412088 216582 412140 216588
rect 412100 215393 412128 216582
rect 412086 215384 412142 215393
rect 412086 215319 412142 215328
rect 412192 199850 412220 379879
rect 413284 379568 413336 379574
rect 413284 379510 413336 379516
rect 412270 367568 412326 367577
rect 412270 367503 412326 367512
rect 412284 200054 412312 367503
rect 412546 361448 412602 361457
rect 412602 361406 412772 361434
rect 412546 361383 412602 361392
rect 412640 202156 412692 202162
rect 412640 202098 412692 202104
rect 412272 200048 412324 200054
rect 412272 199990 412324 199996
rect 412180 199844 412232 199850
rect 412180 199786 412232 199792
rect 412652 198558 412680 202098
rect 412640 198552 412692 198558
rect 412640 198494 412692 198500
rect 411996 196648 412048 196654
rect 411996 196590 412048 196596
rect 412744 146946 412772 361406
rect 412916 359372 412968 359378
rect 412916 359314 412968 359320
rect 412822 334656 412878 334665
rect 412822 334591 412878 334600
rect 412836 149734 412864 334591
rect 412928 189786 412956 359314
rect 413008 343732 413060 343738
rect 413008 343674 413060 343680
rect 413020 192506 413048 343674
rect 413296 300830 413324 379510
rect 413388 353190 413416 391206
rect 413480 390318 413508 400182
rect 413468 390312 413520 390318
rect 413468 390254 413520 390260
rect 413376 353184 413428 353190
rect 413376 353126 413428 353132
rect 413284 300824 413336 300830
rect 413284 300766 413336 300772
rect 413100 273216 413152 273222
rect 413100 273158 413152 273164
rect 413112 195702 413140 273158
rect 413192 211812 413244 211818
rect 413192 211754 413244 211760
rect 413204 198490 413232 211754
rect 413376 204332 413428 204338
rect 413376 204274 413428 204280
rect 413388 198694 413416 204274
rect 413376 198688 413428 198694
rect 413376 198630 413428 198636
rect 413192 198484 413244 198490
rect 413192 198426 413244 198432
rect 413100 195696 413152 195702
rect 413100 195638 413152 195644
rect 413008 192500 413060 192506
rect 413008 192442 413060 192448
rect 412916 189780 412968 189786
rect 412916 189722 412968 189728
rect 412824 149728 412876 149734
rect 412824 149670 412876 149676
rect 412732 146940 412784 146946
rect 412732 146882 412784 146888
rect 411628 141636 411680 141642
rect 411628 141578 411680 141584
rect 410248 140072 410300 140078
rect 413848 140049 413876 418882
rect 414676 398818 414704 420106
rect 414768 408474 414796 420922
rect 414848 420096 414900 420102
rect 414848 420038 414900 420044
rect 414860 411942 414888 420038
rect 414848 411936 414900 411942
rect 414848 411878 414900 411884
rect 414756 408468 414808 408474
rect 414756 408410 414808 408416
rect 414664 398812 414716 398818
rect 414664 398754 414716 398760
rect 415308 362976 415360 362982
rect 415308 362918 415360 362924
rect 414848 360256 414900 360262
rect 414848 360198 414900 360204
rect 414756 357468 414808 357474
rect 414756 357410 414808 357416
rect 414664 310548 414716 310554
rect 414664 310490 414716 310496
rect 414020 276888 414072 276894
rect 414020 276830 414072 276836
rect 413928 204944 413980 204950
rect 413928 204886 413980 204892
rect 413940 204338 413968 204886
rect 413928 204332 413980 204338
rect 413928 204274 413980 204280
rect 414032 195634 414060 276830
rect 414112 267028 414164 267034
rect 414112 266970 414164 266976
rect 414124 198354 414152 266970
rect 414204 262880 414256 262886
rect 414204 262822 414256 262828
rect 414112 198348 414164 198354
rect 414112 198290 414164 198296
rect 414216 198082 414244 262822
rect 414296 258732 414348 258738
rect 414296 258674 414348 258680
rect 414308 198218 414336 258674
rect 414388 254584 414440 254590
rect 414388 254526 414440 254532
rect 414400 198286 414428 254526
rect 414480 241868 414532 241874
rect 414480 241810 414532 241816
rect 414388 198280 414440 198286
rect 414388 198222 414440 198228
rect 414296 198212 414348 198218
rect 414296 198154 414348 198160
rect 414204 198076 414256 198082
rect 414204 198018 414256 198024
rect 414492 195838 414520 241810
rect 414572 223644 414624 223650
rect 414572 223586 414624 223592
rect 414480 195832 414532 195838
rect 414480 195774 414532 195780
rect 414020 195628 414072 195634
rect 414020 195570 414072 195576
rect 414584 195226 414612 223586
rect 414676 213382 414704 310490
rect 414768 273222 414796 357410
rect 414860 276894 414888 360198
rect 414940 283620 414992 283626
rect 414940 283562 414992 283568
rect 414848 276888 414900 276894
rect 414848 276830 414900 276836
rect 414756 273216 414808 273222
rect 414756 273158 414808 273164
rect 414952 227798 414980 283562
rect 415320 279478 415348 362918
rect 416056 291854 416084 422486
rect 416148 294642 416176 422622
rect 418988 422612 419040 422618
rect 418988 422554 419040 422560
rect 418804 421456 418856 421462
rect 418804 421398 418856 421404
rect 417424 421388 417476 421394
rect 417424 421330 417476 421336
rect 416780 380928 416832 380934
rect 416780 380870 416832 380876
rect 416228 331288 416280 331294
rect 416228 331230 416280 331236
rect 416136 294636 416188 294642
rect 416136 294578 416188 294584
rect 416044 291848 416096 291854
rect 416044 291790 416096 291796
rect 415400 289128 415452 289134
rect 415400 289070 415452 289076
rect 415412 288454 415440 289070
rect 415400 288448 415452 288454
rect 415400 288390 415452 288396
rect 415308 279472 415360 279478
rect 415308 279414 415360 279420
rect 414940 227792 414992 227798
rect 414940 227734 414992 227740
rect 415308 224256 415360 224262
rect 415308 224198 415360 224204
rect 415320 223650 415348 224198
rect 415308 223644 415360 223650
rect 415308 223586 415360 223592
rect 414756 217320 414808 217326
rect 414756 217262 414808 217268
rect 414664 213376 414716 213382
rect 414664 213318 414716 213324
rect 414572 195220 414624 195226
rect 414572 195162 414624 195168
rect 414676 192778 414704 213318
rect 414768 198422 414796 217262
rect 415308 203584 415360 203590
rect 415308 203526 415360 203532
rect 415320 203114 415348 203526
rect 414848 203108 414900 203114
rect 414848 203050 414900 203056
rect 415308 203108 415360 203114
rect 415308 203050 415360 203056
rect 414756 198416 414808 198422
rect 414756 198358 414808 198364
rect 414860 192914 414888 203050
rect 415412 199986 415440 288390
rect 415492 274712 415544 274718
rect 415492 274654 415544 274660
rect 415400 199980 415452 199986
rect 415400 199922 415452 199928
rect 415504 198150 415532 274654
rect 415584 270564 415636 270570
rect 415584 270506 415636 270512
rect 415492 198144 415544 198150
rect 415492 198086 415544 198092
rect 415596 198014 415624 270506
rect 415676 263628 415728 263634
rect 415676 263570 415728 263576
rect 415584 198008 415636 198014
rect 415584 197950 415636 197956
rect 415688 195430 415716 263570
rect 416240 240106 416268 331230
rect 416688 275324 416740 275330
rect 416688 275266 416740 275272
rect 416700 274718 416728 275266
rect 416688 274712 416740 274718
rect 416688 274654 416740 274660
rect 416688 271176 416740 271182
rect 416688 271118 416740 271124
rect 416700 270570 416728 271118
rect 416688 270564 416740 270570
rect 416688 270506 416740 270512
rect 416228 240100 416280 240106
rect 416228 240042 416280 240048
rect 416688 238060 416740 238066
rect 416688 238002 416740 238008
rect 416700 237454 416728 238002
rect 415768 237448 415820 237454
rect 415768 237390 415820 237396
rect 416688 237448 416740 237454
rect 416688 237390 416740 237396
rect 415780 195566 415808 237390
rect 415860 233300 415912 233306
rect 415860 233242 415912 233248
rect 415872 195906 415900 233242
rect 415952 229764 416004 229770
rect 415952 229706 416004 229712
rect 415964 229158 415992 229706
rect 415952 229152 416004 229158
rect 415952 229094 416004 229100
rect 415964 195974 415992 229094
rect 415952 195968 416004 195974
rect 415952 195910 416004 195916
rect 415860 195900 415912 195906
rect 415860 195842 415912 195848
rect 415768 195560 415820 195566
rect 415768 195502 415820 195508
rect 415676 195424 415728 195430
rect 415676 195366 415728 195372
rect 414848 192908 414900 192914
rect 414848 192850 414900 192856
rect 414664 192772 414716 192778
rect 414664 192714 414716 192720
rect 416792 192574 416820 380870
rect 416872 279472 416924 279478
rect 416872 279414 416924 279420
rect 416884 192710 416912 279414
rect 416964 268388 417016 268394
rect 416964 268330 417016 268336
rect 416976 267782 417004 268330
rect 416964 267776 417016 267782
rect 416964 267718 417016 267724
rect 416976 195537 417004 267718
rect 417056 259480 417108 259486
rect 417056 259422 417108 259428
rect 416962 195528 417018 195537
rect 417068 195498 417096 259422
rect 417332 256012 417384 256018
rect 417332 255954 417384 255960
rect 417344 255338 417372 255954
rect 417148 255332 417200 255338
rect 417148 255274 417200 255280
rect 417332 255332 417384 255338
rect 417332 255274 417384 255280
rect 417160 195770 417188 255274
rect 417332 246356 417384 246362
rect 417332 246298 417384 246304
rect 417344 245682 417372 246298
rect 417332 245676 417384 245682
rect 417332 245618 417384 245624
rect 417344 238754 417372 245618
rect 417252 238726 417372 238754
rect 417148 195764 417200 195770
rect 417148 195706 417200 195712
rect 416962 195463 417018 195472
rect 417056 195492 417108 195498
rect 417056 195434 417108 195440
rect 417252 195362 417280 238726
rect 417240 195356 417292 195362
rect 417240 195298 417292 195304
rect 416872 192704 416924 192710
rect 416872 192646 416924 192652
rect 416780 192568 416832 192574
rect 416780 192510 416832 192516
rect 417436 142934 417464 421330
rect 417516 409896 417568 409902
rect 417516 409838 417568 409844
rect 417528 198393 417556 409838
rect 417700 385688 417752 385694
rect 417700 385630 417752 385636
rect 417608 338156 417660 338162
rect 417608 338098 417660 338104
rect 417620 247722 417648 338098
rect 417712 338094 417740 385630
rect 417700 338088 417752 338094
rect 417700 338030 417752 338036
rect 417700 330540 417752 330546
rect 417700 330482 417752 330488
rect 417608 247716 417660 247722
rect 417608 247658 417660 247664
rect 417712 244254 417740 330482
rect 417792 322244 417844 322250
rect 417792 322186 417844 322192
rect 417804 309126 417832 322186
rect 417792 309120 417844 309126
rect 417792 309062 417844 309068
rect 418160 287088 418212 287094
rect 418160 287030 418212 287036
rect 417700 244248 417752 244254
rect 417700 244190 417752 244196
rect 417514 198384 417570 198393
rect 417514 198319 417570 198328
rect 418172 192642 418200 287030
rect 418252 283688 418304 283694
rect 418252 283630 418304 283636
rect 418264 282946 418292 283630
rect 418252 282940 418304 282946
rect 418252 282882 418304 282888
rect 418264 195090 418292 282882
rect 418344 280832 418396 280838
rect 418344 280774 418396 280780
rect 418356 280226 418384 280774
rect 418344 280220 418396 280226
rect 418344 280162 418396 280168
rect 418356 197946 418384 280162
rect 418344 197940 418396 197946
rect 418344 197882 418396 197888
rect 418252 195084 418304 195090
rect 418252 195026 418304 195032
rect 418160 192636 418212 192642
rect 418160 192578 418212 192584
rect 417424 142928 417476 142934
rect 417424 142870 417476 142876
rect 418816 142866 418844 421398
rect 418896 411324 418948 411330
rect 418896 411266 418948 411272
rect 418908 143546 418936 411266
rect 419000 298110 419028 422554
rect 419172 332648 419224 332654
rect 419172 332590 419224 332596
rect 419080 314696 419132 314702
rect 419080 314638 419132 314644
rect 418988 298104 419040 298110
rect 418988 298046 419040 298052
rect 419092 220114 419120 314638
rect 419184 241874 419212 332590
rect 419172 241868 419224 241874
rect 419172 241810 419224 241816
rect 419080 220108 419132 220114
rect 419080 220050 419132 220056
rect 418896 143540 418948 143546
rect 418896 143482 418948 143488
rect 418804 142860 418856 142866
rect 418804 142802 418856 142808
rect 418908 142154 418936 143482
rect 418632 142126 418936 142154
rect 410248 140014 410300 140020
rect 413834 140040 413890 140049
rect 413834 139975 413890 139984
rect 418632 139890 418660 142126
rect 419552 141506 419580 422826
rect 431316 422476 431368 422482
rect 431316 422418 431368 422424
rect 420184 422408 420236 422414
rect 420184 422350 420236 422356
rect 420196 294710 420224 422350
rect 429200 421184 429252 421190
rect 429200 421126 429252 421132
rect 421656 420028 421708 420034
rect 421656 419970 421708 419976
rect 420368 350600 420420 350606
rect 420368 350542 420420 350548
rect 420276 320884 420328 320890
rect 420276 320826 420328 320832
rect 420184 294704 420236 294710
rect 420184 294646 420236 294652
rect 419632 293276 419684 293282
rect 419632 293218 419684 293224
rect 419644 292602 419672 293218
rect 419632 292596 419684 292602
rect 419632 292538 419684 292544
rect 419644 292074 419672 292538
rect 419644 292046 419764 292074
rect 419632 291916 419684 291922
rect 419632 291858 419684 291864
rect 419644 291242 419672 291858
rect 419632 291236 419684 291242
rect 419632 291178 419684 291184
rect 419644 192982 419672 291178
rect 419736 199578 419764 292046
rect 419816 284980 419868 284986
rect 419816 284922 419868 284928
rect 419828 284374 419856 284922
rect 419816 284368 419868 284374
rect 419816 284310 419868 284316
rect 419828 199782 419856 284310
rect 420288 233306 420316 320826
rect 420380 263634 420408 350542
rect 421564 313336 421616 313342
rect 421564 313278 421616 313284
rect 420920 309800 420972 309806
rect 420920 309742 420972 309748
rect 420932 309194 420960 309742
rect 420920 309188 420972 309194
rect 420920 309130 420972 309136
rect 420368 263628 420420 263634
rect 420368 263570 420420 263576
rect 420276 233300 420328 233306
rect 420276 233242 420328 233248
rect 419816 199776 419868 199782
rect 419816 199718 419868 199724
rect 419724 199572 419776 199578
rect 419724 199514 419776 199520
rect 419632 192976 419684 192982
rect 419632 192918 419684 192924
rect 420932 192846 420960 309130
rect 421012 304292 421064 304298
rect 421012 304234 421064 304240
rect 421024 303686 421052 304234
rect 421012 303680 421064 303686
rect 421012 303622 421064 303628
rect 421024 195158 421052 303622
rect 421012 195152 421064 195158
rect 421012 195094 421064 195100
rect 420920 192840 420972 192846
rect 420920 192782 420972 192788
rect 421576 149734 421604 313278
rect 421668 298042 421696 419970
rect 424416 419960 424468 419966
rect 424416 419902 424468 419908
rect 422944 376780 422996 376786
rect 422944 376722 422996 376728
rect 421932 375420 421984 375426
rect 421932 375362 421984 375368
rect 421840 328500 421892 328506
rect 421840 328442 421892 328448
rect 421748 313336 421800 313342
rect 421748 313278 421800 313284
rect 421656 298036 421708 298042
rect 421656 297978 421708 297984
rect 421760 217326 421788 313278
rect 421852 237386 421880 328442
rect 421944 296682 421972 375362
rect 422956 297974 422984 376722
rect 423128 347812 423180 347818
rect 423128 347754 423180 347760
rect 423036 342372 423088 342378
rect 423036 342314 423088 342320
rect 422944 297968 422996 297974
rect 422944 297910 422996 297916
rect 421932 296676 421984 296682
rect 421932 296618 421984 296624
rect 422944 295996 422996 296002
rect 422944 295938 422996 295944
rect 421840 237380 421892 237386
rect 421840 237322 421892 237328
rect 421748 217320 421800 217326
rect 421748 217262 421800 217268
rect 422956 200802 422984 295938
rect 423048 254590 423076 342314
rect 423140 259486 423168 347754
rect 424324 311908 424376 311914
rect 424324 311850 424376 311856
rect 423128 259480 423180 259486
rect 423128 259422 423180 259428
rect 423036 254584 423088 254590
rect 423036 254526 423088 254532
rect 422944 200796 422996 200802
rect 422944 200738 422996 200744
rect 424336 151094 424364 311850
rect 424428 297838 424456 419902
rect 428556 419892 428608 419898
rect 428556 419834 428608 419840
rect 425888 419756 425940 419762
rect 425888 419698 425940 419704
rect 425704 398880 425756 398886
rect 425704 398822 425756 398828
rect 424600 369912 424652 369918
rect 424600 369854 424652 369860
rect 424508 353320 424560 353326
rect 424508 353262 424560 353268
rect 424416 297832 424468 297838
rect 424416 297774 424468 297780
rect 424520 267034 424548 353262
rect 424612 287094 424640 369854
rect 424692 307080 424744 307086
rect 424692 307022 424744 307028
rect 424600 287088 424652 287094
rect 424600 287030 424652 287036
rect 424508 267028 424560 267034
rect 424508 266970 424560 266976
rect 424704 225622 424732 307022
rect 424692 225616 424744 225622
rect 424692 225558 424744 225564
rect 425716 198830 425744 398822
rect 425796 317484 425848 317490
rect 425796 317426 425848 317432
rect 425704 198824 425756 198830
rect 425704 198766 425756 198772
rect 424324 151088 424376 151094
rect 424324 151030 424376 151036
rect 421564 149728 421616 149734
rect 421564 149670 421616 149676
rect 425808 148374 425836 317426
rect 425900 297770 425928 419698
rect 426072 371340 426124 371346
rect 426072 371282 426124 371288
rect 425980 336796 426032 336802
rect 425980 336738 426032 336744
rect 425888 297764 425940 297770
rect 425888 297706 425940 297712
rect 425992 246362 426020 336738
rect 426084 289134 426112 371282
rect 427084 354748 427136 354754
rect 427084 354690 427136 354696
rect 426072 289128 426124 289134
rect 426072 289070 426124 289076
rect 427096 268394 427124 354690
rect 427176 326392 427228 326398
rect 427176 326334 427228 326340
rect 427084 268388 427136 268394
rect 427084 268330 427136 268336
rect 427188 252550 427216 326334
rect 428464 316056 428516 316062
rect 428464 315998 428516 316004
rect 427176 252544 427228 252550
rect 427176 252486 427228 252492
rect 425980 246356 426032 246362
rect 425980 246298 426032 246304
rect 428476 153882 428504 315998
rect 428568 297906 428596 419834
rect 428832 380928 428884 380934
rect 428832 380870 428884 380876
rect 428740 356108 428792 356114
rect 428740 356050 428792 356056
rect 428648 305040 428700 305046
rect 428648 304982 428700 304988
rect 428556 297900 428608 297906
rect 428556 297842 428608 297848
rect 428660 207670 428688 304982
rect 428752 271182 428780 356050
rect 428844 302190 428872 380870
rect 428832 302184 428884 302190
rect 428832 302126 428884 302132
rect 428832 300144 428884 300150
rect 428832 300086 428884 300092
rect 428740 271176 428792 271182
rect 428740 271118 428792 271124
rect 428844 229770 428872 300086
rect 428832 229764 428884 229770
rect 428832 229706 428884 229712
rect 428648 207664 428700 207670
rect 428648 207606 428700 207612
rect 428464 153876 428516 153882
rect 428464 153818 428516 153824
rect 429212 151814 429240 421126
rect 430120 383784 430172 383790
rect 430120 383726 430172 383732
rect 430028 346452 430080 346458
rect 430028 346394 430080 346400
rect 429936 345092 429988 345098
rect 429936 345034 429988 345040
rect 429844 318844 429896 318850
rect 429844 318786 429896 318792
rect 429856 224262 429884 318786
rect 429948 256018 429976 345034
rect 430040 258738 430068 346394
rect 430132 306338 430160 383726
rect 431224 325712 431276 325718
rect 431224 325654 431276 325660
rect 430120 306332 430172 306338
rect 430120 306274 430172 306280
rect 430028 258732 430080 258738
rect 430028 258674 430080 258680
rect 429936 256012 429988 256018
rect 429936 255954 429988 255960
rect 430028 256012 430080 256018
rect 430028 255954 430080 255960
rect 429844 224256 429896 224262
rect 429844 224198 429896 224204
rect 430040 203590 430068 255954
rect 430028 203584 430080 203590
rect 430028 203526 430080 203532
rect 431236 153202 431264 325654
rect 431328 297974 431356 422418
rect 435364 422340 435416 422346
rect 435364 422282 435416 422288
rect 432604 401668 432656 401674
rect 432604 401610 432656 401616
rect 431592 367124 431644 367130
rect 431592 367066 431644 367072
rect 431500 329928 431552 329934
rect 431500 329870 431552 329876
rect 431408 301504 431460 301510
rect 431408 301446 431460 301452
rect 431316 297968 431368 297974
rect 431316 297910 431368 297916
rect 431420 209098 431448 301446
rect 431512 238066 431540 329870
rect 431604 284986 431632 367066
rect 431960 317416 432012 317422
rect 431960 317358 432012 317364
rect 431972 309806 432000 317358
rect 431960 309800 432012 309806
rect 431960 309742 432012 309748
rect 431592 284980 431644 284986
rect 431592 284922 431644 284928
rect 431500 238060 431552 238066
rect 431500 238002 431552 238008
rect 431408 209092 431460 209098
rect 431408 209034 431460 209040
rect 432616 198626 432644 401610
rect 432972 374332 433024 374338
rect 432972 374274 433024 374280
rect 432880 365764 432932 365770
rect 432880 365706 432932 365712
rect 432696 307828 432748 307834
rect 432696 307770 432748 307776
rect 432708 211818 432736 307770
rect 432788 302252 432840 302258
rect 432788 302194 432840 302200
rect 432800 216646 432828 302194
rect 432892 283694 432920 365706
rect 432984 293282 433012 374274
rect 433984 364608 434036 364614
rect 433984 364550 434036 364556
rect 432972 293276 433024 293282
rect 432972 293218 433024 293224
rect 432880 283688 432932 283694
rect 432880 283630 432932 283636
rect 433996 280838 434024 364550
rect 434076 311908 434128 311914
rect 434076 311850 434128 311856
rect 433984 280832 434036 280838
rect 433984 280774 434036 280780
rect 434088 231130 434116 311850
rect 434076 231124 434128 231130
rect 434076 231066 434128 231072
rect 432788 216640 432840 216646
rect 432788 216582 432840 216588
rect 432696 211812 432748 211818
rect 432696 211754 432748 211760
rect 432604 198620 432656 198626
rect 432604 198562 432656 198568
rect 431224 153196 431276 153202
rect 431224 153138 431276 153144
rect 429212 151786 430160 151814
rect 425796 148368 425848 148374
rect 425796 148310 425848 148316
rect 419540 141500 419592 141506
rect 419540 141442 419592 141448
rect 406028 139862 406134 139890
rect 418278 139862 418660 139890
rect 430132 139890 430160 151786
rect 435376 141506 435404 422282
rect 438124 421116 438176 421122
rect 438124 421058 438176 421064
rect 437480 409828 437532 409834
rect 437480 409770 437532 409776
rect 437492 409193 437520 409770
rect 437478 409184 437534 409193
rect 437478 409119 437534 409128
rect 437480 408468 437532 408474
rect 437480 408410 437532 408416
rect 437492 407561 437520 408410
rect 437478 407552 437534 407561
rect 437478 407487 437534 407496
rect 437480 407108 437532 407114
rect 437480 407050 437532 407056
rect 437492 405929 437520 407050
rect 437478 405920 437534 405929
rect 437478 405855 437534 405864
rect 437480 404320 437532 404326
rect 437478 404288 437480 404297
rect 437532 404288 437534 404297
rect 437478 404223 437534 404232
rect 437478 402656 437534 402665
rect 437478 402591 437534 402600
rect 437492 401674 437520 402591
rect 437480 401668 437532 401674
rect 437480 401610 437532 401616
rect 437478 401024 437534 401033
rect 437478 400959 437534 400968
rect 437492 400246 437520 400959
rect 437480 400240 437532 400246
rect 437480 400182 437532 400188
rect 437478 399392 437534 399401
rect 437478 399327 437534 399336
rect 437492 398886 437520 399327
rect 437480 398880 437532 398886
rect 437480 398822 437532 398828
rect 437572 398812 437624 398818
rect 437572 398754 437624 398760
rect 437584 397769 437612 398754
rect 437570 397760 437626 397769
rect 437570 397695 437626 397704
rect 436742 396128 436798 396137
rect 436742 396063 436798 396072
rect 435456 389224 435508 389230
rect 435456 389166 435508 389172
rect 435468 198762 435496 389166
rect 435824 382288 435876 382294
rect 435824 382230 435876 382236
rect 435640 349172 435692 349178
rect 435640 349114 435692 349120
rect 435548 339516 435600 339522
rect 435548 339458 435600 339464
rect 435560 250510 435588 339458
rect 435652 262886 435680 349114
rect 435836 304298 435864 382230
rect 435824 304292 435876 304298
rect 435824 304234 435876 304240
rect 435732 303680 435784 303686
rect 435732 303622 435784 303628
rect 435640 262880 435692 262886
rect 435640 262822 435692 262828
rect 435548 250504 435600 250510
rect 435548 250446 435600 250452
rect 435744 222154 435772 303622
rect 435732 222148 435784 222154
rect 435732 222090 435784 222096
rect 436756 198966 436784 396063
rect 437570 394496 437626 394505
rect 437570 394431 437626 394440
rect 437480 393304 437532 393310
rect 437480 393246 437532 393252
rect 437492 392873 437520 393246
rect 437478 392864 437534 392873
rect 437478 392799 437534 392808
rect 437584 391270 437612 394431
rect 437572 391264 437624 391270
rect 437478 391232 437534 391241
rect 437572 391206 437624 391212
rect 437478 391167 437534 391176
rect 437492 385694 437520 391167
rect 437754 389600 437810 389609
rect 437754 389535 437810 389544
rect 437768 389230 437796 389535
rect 437756 389224 437808 389230
rect 437756 389166 437808 389172
rect 437480 385688 437532 385694
rect 437480 385630 437532 385636
rect 437478 384568 437534 384577
rect 437478 384503 437534 384512
rect 437492 383790 437520 384503
rect 437480 383784 437532 383790
rect 437480 383726 437532 383732
rect 437938 382936 437994 382945
rect 437938 382871 437994 382880
rect 437952 382294 437980 382871
rect 437940 382288 437992 382294
rect 437940 382230 437992 382236
rect 437478 381304 437534 381313
rect 437478 381239 437534 381248
rect 437492 380934 437520 381239
rect 437480 380928 437532 380934
rect 437480 380870 437532 380876
rect 437478 379672 437534 379681
rect 437478 379607 437534 379616
rect 437492 379574 437520 379607
rect 437480 379568 437532 379574
rect 437480 379510 437532 379516
rect 437478 378040 437534 378049
rect 437478 377975 437534 377984
rect 437492 376786 437520 377975
rect 437480 376780 437532 376786
rect 437480 376722 437532 376728
rect 437478 376408 437534 376417
rect 437478 376343 437534 376352
rect 437492 375426 437520 376343
rect 437480 375420 437532 375426
rect 437480 375362 437532 375368
rect 437478 374776 437534 374785
rect 437478 374711 437534 374720
rect 437492 374338 437520 374711
rect 437480 374332 437532 374338
rect 437480 374274 437532 374280
rect 437018 373144 437074 373153
rect 437018 373079 437074 373088
rect 436926 359952 436982 359961
rect 436926 359887 436982 359896
rect 436834 304192 436890 304201
rect 436834 304127 436890 304136
rect 436848 204950 436876 304127
rect 436940 275330 436968 359887
rect 437032 291922 437060 373079
rect 437478 371512 437534 371521
rect 437478 371447 437534 371456
rect 437492 371346 437520 371447
rect 437480 371340 437532 371346
rect 437480 371282 437532 371288
rect 437480 369912 437532 369918
rect 437478 369880 437480 369889
rect 437532 369880 437534 369889
rect 437478 369815 437534 369824
rect 437478 368248 437534 368257
rect 437478 368183 437534 368192
rect 437492 367130 437520 368183
rect 437480 367124 437532 367130
rect 437480 367066 437532 367072
rect 437478 366480 437534 366489
rect 437478 366415 437534 366424
rect 437492 365770 437520 366415
rect 437480 365764 437532 365770
rect 437480 365706 437532 365712
rect 437478 364848 437534 364857
rect 437478 364783 437534 364792
rect 437492 364614 437520 364783
rect 437480 364608 437532 364614
rect 437480 364550 437532 364556
rect 437478 363216 437534 363225
rect 437478 363151 437534 363160
rect 437492 362982 437520 363151
rect 437480 362976 437532 362982
rect 437480 362918 437532 362924
rect 437478 361584 437534 361593
rect 437478 361519 437534 361528
rect 437492 360262 437520 361519
rect 437480 360256 437532 360262
rect 437480 360198 437532 360204
rect 437478 358320 437534 358329
rect 437478 358255 437534 358264
rect 437492 357474 437520 358255
rect 437480 357468 437532 357474
rect 437480 357410 437532 357416
rect 437478 356688 437534 356697
rect 437478 356623 437534 356632
rect 437492 356114 437520 356623
rect 437480 356108 437532 356114
rect 437480 356050 437532 356056
rect 437478 355056 437534 355065
rect 437478 354991 437534 355000
rect 437492 354754 437520 354991
rect 437480 354748 437532 354754
rect 437480 354690 437532 354696
rect 437478 353424 437534 353433
rect 437478 353359 437534 353368
rect 437492 353326 437520 353359
rect 437480 353320 437532 353326
rect 437480 353262 437532 353268
rect 437478 351792 437534 351801
rect 437478 351727 437534 351736
rect 437492 350606 437520 351727
rect 437480 350600 437532 350606
rect 437480 350542 437532 350548
rect 437478 350160 437534 350169
rect 437478 350095 437534 350104
rect 437492 349178 437520 350095
rect 437480 349172 437532 349178
rect 437480 349114 437532 349120
rect 437478 348528 437534 348537
rect 437478 348463 437534 348472
rect 437492 347818 437520 348463
rect 437480 347812 437532 347818
rect 437480 347754 437532 347760
rect 437478 346896 437534 346905
rect 437478 346831 437534 346840
rect 437492 346458 437520 346831
rect 437480 346452 437532 346458
rect 437480 346394 437532 346400
rect 437478 345264 437534 345273
rect 437478 345199 437534 345208
rect 437492 345098 437520 345199
rect 437480 345092 437532 345098
rect 437480 345034 437532 345040
rect 437478 343496 437534 343505
rect 437478 343431 437534 343440
rect 437492 342378 437520 343431
rect 437480 342372 437532 342378
rect 437480 342314 437532 342320
rect 437846 340232 437902 340241
rect 437846 340167 437902 340176
rect 437860 339522 437888 340167
rect 437848 339516 437900 339522
rect 437848 339458 437900 339464
rect 437478 338600 437534 338609
rect 437478 338535 437534 338544
rect 437492 338162 437520 338535
rect 437480 338156 437532 338162
rect 437480 338098 437532 338104
rect 437478 336968 437534 336977
rect 437478 336903 437534 336912
rect 437492 336802 437520 336903
rect 437480 336796 437532 336802
rect 437480 336738 437532 336744
rect 437570 335336 437626 335345
rect 437570 335271 437626 335280
rect 437478 333704 437534 333713
rect 437478 333639 437534 333648
rect 437492 332654 437520 333639
rect 437480 332648 437532 332654
rect 437480 332590 437532 332596
rect 437478 332072 437534 332081
rect 437478 332007 437534 332016
rect 437492 331294 437520 332007
rect 437480 331288 437532 331294
rect 437480 331230 437532 331236
rect 437584 330546 437612 335271
rect 437572 330540 437624 330546
rect 437572 330482 437624 330488
rect 437478 330440 437534 330449
rect 437478 330375 437534 330384
rect 437492 329934 437520 330375
rect 437480 329928 437532 329934
rect 437480 329870 437532 329876
rect 437478 328808 437534 328817
rect 437478 328743 437534 328752
rect 437492 328506 437520 328743
rect 437480 328500 437532 328506
rect 437480 328442 437532 328448
rect 437478 327176 437534 327185
rect 437478 327111 437534 327120
rect 437492 320890 437520 327111
rect 437480 320884 437532 320890
rect 437480 320826 437532 320832
rect 437478 318880 437534 318889
rect 437478 318815 437480 318824
rect 437532 318815 437534 318824
rect 437480 318786 437532 318792
rect 437478 315616 437534 315625
rect 437478 315551 437534 315560
rect 437492 314702 437520 315551
rect 437480 314696 437532 314702
rect 437480 314638 437532 314644
rect 437478 313984 437534 313993
rect 437478 313919 437534 313928
rect 437492 313342 437520 313919
rect 437480 313336 437532 313342
rect 437480 313278 437532 313284
rect 438030 312352 438086 312361
rect 438030 312287 438086 312296
rect 437478 310720 437534 310729
rect 437478 310655 437534 310664
rect 437492 310554 437520 310655
rect 437480 310548 437532 310554
rect 437480 310490 437532 310496
rect 437478 309088 437534 309097
rect 437478 309023 437534 309032
rect 437492 307834 437520 309023
rect 437480 307828 437532 307834
rect 437480 307770 437532 307776
rect 437570 307456 437626 307465
rect 437570 307391 437626 307400
rect 437478 305824 437534 305833
rect 437478 305759 437534 305768
rect 437492 305046 437520 305759
rect 437480 305040 437532 305046
rect 437480 304982 437532 304988
rect 437584 301510 437612 307391
rect 438044 302258 438072 312287
rect 438032 302252 438084 302258
rect 438032 302194 438084 302200
rect 437572 301504 437624 301510
rect 437572 301446 437624 301452
rect 437020 291916 437072 291922
rect 437020 291858 437072 291864
rect 436928 275324 436980 275330
rect 436928 275266 436980 275272
rect 436836 204944 436888 204950
rect 436836 204886 436888 204892
rect 436744 198960 436796 198966
rect 436744 198902 436796 198908
rect 435456 198756 435508 198762
rect 435456 198698 435508 198704
rect 438136 141574 438164 421058
rect 445772 411398 445800 428606
rect 445956 426018 445984 496839
rect 447152 426086 447180 496975
rect 447230 496904 447286 496913
rect 447230 496839 447286 496848
rect 448518 496904 448574 496913
rect 448518 496839 448574 496848
rect 447244 472734 447272 496839
rect 447232 472728 447284 472734
rect 447232 472670 447284 472676
rect 448532 446486 448560 496839
rect 448624 475386 448652 496975
rect 449898 496904 449954 496913
rect 449898 496839 449954 496848
rect 448612 475380 448664 475386
rect 448612 475322 448664 475328
rect 448520 446480 448572 446486
rect 448520 446422 448572 446428
rect 449912 426222 449940 496839
rect 450004 479602 450032 496975
rect 451278 496904 451334 496913
rect 451278 496839 451334 496848
rect 449992 479596 450044 479602
rect 449992 479538 450044 479544
rect 451292 474094 451320 496839
rect 451280 474088 451332 474094
rect 451280 474030 451332 474036
rect 452672 430030 452700 496975
rect 452750 496904 452806 496913
rect 452750 496839 452806 496848
rect 454038 496904 454094 496913
rect 454038 496839 454094 496848
rect 452764 469878 452792 496839
rect 452752 469872 452804 469878
rect 452752 469814 452804 469820
rect 454052 447914 454080 496839
rect 454696 465730 454724 498063
rect 455800 494834 455828 498063
rect 462318 498063 462320 498072
rect 457444 498034 457496 498040
rect 462372 498063 462374 498072
rect 462320 498034 462372 498040
rect 456798 497312 456854 497321
rect 456798 497247 456854 497256
rect 456812 497010 456840 497247
rect 456800 497004 456852 497010
rect 456800 496946 456852 496952
rect 456890 496904 456946 496913
rect 456890 496839 456946 496848
rect 455788 494828 455840 494834
rect 455788 494770 455840 494776
rect 454684 465724 454736 465730
rect 454684 465666 454736 465672
rect 456904 449274 456932 496839
rect 456892 449268 456944 449274
rect 456892 449210 456944 449216
rect 454040 447908 454092 447914
rect 454040 447850 454092 447856
rect 457456 432750 457484 498034
rect 458270 497040 458326 497049
rect 458270 496975 458326 496984
rect 498198 497040 498254 497049
rect 498198 496975 498254 496984
rect 458178 496904 458234 496913
rect 458178 496839 458234 496848
rect 457444 432744 457496 432750
rect 457444 432686 457496 432692
rect 458192 431390 458220 496839
rect 458284 451994 458312 496975
rect 498212 496942 498240 496975
rect 494704 496936 494756 496942
rect 460938 496904 460994 496913
rect 460938 496839 460994 496848
rect 465078 496904 465134 496913
rect 465078 496839 465134 496848
rect 467838 496904 467894 496913
rect 467838 496839 467894 496848
rect 470598 496904 470654 496913
rect 470598 496839 470654 496848
rect 473358 496904 473414 496913
rect 473358 496839 473414 496848
rect 474738 496904 474794 496913
rect 474738 496839 474794 496848
rect 477498 496904 477554 496913
rect 480258 496904 480314 496913
rect 477498 496839 477554 496848
rect 479524 496868 479576 496874
rect 458272 451988 458324 451994
rect 458272 451930 458324 451936
rect 460952 434110 460980 496839
rect 465092 435470 465120 496839
rect 465080 435464 465132 435470
rect 465080 435406 465132 435412
rect 460940 434104 460992 434110
rect 460940 434046 460992 434052
rect 458180 431384 458232 431390
rect 458180 431326 458232 431332
rect 452660 430024 452712 430030
rect 452660 429966 452712 429972
rect 449900 426216 449952 426222
rect 449900 426158 449952 426164
rect 447140 426080 447192 426086
rect 447140 426022 447192 426028
rect 445944 426012 445996 426018
rect 445944 425954 445996 425960
rect 467852 424454 467880 496839
rect 470612 424590 470640 496839
rect 470600 424584 470652 424590
rect 470600 424526 470652 424532
rect 473372 424522 473400 496839
rect 474752 424726 474780 496839
rect 474740 424720 474792 424726
rect 474740 424662 474792 424668
rect 477512 424658 477540 496839
rect 480258 496839 480314 496848
rect 483018 496904 483074 496913
rect 483018 496839 483074 496848
rect 485778 496904 485834 496913
rect 485778 496839 485834 496848
rect 488538 496904 488594 496913
rect 488538 496839 488594 496848
rect 489918 496904 489974 496913
rect 489918 496839 489974 496848
rect 492678 496904 492734 496913
rect 498200 496936 498252 496942
rect 494704 496878 494756 496884
rect 495438 496904 495494 496913
rect 492678 496839 492734 496848
rect 479524 496810 479576 496816
rect 479536 440978 479564 496810
rect 479524 440972 479576 440978
rect 479524 440914 479576 440920
rect 480272 424862 480300 496839
rect 480260 424856 480312 424862
rect 480260 424798 480312 424804
rect 483032 424794 483060 496839
rect 485792 424930 485820 496839
rect 488552 424998 488580 496839
rect 489932 436898 489960 496839
rect 492692 438258 492720 496839
rect 494716 439618 494744 496878
rect 498200 496878 498252 496884
rect 500958 496904 501014 496913
rect 495438 496839 495440 496848
rect 495492 496839 495494 496848
rect 497464 496868 497516 496874
rect 495440 496810 495492 496816
rect 500958 496839 501014 496848
rect 502338 496904 502394 496913
rect 502338 496839 502394 496848
rect 505098 496904 505154 496913
rect 505098 496839 505100 496848
rect 497464 496810 497516 496816
rect 497476 445126 497504 496810
rect 497464 445120 497516 445126
rect 497464 445062 497516 445068
rect 500972 442338 501000 496839
rect 502352 443766 502380 496839
rect 505152 496839 505154 496848
rect 505100 496810 505152 496816
rect 502340 443760 502392 443766
rect 502340 443702 502392 443708
rect 500960 442332 501012 442338
rect 500960 442274 501012 442280
rect 494704 439612 494756 439618
rect 494704 439554 494756 439560
rect 492680 438252 492732 438258
rect 492680 438194 492732 438200
rect 489920 436892 489972 436898
rect 489920 436834 489972 436840
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 560944 430636 560996 430642
rect 560944 430578 560996 430584
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 488540 424992 488592 424998
rect 488540 424934 488592 424940
rect 485780 424924 485832 424930
rect 485780 424866 485832 424872
rect 483020 424788 483072 424794
rect 483020 424730 483072 424736
rect 477500 424652 477552 424658
rect 477500 424594 477552 424600
rect 473360 424516 473412 424522
rect 473360 424458 473412 424464
rect 467840 424448 467892 424454
rect 467840 424390 467892 424396
rect 552020 421592 552072 421598
rect 552020 421534 552072 421540
rect 551284 421048 551336 421054
rect 551284 420990 551336 420996
rect 482284 420368 482336 420374
rect 482284 420310 482336 420316
rect 470140 412004 470192 412010
rect 470140 411946 470192 411952
rect 439504 411392 439556 411398
rect 439504 411334 439556 411340
rect 445760 411392 445812 411398
rect 445760 411334 445812 411340
rect 438306 387832 438362 387841
rect 438306 387767 438362 387776
rect 438216 383716 438268 383722
rect 438216 383658 438268 383664
rect 438228 141642 438256 383658
rect 438320 317422 438348 387767
rect 438398 386200 438454 386209
rect 438398 386135 438454 386144
rect 438412 322250 438440 386135
rect 438490 341864 438546 341873
rect 438490 341799 438546 341808
rect 438504 326398 438532 341799
rect 438492 326392 438544 326398
rect 438492 326334 438544 326340
rect 438766 325544 438822 325553
rect 438766 325479 438822 325488
rect 438582 323912 438638 323921
rect 438582 323847 438638 323856
rect 438400 322244 438452 322250
rect 438400 322186 438452 322192
rect 438490 322144 438546 322153
rect 438490 322079 438546 322088
rect 438398 320512 438454 320521
rect 438398 320447 438454 320456
rect 438308 317416 438360 317422
rect 438308 317358 438360 317364
rect 438412 307086 438440 320447
rect 438400 307080 438452 307086
rect 438400 307022 438452 307028
rect 438306 302560 438362 302569
rect 438306 302495 438362 302504
rect 438320 256018 438348 302495
rect 438398 300928 438454 300937
rect 438398 300863 438454 300872
rect 438412 296002 438440 300863
rect 438400 295996 438452 296002
rect 438400 295938 438452 295944
rect 438504 283626 438532 322079
rect 438596 300150 438624 323847
rect 438674 317248 438730 317257
rect 438674 317183 438730 317192
rect 438688 303686 438716 317183
rect 438780 311914 438808 325479
rect 438768 311908 438820 311914
rect 438768 311850 438820 311856
rect 438676 303680 438728 303686
rect 438676 303622 438728 303628
rect 438584 300144 438636 300150
rect 438584 300086 438636 300092
rect 438492 283620 438544 283626
rect 438492 283562 438544 283568
rect 438308 256012 438360 256018
rect 438308 255954 438360 255960
rect 439516 147014 439544 411334
rect 445772 409986 445800 411334
rect 458272 411324 458324 411330
rect 458272 411266 458324 411272
rect 445772 409958 446108 409986
rect 458284 409850 458312 411266
rect 470152 409986 470180 411946
rect 482296 409986 482324 420310
rect 550640 419824 550692 419830
rect 550640 419766 550692 419772
rect 494520 419688 494572 419694
rect 494520 419630 494572 419636
rect 494532 409986 494560 419630
rect 506756 418804 506808 418810
rect 506756 418746 506808 418752
rect 506768 409986 506796 418746
rect 549904 418192 549956 418198
rect 549904 418134 549956 418140
rect 531320 417444 531372 417450
rect 531320 417386 531372 417392
rect 531332 409986 531360 417386
rect 543740 411936 543792 411942
rect 543740 411878 543792 411884
rect 543752 409986 543780 411878
rect 470152 409958 470488 409986
rect 482296 409958 482724 409986
rect 494532 409958 494960 409986
rect 506768 409958 507196 409986
rect 531332 409958 531668 409986
rect 543752 409958 543904 409986
rect 458252 409822 458312 409850
rect 519084 409896 519136 409902
rect 519136 409844 519432 409850
rect 519084 409838 519432 409844
rect 519096 409822 519432 409838
rect 439688 371272 439740 371278
rect 439688 371214 439740 371220
rect 439596 329860 439648 329866
rect 439596 329802 439648 329808
rect 439608 147014 439636 329802
rect 439700 293962 439728 371214
rect 439780 342304 439832 342310
rect 439780 342246 439832 342252
rect 439792 300830 439820 342246
rect 439872 324352 439924 324358
rect 439872 324294 439924 324300
rect 439780 300824 439832 300830
rect 439780 300766 439832 300772
rect 439884 300762 439912 324294
rect 439872 300756 439924 300762
rect 439872 300698 439924 300704
rect 443012 300070 444268 300098
rect 452732 300070 452792 300098
rect 439688 293956 439740 293962
rect 439688 293898 439740 293904
rect 441620 293956 441672 293962
rect 441620 293898 441672 293904
rect 441632 151814 441660 293898
rect 443012 179382 443040 300070
rect 452764 296714 452792 300070
rect 452672 296686 452792 296714
rect 460952 300070 461196 300098
rect 469232 300070 469660 300098
rect 477512 300070 478124 300098
rect 485792 300070 486588 300098
rect 494716 300070 495052 300098
rect 503180 300070 503516 300098
rect 511980 300070 512040 300098
rect 452672 193186 452700 296686
rect 460952 219434 460980 300070
rect 469232 233238 469260 300070
rect 477512 296002 477540 300070
rect 477500 295996 477552 296002
rect 477500 295938 477552 295944
rect 469220 233232 469272 233238
rect 469220 233174 469272 233180
rect 460940 219428 460992 219434
rect 460940 219370 460992 219376
rect 452660 193180 452712 193186
rect 452660 193122 452712 193128
rect 466460 182844 466512 182850
rect 466460 182786 466512 182792
rect 443000 179376 443052 179382
rect 443000 179318 443052 179324
rect 466472 151814 466500 182786
rect 441632 151786 442304 151814
rect 466472 151786 466776 151814
rect 439504 147008 439556 147014
rect 439504 146950 439556 146956
rect 439596 147008 439648 147014
rect 439596 146950 439648 146956
rect 438216 141636 438268 141642
rect 438216 141578 438268 141584
rect 438124 141568 438176 141574
rect 438124 141510 438176 141516
rect 435364 141500 435416 141506
rect 435364 141442 435416 141448
rect 442276 139890 442304 151786
rect 454684 142928 454736 142934
rect 454684 142870 454736 142876
rect 454696 139890 454724 142870
rect 466748 139890 466776 151786
rect 485792 146946 485820 300070
rect 494716 297770 494744 300070
rect 503180 297838 503208 300070
rect 512012 297906 512040 300070
rect 520292 300070 520444 300098
rect 528756 300070 528908 300098
rect 536852 300070 537372 300098
rect 545500 300070 545836 300098
rect 520292 297974 520320 300070
rect 522304 298172 522356 298178
rect 522304 298114 522356 298120
rect 520280 297968 520332 297974
rect 520280 297910 520332 297916
rect 512000 297900 512052 297906
rect 512000 297842 512052 297848
rect 503168 297832 503220 297838
rect 503168 297774 503220 297780
rect 494704 297764 494756 297770
rect 494704 297706 494756 297712
rect 512000 294704 512052 294710
rect 512000 294646 512052 294652
rect 510802 198112 510858 198121
rect 510802 198047 510858 198056
rect 510618 197976 510674 197985
rect 510618 197911 510674 197920
rect 503720 195288 503772 195294
rect 503720 195230 503772 195236
rect 485780 146940 485832 146946
rect 485780 146882 485832 146888
rect 479156 142860 479208 142866
rect 479156 142802 479208 142808
rect 479168 139890 479196 142802
rect 491298 142760 491354 142769
rect 491298 142695 491354 142704
rect 491312 139890 491340 142695
rect 503732 139890 503760 195230
rect 509240 191140 509292 191146
rect 509240 191082 509292 191088
rect 430132 139862 430514 139890
rect 442276 139862 442750 139890
rect 454696 139862 454986 139890
rect 466748 139862 467222 139890
rect 479168 139862 479458 139890
rect 491312 139862 491694 139890
rect 503732 139862 503930 139890
rect 401140 139596 401192 139602
rect 401140 139538 401192 139544
rect 401048 137896 401100 137902
rect 401048 137838 401100 137844
rect 400956 121440 401008 121446
rect 400956 121382 401008 121388
rect 400600 74506 400904 74534
rect 400600 70417 400628 74506
rect 400586 70408 400642 70417
rect 400586 70343 400642 70352
rect 509252 37262 509280 191082
rect 509332 141636 509384 141642
rect 509332 141578 509384 141584
rect 509240 37256 509292 37262
rect 509240 37198 509292 37204
rect 399758 35864 399814 35873
rect 399758 35799 399814 35808
rect 399772 34542 399800 35799
rect 399760 34536 399812 34542
rect 399760 34478 399812 34484
rect 404188 30110 404294 30138
rect 412758 30110 413048 30138
rect 421222 30110 421512 30138
rect 429686 30110 429976 30138
rect 438150 30110 438440 30138
rect 446614 30110 446904 30138
rect 399208 28824 399260 28830
rect 399208 28766 399260 28772
rect 398288 28756 398340 28762
rect 398288 28698 398340 28704
rect 404188 28558 404216 30110
rect 413020 28830 413048 30110
rect 413008 28824 413060 28830
rect 413008 28766 413060 28772
rect 421484 28762 421512 30110
rect 429948 29170 429976 30110
rect 438412 29238 438440 30110
rect 446876 29306 446904 30110
rect 454696 30110 455078 30138
rect 463160 30110 463542 30138
rect 472006 30110 472112 30138
rect 446864 29300 446916 29306
rect 446864 29242 446916 29248
rect 438400 29232 438452 29238
rect 438400 29174 438452 29180
rect 429936 29164 429988 29170
rect 429936 29106 429988 29112
rect 454696 28937 454724 30110
rect 454682 28928 454738 28937
rect 454682 28863 454738 28872
rect 421472 28756 421524 28762
rect 421472 28698 421524 28704
rect 463160 28626 463188 30110
rect 463148 28620 463200 28626
rect 463148 28562 463200 28568
rect 404176 28552 404228 28558
rect 404176 28494 404228 28500
rect 472084 28354 472112 30110
rect 480364 30110 480470 30138
rect 488934 30110 489224 30138
rect 497398 30110 497688 30138
rect 505862 30110 506152 30138
rect 480364 28694 480392 30110
rect 489196 28694 489224 30110
rect 497660 28898 497688 30110
rect 506124 28966 506152 30110
rect 506112 28960 506164 28966
rect 506112 28902 506164 28908
rect 497648 28892 497700 28898
rect 497648 28834 497700 28840
rect 509344 28694 509372 141578
rect 509424 141568 509476 141574
rect 509424 141510 509476 141516
rect 509436 28898 509464 141510
rect 510632 78577 510660 197911
rect 510712 141500 510764 141506
rect 510712 141442 510764 141448
rect 510618 78568 510674 78577
rect 510618 78503 510674 78512
rect 509516 37256 509568 37262
rect 509514 37224 509516 37233
rect 509568 37224 509570 37233
rect 509514 37159 509570 37168
rect 510724 28966 510752 141442
rect 510816 106185 510844 198047
rect 510896 155236 510948 155242
rect 510896 155178 510948 155184
rect 510802 106176 510858 106185
rect 510802 106111 510858 106120
rect 510908 64705 510936 155178
rect 512012 92449 512040 294646
rect 512184 294636 512236 294642
rect 512184 294578 512236 294584
rect 512092 291848 512144 291854
rect 512092 291790 512144 291796
rect 512104 119921 512132 291790
rect 512196 133657 512224 294578
rect 515404 271924 515456 271930
rect 515404 271866 515456 271872
rect 512276 147008 512328 147014
rect 512276 146950 512328 146956
rect 512182 133648 512238 133657
rect 512182 133583 512238 133592
rect 512090 119912 512146 119921
rect 512090 119847 512146 119856
rect 511998 92440 512054 92449
rect 511998 92375 512054 92384
rect 510894 64696 510950 64705
rect 510894 64631 510950 64640
rect 512288 50969 512316 146950
rect 512274 50960 512330 50969
rect 512274 50895 512330 50904
rect 515416 29034 515444 271866
rect 520924 244316 520976 244322
rect 520924 244258 520976 244264
rect 519544 205692 519596 205698
rect 519544 205634 519596 205640
rect 518164 141432 518216 141438
rect 518164 141374 518216 141380
rect 518176 46918 518204 141374
rect 518164 46912 518216 46918
rect 518164 46854 518216 46860
rect 519556 29102 519584 205634
rect 520936 29238 520964 244258
rect 522316 29306 522344 298114
rect 528756 298042 528784 300070
rect 528744 298036 528796 298042
rect 528744 297978 528796 297984
rect 536852 202162 536880 300070
rect 545500 298110 545528 300070
rect 545488 298104 545540 298110
rect 545488 298046 545540 298052
rect 544384 295996 544436 296002
rect 544384 295938 544436 295944
rect 536840 202156 536892 202162
rect 536840 202098 536892 202104
rect 544396 86970 544424 295938
rect 544384 86964 544436 86970
rect 544384 86906 544436 86912
rect 522304 29300 522356 29306
rect 522304 29242 522356 29248
rect 520924 29232 520976 29238
rect 520924 29174 520976 29180
rect 519544 29096 519596 29102
rect 519544 29038 519596 29044
rect 515404 29028 515456 29034
rect 515404 28970 515456 28976
rect 510712 28960 510764 28966
rect 510712 28902 510764 28908
rect 509424 28892 509476 28898
rect 509424 28834 509476 28840
rect 549916 28762 549944 418134
rect 550652 403073 550680 419766
rect 550638 403064 550694 403073
rect 550638 402999 550694 403008
rect 550546 306504 550602 306513
rect 550546 306439 550602 306448
rect 550560 300762 550588 306439
rect 550548 300756 550600 300762
rect 550548 300698 550600 300704
rect 551296 113150 551324 420990
rect 552032 361865 552060 421534
rect 552204 421524 552256 421530
rect 552204 421466 552256 421472
rect 552112 419552 552164 419558
rect 552112 419494 552164 419500
rect 552018 361856 552074 361865
rect 552018 361791 552074 361800
rect 552018 334384 552074 334393
rect 552018 334319 552074 334328
rect 551376 324352 551428 324358
rect 551376 324294 551428 324300
rect 551284 113144 551336 113150
rect 551284 113086 551336 113092
rect 549904 28756 549956 28762
rect 549904 28698 549956 28704
rect 480352 28688 480404 28694
rect 480352 28630 480404 28636
rect 489184 28688 489236 28694
rect 489184 28630 489236 28636
rect 509332 28688 509384 28694
rect 551388 28665 551416 324294
rect 552032 199442 552060 334319
rect 552124 320657 552152 419494
rect 552216 375601 552244 421466
rect 552296 419620 552348 419626
rect 552296 419562 552348 419568
rect 552308 389337 552336 419562
rect 552294 389328 552350 389337
rect 552294 389263 552350 389272
rect 554044 378208 554096 378214
rect 554044 378150 554096 378156
rect 552202 375592 552258 375601
rect 552202 375527 552258 375536
rect 552202 348120 552258 348129
rect 552202 348055 552258 348064
rect 552110 320648 552166 320657
rect 552110 320583 552166 320592
rect 552216 300830 552244 348055
rect 552204 300824 552256 300830
rect 552204 300766 552256 300772
rect 552020 199436 552072 199442
rect 552020 199378 552072 199384
rect 554056 28830 554084 378150
rect 558184 364404 558236 364410
rect 558184 364346 558236 364352
rect 556804 311908 556856 311914
rect 556804 311850 556856 311856
rect 555424 258120 555476 258126
rect 555424 258062 555476 258068
rect 554044 28824 554096 28830
rect 554044 28766 554096 28772
rect 509332 28630 509384 28636
rect 551374 28656 551430 28665
rect 551374 28591 551430 28600
rect 472072 28348 472124 28354
rect 472072 28290 472124 28296
rect 555436 28014 555464 258062
rect 556816 28801 556844 311850
rect 556802 28792 556858 28801
rect 556802 28727 556858 28736
rect 558196 28558 558224 364346
rect 560956 29170 560984 430578
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580184 418198 580212 418231
rect 580172 418192 580224 418198
rect 580172 418134 580224 418140
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580184 364410 580212 365055
rect 580172 364404 580224 364410
rect 580172 364346 580224 364352
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580184 311914 580212 312015
rect 580172 311908 580224 311914
rect 580172 311850 580224 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 579802 272232 579858 272241
rect 579802 272167 579858 272176
rect 579816 271930 579844 272167
rect 579804 271924 579856 271930
rect 579804 271866 579856 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 579802 245576 579858 245585
rect 579802 245511 579858 245520
rect 579816 244322 579844 245511
rect 579804 244316 579856 244322
rect 579804 244258 579856 244264
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580170 205728 580226 205737
rect 580170 205663 580172 205672
rect 580224 205663 580226 205672
rect 580172 205634 580224 205640
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580184 165646 580212 165815
rect 580172 165640 580224 165646
rect 580172 165582 580224 165588
rect 580632 153876 580684 153882
rect 580632 153818 580684 153824
rect 580172 153196 580224 153202
rect 580172 153138 580224 153144
rect 580184 152697 580212 153138
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580540 151088 580592 151094
rect 580540 151030 580592 151036
rect 580356 149728 580408 149734
rect 580356 149670 580408 149676
rect 580264 148368 580316 148374
rect 580264 148310 580316 148316
rect 562324 146940 562376 146946
rect 562324 146882 562376 146888
rect 562336 126954 562364 146882
rect 562324 126948 562376 126954
rect 562324 126890 562376 126896
rect 579712 126948 579764 126954
rect 579712 126890 579764 126896
rect 579724 126041 579752 126890
rect 579710 126032 579766 126041
rect 579710 125967 579766 125976
rect 579712 113144 579764 113150
rect 579712 113086 579764 113092
rect 579724 112849 579752 113086
rect 579710 112840 579766 112849
rect 579710 112775 579766 112784
rect 579988 86964 580040 86970
rect 579988 86906 580040 86912
rect 580000 86193 580028 86906
rect 579986 86184 580042 86193
rect 579986 86119 580042 86128
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 560944 29164 560996 29170
rect 560944 29106 560996 29112
rect 558184 28552 558236 28558
rect 558184 28494 558236 28500
rect 555424 28008 555476 28014
rect 555424 27950 555476 27956
rect 398012 27940 398064 27946
rect 398012 27882 398064 27888
rect 580276 19825 580304 148310
rect 580368 59673 580396 149670
rect 580448 144220 580500 144226
rect 580448 144162 580500 144168
rect 580460 73001 580488 144162
rect 580552 99521 580580 151030
rect 580644 139369 580672 153818
rect 580630 139360 580686 139369
rect 580630 139295 580686 139304
rect 580538 99512 580594 99521
rect 580538 99447 580594 99456
rect 580446 72992 580502 73001
rect 580446 72927 580502 72936
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580262 19816 580318 19825
rect 580262 19751 580318 19760
rect 284944 6860 284996 6866
rect 284944 6802 284996 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 1646 354 1758 480
rect 1412 326 1758 354
rect 542 -960 654 326
rect 1646 -960 1758 326
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 48042 536832 48098 536888
rect 47950 533704 48006 533760
rect 47858 530984 47914 531040
rect 47766 508000 47822 508056
rect 396630 536852 396686 536888
rect 396630 536832 396632 536852
rect 396632 536832 396684 536852
rect 396684 536832 396686 536852
rect 48226 535880 48282 535936
rect 48134 532752 48190 532808
rect 49514 529930 49570 529986
rect 49422 528162 49478 528218
rect 49330 508272 49386 508328
rect 49606 509938 49662 509994
rect 67546 498072 67602 498128
rect 73342 498072 73398 498128
rect 74354 498072 74410 498128
rect 78586 498072 78642 498128
rect 79874 498072 79930 498128
rect 81254 498072 81310 498128
rect 85946 498072 86002 498128
rect 86498 498072 86554 498128
rect 89534 498072 89590 498128
rect 92294 498072 92350 498128
rect 96526 498072 96582 498128
rect 103426 498072 103482 498128
rect 104806 498072 104862 498128
rect 113546 498072 113602 498128
rect 116858 498072 116914 498128
rect 118606 498072 118662 498128
rect 121366 498072 121422 498128
rect 126886 498072 126942 498128
rect 129646 498072 129702 498128
rect 146206 498072 146262 498128
rect 150990 498072 151046 498128
rect 154486 498072 154542 498128
rect 66166 496848 66222 496904
rect 73066 497392 73122 497448
rect 68926 496848 68982 496904
rect 70306 496848 70362 496904
rect 71686 496848 71742 496904
rect 75826 496848 75882 496904
rect 77206 496848 77262 496904
rect 78310 496868 78366 496904
rect 78310 496848 78312 496868
rect 78312 496848 78364 496868
rect 78364 496848 78366 496868
rect 81162 496984 81218 497040
rect 96342 497800 96398 497856
rect 84014 496984 84070 497040
rect 88154 496984 88210 497040
rect 93674 496984 93730 497040
rect 81254 496848 81310 496904
rect 82726 496848 82782 496904
rect 84106 496848 84162 496904
rect 85486 496848 85542 496904
rect 88246 496848 88302 496904
rect 89166 496848 89222 496904
rect 91006 496848 91062 496904
rect 91190 496848 91246 496904
rect 93766 496848 93822 496904
rect 95146 496848 95202 496904
rect 96434 496984 96490 497040
rect 99286 496984 99342 497040
rect 101954 496984 102010 497040
rect 97906 496848 97962 496904
rect 99194 496848 99250 496904
rect 100666 496848 100722 496904
rect 102046 496848 102102 496904
rect 103334 496848 103390 496904
rect 104714 496848 104770 496904
rect 106094 496984 106150 497040
rect 108854 496984 108910 497040
rect 106186 496848 106242 496904
rect 107566 496848 107622 496904
rect 108946 496848 109002 496904
rect 110326 496848 110382 496904
rect 111706 496848 111762 496904
rect 124126 496848 124182 496904
rect 28906 349968 28962 350024
rect 131026 496848 131082 496904
rect 131210 399064 131266 399120
rect 131210 398520 131266 398576
rect 131486 397296 131542 397352
rect 131302 396752 131358 396808
rect 131210 396228 131266 396264
rect 131210 396208 131212 396228
rect 131212 396208 131264 396228
rect 131264 396208 131266 396228
rect 131210 395528 131266 395584
rect 131302 394984 131358 395040
rect 131210 394440 131266 394496
rect 131210 393216 131266 393272
rect 131302 392128 131358 392184
rect 131210 391448 131266 391504
rect 131118 390360 131174 390416
rect 131486 390904 131542 390960
rect 131486 389816 131542 389872
rect 131210 389136 131266 389192
rect 131302 388592 131358 388648
rect 131210 388048 131266 388104
rect 131118 387368 131174 387424
rect 131210 386824 131266 386880
rect 131302 386280 131358 386336
rect 131118 385736 131174 385792
rect 131210 385092 131212 385112
rect 131212 385092 131264 385112
rect 131264 385092 131266 385112
rect 131210 385056 131266 385092
rect 131118 384512 131174 384568
rect 131210 383968 131266 384024
rect 131118 383424 131174 383480
rect 131210 382744 131266 382800
rect 131486 382200 131542 382256
rect 131210 380996 131266 381032
rect 131210 380976 131212 380996
rect 131212 380976 131264 380996
rect 131264 380976 131266 380996
rect 131210 380432 131266 380488
rect 131486 379888 131542 379944
rect 131118 379344 131174 379400
rect 131302 378664 131358 378720
rect 131210 378120 131266 378176
rect 131118 377576 131174 377632
rect 131210 377032 131266 377088
rect 131210 376352 131266 376408
rect 131486 375808 131542 375864
rect 131210 375264 131266 375320
rect 131118 374584 131174 374640
rect 131210 374060 131266 374096
rect 131210 374040 131212 374060
rect 131212 374040 131264 374060
rect 131264 374040 131266 374060
rect 131210 373496 131266 373552
rect 131486 372952 131542 373008
rect 131118 372272 131174 372328
rect 131210 371728 131266 371784
rect 131118 370640 131174 370696
rect 131210 369980 131266 370016
rect 131210 369960 131212 369980
rect 131212 369960 131264 369980
rect 131264 369960 131266 369980
rect 131210 369416 131266 369472
rect 131486 368872 131542 368928
rect 131210 368192 131266 368248
rect 131118 367648 131174 367704
rect 131210 367124 131266 367160
rect 131210 367104 131212 367124
rect 131212 367104 131264 367124
rect 131264 367104 131266 367124
rect 131210 365880 131266 365936
rect 131118 365336 131174 365392
rect 131210 364792 131266 364848
rect 131486 364248 131542 364304
rect 131118 363568 131174 363624
rect 131210 363044 131266 363080
rect 131210 363024 131212 363044
rect 131212 363024 131264 363044
rect 131264 363024 131266 363044
rect 131118 362480 131174 362536
rect 131210 361800 131266 361856
rect 131118 361256 131174 361312
rect 131210 360204 131212 360224
rect 131212 360204 131264 360224
rect 131264 360204 131266 360224
rect 131210 360168 131266 360204
rect 131210 358944 131266 359000
rect 131118 358400 131174 358456
rect 131210 357856 131266 357912
rect 131302 357176 131358 357232
rect 131118 356632 131174 356688
rect 131210 356088 131266 356144
rect 131302 355408 131358 355464
rect 131210 354864 131266 354920
rect 131118 354320 131174 354376
rect 131210 353776 131266 353832
rect 131210 353096 131266 353152
rect 131118 352552 131174 352608
rect 131486 352008 131542 352064
rect 131118 351464 131174 351520
rect 131210 350784 131266 350840
rect 131118 350240 131174 350296
rect 131210 349696 131266 349752
rect 131210 349016 131266 349072
rect 131302 348472 131358 348528
rect 131486 347928 131542 347984
rect 131118 347384 131174 347440
rect 131210 346704 131266 346760
rect 131210 346160 131266 346216
rect 131118 345616 131174 345672
rect 131210 345092 131266 345128
rect 131210 345072 131212 345092
rect 131212 345072 131264 345092
rect 131264 345072 131266 345092
rect 131302 344392 131358 344448
rect 131210 343848 131266 343904
rect 131210 343304 131266 343360
rect 131486 342624 131542 342680
rect 131118 342080 131174 342136
rect 131302 341536 131358 341592
rect 131210 341028 131212 341048
rect 131212 341028 131264 341048
rect 131264 341028 131266 341048
rect 131210 340992 131266 341028
rect 131302 340312 131358 340368
rect 131210 339768 131266 339824
rect 131118 339224 131174 339280
rect 131210 338680 131266 338736
rect 131486 338000 131542 338056
rect 131210 336932 131266 336968
rect 131210 336912 131212 336932
rect 131212 336912 131264 336932
rect 131264 336912 131266 336932
rect 131118 336232 131174 336288
rect 131210 335688 131266 335744
rect 131210 335144 131266 335200
rect 131118 333920 131174 333976
rect 131302 333376 131358 333432
rect 131210 332832 131266 332888
rect 131486 331608 131542 331664
rect 131118 331064 131174 331120
rect 131210 329860 131266 329896
rect 131210 329840 131212 329860
rect 131212 329840 131264 329860
rect 131264 329840 131266 329860
rect 131210 329296 131266 329352
rect 131302 328752 131358 328808
rect 131118 328208 131174 328264
rect 131210 327528 131266 327584
rect 131302 326440 131358 326496
rect 131210 325896 131266 325952
rect 131210 325216 131266 325272
rect 131486 324672 131542 324728
rect 131118 324128 131174 324184
rect 131486 323448 131542 323504
rect 131210 322940 131212 322960
rect 131212 322940 131264 322960
rect 131264 322940 131266 322960
rect 131210 322904 131266 322940
rect 131118 322360 131174 322416
rect 131210 321816 131266 321872
rect 131118 321136 131174 321192
rect 131210 320592 131266 320648
rect 131210 318844 131266 318880
rect 131210 318824 131212 318844
rect 131212 318824 131264 318844
rect 131264 318824 131266 318844
rect 131486 317736 131542 317792
rect 131210 316512 131266 316568
rect 131486 315968 131542 316024
rect 131210 315424 131266 315480
rect 131302 314744 131358 314800
rect 131118 314200 131174 314256
rect 131210 313656 131266 313712
rect 131302 313112 131358 313168
rect 131118 312432 131174 312488
rect 131210 311908 131266 311944
rect 131210 311888 131212 311908
rect 131212 311888 131264 311908
rect 131264 311888 131266 311908
rect 131210 311344 131266 311400
rect 131118 310120 131174 310176
rect 131486 310664 131542 310720
rect 131210 309576 131266 309632
rect 131118 309032 131174 309088
rect 131486 308352 131542 308408
rect 131210 307808 131266 307864
rect 131118 307264 131174 307320
rect 131210 306720 131266 306776
rect 131118 306040 131174 306096
rect 131486 305496 131542 305552
rect 131210 304988 131212 305008
rect 131212 304988 131264 305008
rect 131264 304988 131266 305008
rect 131210 304952 131266 304988
rect 131302 304272 131358 304328
rect 131210 303728 131266 303784
rect 131118 303184 131174 303240
rect 131210 302640 131266 302696
rect 131486 301960 131542 302016
rect 131210 300908 131212 300928
rect 131212 300908 131264 300928
rect 131264 300908 131266 300928
rect 131210 300872 131266 300908
rect 131118 300056 131174 300112
rect 131946 400152 132002 400208
rect 131946 397840 132002 397896
rect 132038 393760 132094 393816
rect 132038 392672 132094 392728
rect 132222 381656 132278 381712
rect 131946 371184 132002 371240
rect 132222 366560 132278 366616
rect 132130 360712 132186 360768
rect 132038 359488 132094 359544
rect 132038 337456 132094 337512
rect 132222 334600 132278 334656
rect 132222 332288 132278 332344
rect 132222 330520 132278 330576
rect 132222 326984 132278 327040
rect 131946 320048 132002 320104
rect 132222 319504 132278 319560
rect 132130 318280 132186 318336
rect 132038 301416 132094 301472
rect 132222 317056 132278 317112
rect 133786 496848 133842 496904
rect 136546 496848 136602 496904
rect 139306 496848 139362 496904
rect 142066 496848 142122 496904
rect 143446 496848 143502 496904
rect 148966 496848 149022 496904
rect 157246 496848 157302 496904
rect 168286 195336 168342 195392
rect 167366 195200 167422 195256
rect 168102 145560 168158 145616
rect 167366 136584 167422 136640
rect 166906 117816 166962 117872
rect 166998 96464 167054 96520
rect 167734 139576 167790 139632
rect 167642 111288 167698 111344
rect 167734 106392 167790 106448
rect 167826 98232 167882 98288
rect 168102 139440 168158 139496
rect 167918 89936 167974 89992
rect 168010 88304 168066 88360
rect 168286 139848 168342 139904
rect 168194 134272 168250 134328
rect 168838 126112 168894 126168
rect 168930 124480 168986 124536
rect 169206 119584 169262 119640
rect 169114 116184 169170 116240
rect 168286 114552 168342 114608
rect 169298 112920 169354 112976
rect 169482 139576 169538 139632
rect 169390 109656 169446 109712
rect 169482 108024 169538 108080
rect 169574 101496 169630 101552
rect 169850 139168 169906 139224
rect 169758 131008 169814 131064
rect 169666 99864 169722 99920
rect 170310 139712 170366 139768
rect 170310 135632 170366 135688
rect 170218 133184 170274 133240
rect 170126 104896 170182 104952
rect 170034 103264 170090 103320
rect 169942 95104 169998 95160
rect 168194 86672 168250 86728
rect 168102 83408 168158 83464
rect 168102 81776 168158 81832
rect 167458 80144 167514 80200
rect 168010 75248 168066 75304
rect 167274 73480 167330 73536
rect 167182 43968 167238 44024
rect 78678 28872 78734 28928
rect 167642 71848 167698 71904
rect 167734 68584 167790 68640
rect 167366 53896 167422 53952
rect 167550 48864 167606 48920
rect 167458 47232 167514 47288
rect 167918 70216 167974 70272
rect 167826 41792 167882 41848
rect 168194 76880 168250 76936
rect 169758 66952 169814 67008
rect 168286 65320 168342 65376
rect 169666 62056 169722 62112
rect 169482 58792 169538 58848
rect 169390 52128 169446 52184
rect 168286 41384 168342 41440
rect 168010 39072 168066 39128
rect 168286 39888 168342 39944
rect 168286 37440 168342 37496
rect 168286 35264 168342 35320
rect 169574 55528 169630 55584
rect 169850 50496 169906 50552
rect 169942 45736 169998 45792
rect 170586 33632 170642 33688
rect 170494 32000 170550 32056
rect 170402 31048 170458 31104
rect 170586 30232 170642 30288
rect 170494 29688 170550 29744
rect 181442 198600 181498 198656
rect 180062 198464 180118 198520
rect 186318 418376 186374 418432
rect 186318 415248 186374 415304
rect 186870 413072 186926 413128
rect 186318 412120 186374 412176
rect 186318 411032 186374 411088
rect 186410 409944 186466 410000
rect 186318 406816 186374 406872
rect 186318 403688 186374 403744
rect 186318 401548 186320 401568
rect 186320 401548 186372 401568
rect 186372 401548 186374 401568
rect 186318 401512 186374 401548
rect 186318 395256 186374 395312
rect 186318 393080 186374 393136
rect 186318 391040 186374 391096
rect 186318 388864 186374 388920
rect 186410 387912 186466 387968
rect 186318 385736 186374 385792
rect 186410 379480 186466 379536
rect 186318 378392 186374 378448
rect 186318 377304 186374 377360
rect 186318 376216 186374 376272
rect 186410 375284 186466 375320
rect 186410 375264 186412 375284
rect 186412 375264 186464 375284
rect 186464 375264 186466 375284
rect 186318 374176 186374 374232
rect 186318 373088 186374 373144
rect 186318 372000 186374 372056
rect 186318 371048 186374 371104
rect 186410 369960 186466 370016
rect 186318 368872 186374 368928
rect 186318 367784 186374 367840
rect 186318 366832 186374 366888
rect 186410 365744 186466 365800
rect 186318 364656 186374 364712
rect 186318 363568 186374 363624
rect 186318 362616 186374 362672
rect 186318 361548 186374 361584
rect 186318 361528 186320 361548
rect 186320 361528 186372 361548
rect 186372 361528 186374 361548
rect 186410 360440 186466 360496
rect 186318 359352 186374 359408
rect 186318 357348 186320 357368
rect 186320 357348 186372 357368
rect 186372 357348 186374 357368
rect 186318 357312 186374 357348
rect 186410 356224 186466 356280
rect 186318 355272 186374 355328
rect 186318 354184 186374 354240
rect 186410 353132 186412 353152
rect 186412 353132 186464 353152
rect 186464 353132 186466 353152
rect 186410 353096 186466 353132
rect 186318 352008 186374 352064
rect 186318 351056 186374 351112
rect 186318 349968 186374 350024
rect 186410 348880 186466 348936
rect 186318 347792 186374 347848
rect 186318 346840 186374 346896
rect 186318 345752 186374 345808
rect 186318 344664 186374 344720
rect 186318 343596 186374 343632
rect 186318 343576 186320 343596
rect 186320 343576 186372 343596
rect 186372 343576 186374 343596
rect 186410 342624 186466 342680
rect 186318 341536 186374 341592
rect 186318 340448 186374 340504
rect 186318 339396 186320 339416
rect 186320 339396 186372 339416
rect 186372 339396 186374 339416
rect 186318 339360 186374 339396
rect 186410 338408 186466 338464
rect 186318 337320 186374 337376
rect 186318 336232 186374 336288
rect 186318 335144 186374 335200
rect 186410 334192 186466 334248
rect 186318 333104 186374 333160
rect 186318 332016 186374 332072
rect 186318 330928 186374 330984
rect 186410 329976 186466 330032
rect 186318 328888 186374 328944
rect 186318 327800 186374 327856
rect 186318 326712 186374 326768
rect 186410 325760 186466 325816
rect 186318 324672 186374 324728
rect 186318 323584 186374 323640
rect 186318 322632 186374 322688
rect 186410 321544 186466 321600
rect 186318 320456 186374 320512
rect 186318 319368 186374 319424
rect 186318 318416 186374 318472
rect 186410 317348 186466 317384
rect 186410 317328 186412 317348
rect 186412 317328 186464 317348
rect 186464 317328 186466 317348
rect 186318 316240 186374 316296
rect 186318 315152 186374 315208
rect 186318 314200 186374 314256
rect 186318 313148 186320 313168
rect 186320 313148 186372 313168
rect 186372 313148 186374 313168
rect 186318 313112 186374 313148
rect 186410 312024 186466 312080
rect 186318 310936 186374 310992
rect 186318 309984 186374 310040
rect 186318 308896 186374 308952
rect 186410 307808 186466 307864
rect 186318 306720 186374 306776
rect 186318 305768 186374 305824
rect 186686 304680 186742 304736
rect 186410 303592 186466 303648
rect 186318 302504 186374 302560
rect 186318 301552 186374 301608
rect 186318 300464 186374 300520
rect 186318 299412 186320 299432
rect 186320 299412 186372 299432
rect 186372 299412 186374 299432
rect 186318 299376 186374 299412
rect 186410 298288 186466 298344
rect 186318 297336 186374 297392
rect 186318 296248 186374 296304
rect 186318 295160 186374 295216
rect 186410 294208 186466 294264
rect 186318 293120 186374 293176
rect 186318 292032 186374 292088
rect 186318 290944 186374 291000
rect 186410 289992 186466 290048
rect 186318 288904 186374 288960
rect 186318 287816 186374 287872
rect 186318 286728 186374 286784
rect 186410 285776 186466 285832
rect 186318 284688 186374 284744
rect 186318 283600 186374 283656
rect 186318 282512 186374 282568
rect 186410 281560 186466 281616
rect 186318 280472 186374 280528
rect 186318 279384 186374 279440
rect 186318 278296 186374 278352
rect 186318 277364 186374 277400
rect 186318 277344 186320 277364
rect 186320 277344 186372 277364
rect 186372 277344 186374 277364
rect 186410 276256 186466 276312
rect 186318 275168 186374 275224
rect 186318 274080 186374 274136
rect 186318 273164 186320 273184
rect 186320 273164 186372 273184
rect 186372 273164 186374 273184
rect 186318 273128 186374 273164
rect 186410 272040 186466 272096
rect 186318 270952 186374 271008
rect 186318 269864 186374 269920
rect 186410 268948 186412 268968
rect 186412 268948 186464 268968
rect 186464 268948 186466 268968
rect 186410 268912 186466 268948
rect 186318 267824 186374 267880
rect 186318 266736 186374 266792
rect 186318 265648 186374 265704
rect 186318 264696 186374 264752
rect 186410 263608 186466 263664
rect 186318 262520 186374 262576
rect 186318 261568 186374 261624
rect 186318 260480 186374 260536
rect 186410 259392 186466 259448
rect 186318 258304 186374 258360
rect 186318 257352 186374 257408
rect 186318 256264 186374 256320
rect 186318 255212 186320 255232
rect 186320 255212 186372 255232
rect 186372 255212 186374 255232
rect 186318 255176 186374 255212
rect 186410 254088 186466 254144
rect 186318 253136 186374 253192
rect 186318 252048 186374 252104
rect 186318 250960 186374 251016
rect 186410 249872 186466 249928
rect 186318 248920 186374 248976
rect 186318 247832 186374 247888
rect 186318 246744 186374 246800
rect 186410 245656 186466 245712
rect 186318 244704 186374 244760
rect 186318 243616 186374 243672
rect 186318 242528 186374 242584
rect 186318 241440 186374 241496
rect 186410 240488 186466 240544
rect 186318 239400 186374 239456
rect 186318 238312 186374 238368
rect 186318 237224 186374 237280
rect 186410 236272 186466 236328
rect 186318 235184 186374 235240
rect 186318 234096 186374 234152
rect 186318 233008 186374 233064
rect 186410 232056 186466 232112
rect 186318 230968 186374 231024
rect 186318 229880 186374 229936
rect 186318 228928 186374 228984
rect 186410 227840 186466 227896
rect 186318 226752 186374 226808
rect 186318 225664 186374 225720
rect 186318 224712 186374 224768
rect 186410 223624 186466 223680
rect 186318 222536 186374 222592
rect 186318 221448 186374 221504
rect 186502 220496 186558 220552
rect 186410 219408 186466 219464
rect 186318 218320 186374 218376
rect 186318 217232 186374 217288
rect 186318 216280 186374 216336
rect 186318 215212 186374 215248
rect 186318 215192 186320 215212
rect 186320 215192 186372 215212
rect 186372 215192 186374 215212
rect 186410 214104 186466 214160
rect 186318 213016 186374 213072
rect 186318 212064 186374 212120
rect 186318 210976 186374 211032
rect 186410 209888 186466 209944
rect 186318 208800 186374 208856
rect 186318 207848 186374 207904
rect 186410 206760 186466 206816
rect 186318 205672 186374 205728
rect 186318 204584 186374 204640
rect 186318 203632 186374 203688
rect 186318 202544 186374 202600
rect 186410 201456 186466 201512
rect 186318 200504 186374 200560
rect 187054 402600 187110 402656
rect 187606 416336 187662 416392
rect 187514 414160 187570 414216
rect 187146 394168 187202 394224
rect 187330 396208 187386 396264
rect 187238 389952 187294 390008
rect 187330 386824 187386 386880
rect 187238 381520 187294 381576
rect 187146 380432 187202 380488
rect 187514 407904 187570 407960
rect 187514 400424 187570 400480
rect 187422 384648 187478 384704
rect 187422 358400 187478 358456
rect 188802 405728 188858 405784
rect 188710 404640 188766 404696
rect 188986 397296 189042 397352
rect 189170 408856 189226 408912
rect 189078 391992 189134 392048
rect 189078 382608 189134 382664
rect 189262 399472 189318 399528
rect 189354 398384 189410 398440
rect 190734 420044 190736 420064
rect 190736 420044 190788 420064
rect 190788 420044 190790 420064
rect 190734 420008 190790 420044
rect 396630 535880 396686 535936
rect 396722 533704 396778 533760
rect 396630 532772 396686 532808
rect 396630 532752 396632 532772
rect 396632 532752 396684 532772
rect 396684 532752 396686 532772
rect 396722 530984 396778 531040
rect 396630 529932 396632 529952
rect 396632 529932 396684 529952
rect 396684 529932 396686 529952
rect 396630 529896 396686 529932
rect 396630 528128 396686 528184
rect 396354 509904 396410 509960
rect 397366 508272 397422 508328
rect 396630 508000 396686 508056
rect 351090 420144 351146 420200
rect 370870 422320 370926 422376
rect 380898 420960 380954 421016
rect 419630 498072 419686 498128
rect 433522 498072 433578 498128
rect 440238 498072 440294 498128
rect 454682 498072 454738 498128
rect 455786 498072 455842 498128
rect 400678 420960 400734 421016
rect 190366 417832 190422 417888
rect 409326 413072 409382 413128
rect 252190 197920 252246 197976
rect 260838 192480 260894 192536
rect 191470 28736 191526 28792
rect 199842 28600 199898 28656
rect 233790 28464 233846 28520
rect 242254 28328 242310 28384
rect 279330 29688 279386 29744
rect 281538 133592 281594 133648
rect 280250 92384 280306 92440
rect 282182 78512 282238 78568
rect 282458 119856 282514 119912
rect 282366 106120 282422 106176
rect 282274 64640 282330 64696
rect 280158 37168 280214 37224
rect 280802 29960 280858 30016
rect 280986 29824 281042 29880
rect 282826 50768 282882 50824
rect 292118 198056 292174 198112
rect 360106 198328 360162 198384
rect 387798 198464 387854 198520
rect 392582 139984 392638 140040
rect 392766 139848 392822 139904
rect 393134 59200 393190 59256
rect 395250 195472 395306 195528
rect 394422 63416 394478 63472
rect 395250 139712 395306 139768
rect 393962 30096 394018 30152
rect 396814 96464 396870 96520
rect 396998 53896 397054 53952
rect 397182 43968 397238 44024
rect 397918 139440 397974 139496
rect 397826 135904 397882 135960
rect 397458 134272 397514 134328
rect 397458 132640 397514 132696
rect 397458 129376 397514 129432
rect 397458 124480 397514 124536
rect 397458 122848 397514 122904
rect 397458 119584 397514 119640
rect 397826 116184 397882 116240
rect 398102 117816 398158 117872
rect 398010 114552 398066 114608
rect 397550 112920 397606 112976
rect 397458 104796 397460 104816
rect 397460 104796 397512 104816
rect 397512 104796 397514 104816
rect 397458 104760 397514 104796
rect 397458 101496 397514 101552
rect 397458 98232 397514 98288
rect 397458 94832 397514 94888
rect 398194 109656 398250 109712
rect 398102 93200 398158 93256
rect 397458 91568 397514 91624
rect 397918 89936 397974 89992
rect 397458 88304 397514 88360
rect 397734 86672 397790 86728
rect 397550 85040 397606 85096
rect 397458 81776 397514 81832
rect 398194 80144 398250 80200
rect 397458 78548 397460 78568
rect 397460 78548 397512 78568
rect 397512 78548 397514 78568
rect 397458 78512 397514 78548
rect 398010 76880 398066 76936
rect 398102 75268 398158 75304
rect 398102 75248 398104 75268
rect 398104 75248 398156 75268
rect 398156 75248 398158 75268
rect 397918 71868 397974 71904
rect 397918 71848 397920 71868
rect 397920 71848 397972 71868
rect 397972 71848 397974 71868
rect 397458 66952 397514 67008
rect 397458 60424 397514 60480
rect 397458 59200 397514 59256
rect 397458 57196 397460 57216
rect 397460 57196 397512 57216
rect 397512 57196 397514 57216
rect 397458 57160 397514 57196
rect 397918 50496 397974 50552
rect 397458 48864 397514 48920
rect 397458 47232 397514 47288
rect 397458 42336 397514 42392
rect 397458 40724 397514 40760
rect 397458 40704 397460 40724
rect 397460 40704 397512 40724
rect 397512 40704 397514 40724
rect 397458 39072 397514 39128
rect 397550 37440 397606 37496
rect 397458 34176 397514 34232
rect 397366 33088 397422 33144
rect 397458 32544 397514 32600
rect 397458 30912 397514 30968
rect 398194 73480 398250 73536
rect 398930 199416 398986 199472
rect 398378 131008 398434 131064
rect 398378 99864 398434 99920
rect 398286 71848 398342 71904
rect 398286 70216 398342 70272
rect 398378 68584 398434 68640
rect 398470 65320 398526 65376
rect 398562 58792 398618 58848
rect 398654 52128 398710 52184
rect 398838 111288 398894 111344
rect 398838 76880 398894 76936
rect 398746 47232 398802 47288
rect 398746 45600 398802 45656
rect 399482 144064 399538 144120
rect 399206 68584 399262 68640
rect 399206 62056 399262 62112
rect 399114 55528 399170 55584
rect 398838 42336 398894 42392
rect 399574 127744 399630 127800
rect 399574 83408 399630 83464
rect 399482 62056 399538 62112
rect 399390 50496 399446 50552
rect 399298 37440 399354 37496
rect 400126 142704 400182 142760
rect 400586 126656 400642 126712
rect 400586 121388 400588 121408
rect 400588 121388 400640 121408
rect 400640 121388 400642 121408
rect 400586 121352 400642 121388
rect 400218 103264 400274 103320
rect 403530 198600 403586 198656
rect 404358 196016 404414 196072
rect 409326 410216 409382 410272
rect 409326 404368 409382 404424
rect 409418 398792 409474 398848
rect 415398 496848 415454 496904
rect 416778 496848 416834 496904
rect 418158 496848 418214 496904
rect 419538 496848 419594 496904
rect 409878 355816 409934 355872
rect 410246 369552 410302 369608
rect 410154 363432 410210 363488
rect 410062 333104 410118 333160
rect 409970 320864 410026 320920
rect 409878 307672 409934 307728
rect 409418 236136 409474 236192
rect 409234 196560 409290 196616
rect 409510 227840 409566 227896
rect 409970 305360 410026 305416
rect 410154 299648 410210 299704
rect 410154 295568 410210 295624
rect 410246 252456 410302 252512
rect 410430 394304 410486 394360
rect 410430 392264 410486 392320
rect 410338 224984 410394 225040
rect 410338 221584 410394 221640
rect 410706 414840 410762 414896
rect 410614 400424 410670 400480
rect 410522 373768 410578 373824
rect 411258 371728 411314 371784
rect 411258 365472 411314 365528
rect 411258 359372 411314 359408
rect 411258 359352 411260 359372
rect 411260 359352 411312 359372
rect 411312 359352 411314 359372
rect 411350 357312 411406 357368
rect 411258 353132 411260 353152
rect 411260 353132 411312 353152
rect 411312 353132 411314 353152
rect 411258 353096 411314 353132
rect 410614 349016 410670 349072
rect 410522 307944 410578 308000
rect 410522 299648 410578 299704
rect 410522 244160 410578 244216
rect 411442 346976 411498 347032
rect 411258 344936 411314 344992
rect 411258 342896 411314 342952
rect 411442 340856 411498 340912
rect 410706 338816 410762 338872
rect 411258 336776 411314 336832
rect 411258 330520 411314 330576
rect 411258 326440 411314 326496
rect 411258 324400 411314 324456
rect 411258 318144 411314 318200
rect 411258 316104 411314 316160
rect 411258 314064 411314 314120
rect 411258 312024 411314 312080
rect 411258 309984 411314 310040
rect 411258 303864 411314 303920
rect 411258 297608 411314 297664
rect 411258 293528 411314 293584
rect 411258 291488 411314 291544
rect 411258 289448 411314 289504
rect 411258 287408 411314 287464
rect 411258 285232 411314 285288
rect 411258 283192 411314 283248
rect 411258 281152 411314 281208
rect 411258 279112 411314 279168
rect 411258 277072 411314 277128
rect 411258 275032 411314 275088
rect 411258 272992 411314 273048
rect 411258 270952 411314 271008
rect 411258 268912 411314 268968
rect 411258 266736 411314 266792
rect 411258 264696 411314 264752
rect 411258 262656 411314 262712
rect 411258 260616 411314 260672
rect 411258 258576 411314 258632
rect 411258 256536 411314 256592
rect 411258 254532 411260 254552
rect 411260 254532 411312 254552
rect 411312 254532 411314 254552
rect 411258 254496 411314 254532
rect 410798 252492 410800 252512
rect 410800 252492 410852 252512
rect 410852 252492 410854 252512
rect 410798 252456 410854 252492
rect 411258 250280 411314 250336
rect 411258 246200 411314 246256
rect 410798 244196 410800 244216
rect 410800 244196 410852 244216
rect 410852 244196 410854 244216
rect 410798 244160 410854 244196
rect 411258 242120 411314 242176
rect 411258 240100 411314 240136
rect 411258 240080 411260 240100
rect 411260 240080 411312 240100
rect 411312 240080 411314 240100
rect 411258 238040 411314 238096
rect 411258 233824 411314 233880
rect 411350 231784 411406 231840
rect 411258 229744 411314 229800
rect 411258 223644 411314 223680
rect 411258 223624 411260 223644
rect 411260 223624 411312 223644
rect 411312 223624 411314 223644
rect 410798 221584 410854 221640
rect 411258 217368 411314 217424
rect 411258 213324 411260 213344
rect 411260 213324 411312 213344
rect 411312 213324 411314 213344
rect 411258 213288 411314 213324
rect 411258 211248 411314 211304
rect 411350 207168 411406 207224
rect 411258 205128 411314 205184
rect 411258 203108 411314 203144
rect 411258 203088 411260 203108
rect 411260 203088 411312 203108
rect 411312 203088 411314 203108
rect 411258 201048 411314 201104
rect 432142 497120 432198 497176
rect 426438 496984 426494 497040
rect 427910 496984 427966 497040
rect 430578 496984 430634 497040
rect 420918 496848 420974 496904
rect 422298 496848 422354 496904
rect 423678 496848 423734 496904
rect 425058 496848 425114 496904
rect 426530 496868 426586 496904
rect 426530 496848 426532 496868
rect 426532 496848 426584 496868
rect 426584 496848 426586 496868
rect 427818 496848 427874 496904
rect 433430 496984 433486 497040
rect 429198 496848 429254 496904
rect 430670 496848 430726 496904
rect 433338 496868 433394 496904
rect 433338 496848 433340 496868
rect 433340 496848 433392 496868
rect 433392 496848 433394 496868
rect 434718 496984 434774 497040
rect 437478 496984 437534 497040
rect 434810 496848 434866 496904
rect 436098 496848 436154 496904
rect 437570 496848 437626 496904
rect 438858 496848 438914 496904
rect 441618 496984 441674 497040
rect 443090 496984 443146 497040
rect 445850 496984 445906 497040
rect 447138 496984 447194 497040
rect 448610 496984 448666 497040
rect 449990 496984 450046 497040
rect 452658 496984 452714 497040
rect 440330 496848 440386 496904
rect 441710 496848 441766 496904
rect 442998 496848 443054 496904
rect 444378 496848 444434 496904
rect 445942 496848 445998 496904
rect 412086 418940 412142 418976
rect 412086 418920 412088 418940
rect 412088 418920 412140 418940
rect 412140 418920 412142 418940
rect 412086 416900 412142 416936
rect 412086 416880 412088 416900
rect 412088 416880 412140 416900
rect 412140 416880 412142 416900
rect 411994 396344 412050 396400
rect 411994 390260 411996 390280
rect 411996 390260 412048 390280
rect 412048 390260 412050 390280
rect 411994 390224 412050 390260
rect 411902 388184 411958 388240
rect 411810 386008 411866 386064
rect 411810 383968 411866 384024
rect 411718 381928 411774 381984
rect 412178 379888 412234 379944
rect 411810 375808 411866 375864
rect 411626 351056 411682 351112
rect 411534 322360 411590 322416
rect 411534 301688 411590 301744
rect 411534 225664 411590 225720
rect 410706 193976 410762 194032
rect 410614 193840 410670 193896
rect 411626 209208 411682 209264
rect 411810 248240 411866 248296
rect 411994 219544 412050 219600
rect 412086 215328 412142 215384
rect 412270 367512 412326 367568
rect 412546 361392 412602 361448
rect 412822 334600 412878 334656
rect 416962 195472 417018 195528
rect 417514 198328 417570 198384
rect 413834 139984 413890 140040
rect 437478 409128 437534 409184
rect 437478 407496 437534 407552
rect 437478 405864 437534 405920
rect 437478 404268 437480 404288
rect 437480 404268 437532 404288
rect 437532 404268 437534 404288
rect 437478 404232 437534 404268
rect 437478 402600 437534 402656
rect 437478 400968 437534 401024
rect 437478 399336 437534 399392
rect 437570 397704 437626 397760
rect 436742 396072 436798 396128
rect 437570 394440 437626 394496
rect 437478 392808 437534 392864
rect 437478 391176 437534 391232
rect 437754 389544 437810 389600
rect 437478 384512 437534 384568
rect 437938 382880 437994 382936
rect 437478 381248 437534 381304
rect 437478 379616 437534 379672
rect 437478 377984 437534 378040
rect 437478 376352 437534 376408
rect 437478 374720 437534 374776
rect 437018 373088 437074 373144
rect 436926 359896 436982 359952
rect 436834 304136 436890 304192
rect 437478 371456 437534 371512
rect 437478 369860 437480 369880
rect 437480 369860 437532 369880
rect 437532 369860 437534 369880
rect 437478 369824 437534 369860
rect 437478 368192 437534 368248
rect 437478 366424 437534 366480
rect 437478 364792 437534 364848
rect 437478 363160 437534 363216
rect 437478 361528 437534 361584
rect 437478 358264 437534 358320
rect 437478 356632 437534 356688
rect 437478 355000 437534 355056
rect 437478 353368 437534 353424
rect 437478 351736 437534 351792
rect 437478 350104 437534 350160
rect 437478 348472 437534 348528
rect 437478 346840 437534 346896
rect 437478 345208 437534 345264
rect 437478 343440 437534 343496
rect 437846 340176 437902 340232
rect 437478 338544 437534 338600
rect 437478 336912 437534 336968
rect 437570 335280 437626 335336
rect 437478 333648 437534 333704
rect 437478 332016 437534 332072
rect 437478 330384 437534 330440
rect 437478 328752 437534 328808
rect 437478 327120 437534 327176
rect 437478 318844 437534 318880
rect 437478 318824 437480 318844
rect 437480 318824 437532 318844
rect 437532 318824 437534 318844
rect 437478 315560 437534 315616
rect 437478 313928 437534 313984
rect 438030 312296 438086 312352
rect 437478 310664 437534 310720
rect 437478 309032 437534 309088
rect 437570 307400 437626 307456
rect 437478 305768 437534 305824
rect 447230 496848 447286 496904
rect 448518 496848 448574 496904
rect 449898 496848 449954 496904
rect 451278 496848 451334 496904
rect 452750 496848 452806 496904
rect 454038 496848 454094 496904
rect 462318 498092 462374 498128
rect 462318 498072 462320 498092
rect 462320 498072 462372 498092
rect 462372 498072 462374 498092
rect 456798 497256 456854 497312
rect 456890 496848 456946 496904
rect 458270 496984 458326 497040
rect 498198 496984 498254 497040
rect 458178 496848 458234 496904
rect 460938 496848 460994 496904
rect 465078 496848 465134 496904
rect 467838 496848 467894 496904
rect 470598 496848 470654 496904
rect 473358 496848 473414 496904
rect 474738 496848 474794 496904
rect 477498 496848 477554 496904
rect 480258 496848 480314 496904
rect 483018 496848 483074 496904
rect 485778 496848 485834 496904
rect 488538 496848 488594 496904
rect 489918 496848 489974 496904
rect 492678 496848 492734 496904
rect 495438 496868 495494 496904
rect 495438 496848 495440 496868
rect 495440 496848 495492 496868
rect 495492 496848 495494 496868
rect 500958 496848 501014 496904
rect 502338 496848 502394 496904
rect 505098 496868 505154 496904
rect 505098 496848 505100 496868
rect 505100 496848 505152 496868
rect 505152 496848 505154 496868
rect 580170 431568 580226 431624
rect 438306 387776 438362 387832
rect 438398 386144 438454 386200
rect 438490 341808 438546 341864
rect 438766 325488 438822 325544
rect 438582 323856 438638 323912
rect 438490 322088 438546 322144
rect 438398 320456 438454 320512
rect 438306 302504 438362 302560
rect 438398 300872 438454 300928
rect 438674 317192 438730 317248
rect 510802 198056 510858 198112
rect 510618 197920 510674 197976
rect 491298 142704 491354 142760
rect 400586 70352 400642 70408
rect 399758 35808 399814 35864
rect 454682 28872 454738 28928
rect 510618 78512 510674 78568
rect 509514 37204 509516 37224
rect 509516 37204 509568 37224
rect 509568 37204 509570 37224
rect 509514 37168 509570 37204
rect 510802 106120 510858 106176
rect 512182 133592 512238 133648
rect 512090 119856 512146 119912
rect 511998 92384 512054 92440
rect 510894 64640 510950 64696
rect 512274 50904 512330 50960
rect 550638 403008 550694 403064
rect 550546 306448 550602 306504
rect 552018 361800 552074 361856
rect 552018 334328 552074 334384
rect 552294 389272 552350 389328
rect 552202 375536 552258 375592
rect 552202 348064 552258 348120
rect 552110 320592 552166 320648
rect 551374 28600 551430 28656
rect 556802 28736 556858 28792
rect 580170 418240 580226 418296
rect 580170 378392 580226 378448
rect 580170 365064 580226 365120
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 579802 272176 579858 272232
rect 580170 258848 580226 258904
rect 579802 245520 579858 245576
rect 579986 232328 580042 232384
rect 580170 219000 580226 219056
rect 580170 205692 580226 205728
rect 580170 205672 580172 205692
rect 580172 205672 580224 205692
rect 580224 205672 580226 205692
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 152632 580226 152688
rect 579710 125976 579766 126032
rect 579710 112784 579766 112840
rect 579986 86128 580042 86184
rect 580170 46280 580226 46336
rect 580630 139304 580686 139360
rect 580538 99456 580594 99512
rect 580446 72936 580502 72992
rect 580354 59608 580410 59664
rect 580262 19760 580318 19816
rect 580170 6568 580226 6624
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect 48037 536890 48103 536893
rect 49374 536890 50048 536924
rect 48037 536888 50048 536890
rect 48037 536832 48042 536888
rect 48098 536864 50048 536888
rect 396625 536890 396691 536893
rect 399342 536890 400016 536924
rect 396625 536888 400016 536890
rect 48098 536832 49434 536864
rect 48037 536830 49434 536832
rect 396625 536832 396630 536888
rect 396686 536864 400016 536888
rect 396686 536832 399402 536864
rect 396625 536830 399402 536832
rect 48037 536827 48103 536830
rect 396625 536827 396691 536830
rect 48221 535938 48287 535941
rect 49374 535938 50048 535972
rect 48221 535936 50048 535938
rect 48221 535880 48226 535936
rect 48282 535912 50048 535936
rect 396625 535938 396691 535941
rect 399342 535938 400016 535972
rect 396625 535936 400016 535938
rect 48282 535880 49434 535912
rect 48221 535878 49434 535880
rect 396625 535880 396630 535936
rect 396686 535912 400016 535936
rect 396686 535880 399402 535912
rect 396625 535878 399402 535880
rect 48221 535875 48287 535878
rect 396625 535875 396691 535878
rect 47945 533762 48011 533765
rect 49374 533762 50048 533796
rect 47945 533760 50048 533762
rect 47945 533704 47950 533760
rect 48006 533736 50048 533760
rect 396717 533762 396783 533765
rect 399342 533762 400016 533796
rect 396717 533760 400016 533762
rect 48006 533704 49434 533736
rect 47945 533702 49434 533704
rect 396717 533704 396722 533760
rect 396778 533736 400016 533760
rect 396778 533704 399402 533736
rect 396717 533702 399402 533704
rect 47945 533699 48011 533702
rect 396717 533699 396783 533702
rect 48129 532810 48195 532813
rect 49374 532810 50048 532844
rect 48129 532808 50048 532810
rect 48129 532752 48134 532808
rect 48190 532784 50048 532808
rect 396625 532810 396691 532813
rect 399342 532810 400016 532844
rect 396625 532808 400016 532810
rect 48190 532752 49434 532784
rect 48129 532750 49434 532752
rect 396625 532752 396630 532808
rect 396686 532784 400016 532808
rect 396686 532752 399402 532784
rect 396625 532750 399402 532752
rect 48129 532747 48195 532750
rect 396625 532747 396691 532750
rect 47853 531042 47919 531045
rect 49374 531042 50048 531076
rect 47853 531040 50048 531042
rect 47853 530984 47858 531040
rect 47914 531016 50048 531040
rect 396717 531042 396783 531045
rect 399342 531042 400016 531076
rect 396717 531040 400016 531042
rect 47914 530984 49434 531016
rect 47853 530982 49434 530984
rect 396717 530984 396722 531040
rect 396778 531016 400016 531040
rect 396778 530984 399402 531016
rect 396717 530982 399402 530984
rect 47853 530979 47919 530982
rect 396717 530979 396783 530982
rect 49509 529988 49575 529991
rect 49509 529986 50048 529988
rect 49509 529930 49514 529986
rect 49570 529930 50048 529986
rect 49509 529928 50048 529930
rect 396625 529954 396691 529957
rect 399342 529954 400016 529988
rect 396625 529952 400016 529954
rect 49509 529925 49575 529928
rect 396625 529896 396630 529952
rect 396686 529928 400016 529952
rect 396686 529896 399402 529928
rect 396625 529894 399402 529896
rect 396625 529891 396691 529894
rect 49417 528220 49483 528223
rect 49417 528218 50048 528220
rect 49417 528162 49422 528218
rect 49478 528162 50048 528218
rect 49417 528160 50048 528162
rect 396625 528186 396691 528189
rect 399342 528186 400016 528220
rect 396625 528184 400016 528186
rect 49417 528157 49483 528160
rect 396625 528128 396630 528184
rect 396686 528160 400016 528184
rect 396686 528128 399402 528160
rect 396625 528126 399402 528128
rect 396625 528123 396691 528126
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect 49601 509996 49667 509999
rect 49601 509994 50048 509996
rect 49601 509938 49606 509994
rect 49662 509938 50048 509994
rect 49601 509936 50048 509938
rect 396349 509962 396415 509965
rect 399342 509962 400016 509996
rect 396349 509960 400016 509962
rect 49601 509933 49667 509936
rect 396349 509904 396354 509960
rect 396410 509936 400016 509960
rect 396410 509904 399402 509936
rect 396349 509902 399402 509904
rect 396349 509899 396415 509902
rect 49325 508330 49391 508333
rect 49742 508330 50048 508364
rect 49325 508328 50048 508330
rect 49325 508272 49330 508328
rect 49386 508304 50048 508328
rect 397361 508330 397427 508333
rect 399342 508330 400016 508364
rect 397361 508328 400016 508330
rect 49386 508272 49802 508304
rect 49325 508270 49802 508272
rect 397361 508272 397366 508328
rect 397422 508304 400016 508328
rect 397422 508272 399402 508304
rect 397361 508270 399402 508272
rect 49325 508267 49391 508270
rect 397361 508267 397427 508270
rect 47761 508058 47827 508061
rect 49374 508058 50048 508092
rect 47761 508056 50048 508058
rect 47761 508000 47766 508056
rect 47822 508032 50048 508056
rect 396625 508058 396691 508061
rect 399342 508058 400016 508092
rect 396625 508056 400016 508058
rect 47822 508000 49434 508032
rect 47761 507998 49434 508000
rect 396625 508000 396630 508056
rect 396686 508032 400016 508056
rect 396686 508000 399402 508032
rect 396625 507998 399402 508000
rect 47761 507995 47827 507998
rect 396625 507995 396691 507998
rect -960 501652 480 501892
rect 435766 499700 435772 499764
rect 435836 499762 435842 499764
rect 436040 499762 436046 499764
rect 435836 499702 436046 499762
rect 435836 499700 435842 499702
rect 436040 499700 436046 499702
rect 436110 499700 436116 499764
rect 67214 498204 67220 498268
rect 67284 498204 67290 498268
rect 74206 498204 74212 498268
rect 74276 498204 74282 498268
rect 77702 498204 77708 498268
rect 77772 498204 77778 498268
rect 91870 498204 91876 498268
rect 91940 498204 91946 498268
rect 95918 498204 95924 498268
rect 95988 498204 95994 498268
rect 103278 498204 103284 498268
rect 103348 498204 103354 498268
rect 120942 498204 120948 498268
rect 121012 498204 121018 498268
rect 145966 498204 145972 498268
rect 146036 498204 146042 498268
rect 153326 498204 153332 498268
rect 153396 498204 153402 498268
rect 419574 498204 419580 498268
rect 419644 498204 419650 498268
rect 455638 498204 455644 498268
rect 455708 498204 455714 498268
rect 463550 498204 463556 498268
rect 463620 498204 463626 498268
rect 67222 498130 67282 498204
rect 67541 498130 67607 498133
rect 67222 498128 67607 498130
rect 67222 498072 67546 498128
rect 67602 498072 67607 498128
rect 67222 498070 67607 498072
rect 67541 498067 67607 498070
rect 73102 498068 73108 498132
rect 73172 498130 73178 498132
rect 73337 498130 73403 498133
rect 73172 498128 73403 498130
rect 73172 498072 73342 498128
rect 73398 498072 73403 498128
rect 73172 498070 73403 498072
rect 74214 498130 74274 498204
rect 74349 498130 74415 498133
rect 74214 498128 74415 498130
rect 74214 498072 74354 498128
rect 74410 498072 74415 498128
rect 74214 498070 74415 498072
rect 77710 498130 77770 498204
rect 78581 498130 78647 498133
rect 77710 498128 78647 498130
rect 77710 498072 78586 498128
rect 78642 498072 78647 498128
rect 77710 498070 78647 498072
rect 73172 498068 73178 498070
rect 73337 498067 73403 498070
rect 74349 498067 74415 498070
rect 78581 498067 78647 498070
rect 78806 498068 78812 498132
rect 78876 498130 78882 498132
rect 79869 498130 79935 498133
rect 78876 498128 79935 498130
rect 78876 498072 79874 498128
rect 79930 498072 79935 498128
rect 78876 498070 79935 498072
rect 78876 498068 78882 498070
rect 79869 498067 79935 498070
rect 80094 498068 80100 498132
rect 80164 498130 80170 498132
rect 81249 498130 81315 498133
rect 80164 498128 81315 498130
rect 80164 498072 81254 498128
rect 81310 498072 81315 498128
rect 80164 498070 81315 498072
rect 80164 498068 80170 498070
rect 81249 498067 81315 498070
rect 85798 498068 85804 498132
rect 85868 498130 85874 498132
rect 85941 498130 86007 498133
rect 85868 498128 86007 498130
rect 85868 498072 85946 498128
rect 86002 498072 86007 498128
rect 85868 498070 86007 498072
rect 85868 498068 85874 498070
rect 85941 498067 86007 498070
rect 86166 498068 86172 498132
rect 86236 498130 86242 498132
rect 86493 498130 86559 498133
rect 89529 498132 89595 498133
rect 89478 498130 89484 498132
rect 86236 498128 86559 498130
rect 86236 498072 86498 498128
rect 86554 498072 86559 498128
rect 86236 498070 86559 498072
rect 89438 498070 89484 498130
rect 89548 498128 89595 498132
rect 89590 498072 89595 498128
rect 86236 498068 86242 498070
rect 86493 498067 86559 498070
rect 89478 498068 89484 498070
rect 89548 498068 89595 498072
rect 91878 498130 91938 498204
rect 92289 498130 92355 498133
rect 91878 498128 92355 498130
rect 91878 498072 92294 498128
rect 92350 498072 92355 498128
rect 91878 498070 92355 498072
rect 95926 498130 95986 498204
rect 96521 498130 96587 498133
rect 95926 498128 96587 498130
rect 95926 498072 96526 498128
rect 96582 498072 96587 498128
rect 95926 498070 96587 498072
rect 103286 498130 103346 498204
rect 103421 498130 103487 498133
rect 103286 498128 103487 498130
rect 103286 498072 103426 498128
rect 103482 498072 103487 498128
rect 103286 498070 103487 498072
rect 89529 498067 89595 498068
rect 92289 498067 92355 498070
rect 96521 498067 96587 498070
rect 103421 498067 103487 498070
rect 103646 498068 103652 498132
rect 103716 498130 103722 498132
rect 104801 498130 104867 498133
rect 103716 498128 104867 498130
rect 103716 498072 104806 498128
rect 104862 498072 104867 498128
rect 103716 498070 104867 498072
rect 103716 498068 103722 498070
rect 104801 498067 104867 498070
rect 113398 498068 113404 498132
rect 113468 498130 113474 498132
rect 113541 498130 113607 498133
rect 113468 498128 113607 498130
rect 113468 498072 113546 498128
rect 113602 498072 113607 498128
rect 113468 498070 113607 498072
rect 113468 498068 113474 498070
rect 113541 498067 113607 498070
rect 115974 498068 115980 498132
rect 116044 498130 116050 498132
rect 116853 498130 116919 498133
rect 116044 498128 116919 498130
rect 116044 498072 116858 498128
rect 116914 498072 116919 498128
rect 116044 498070 116919 498072
rect 116044 498068 116050 498070
rect 116853 498067 116919 498070
rect 118366 498068 118372 498132
rect 118436 498130 118442 498132
rect 118601 498130 118667 498133
rect 118436 498128 118667 498130
rect 118436 498072 118606 498128
rect 118662 498072 118667 498128
rect 118436 498070 118667 498072
rect 120950 498130 121010 498204
rect 121361 498130 121427 498133
rect 120950 498128 121427 498130
rect 120950 498072 121366 498128
rect 121422 498072 121427 498128
rect 120950 498070 121427 498072
rect 118436 498068 118442 498070
rect 118601 498067 118667 498070
rect 121361 498067 121427 498070
rect 125910 498068 125916 498132
rect 125980 498130 125986 498132
rect 126881 498130 126947 498133
rect 125980 498128 126947 498130
rect 125980 498072 126886 498128
rect 126942 498072 126947 498128
rect 125980 498070 126947 498072
rect 125980 498068 125986 498070
rect 126881 498067 126947 498070
rect 128486 498068 128492 498132
rect 128556 498130 128562 498132
rect 129641 498130 129707 498133
rect 128556 498128 129707 498130
rect 128556 498072 129646 498128
rect 129702 498072 129707 498128
rect 128556 498070 129707 498072
rect 145974 498130 146034 498204
rect 146201 498130 146267 498133
rect 150985 498132 151051 498133
rect 150934 498130 150940 498132
rect 145974 498128 146267 498130
rect 145974 498072 146206 498128
rect 146262 498072 146267 498128
rect 145974 498070 146267 498072
rect 150894 498070 150940 498130
rect 151004 498128 151051 498132
rect 151046 498072 151051 498128
rect 128556 498068 128562 498070
rect 129641 498067 129707 498070
rect 146201 498067 146267 498070
rect 150934 498068 150940 498070
rect 151004 498068 151051 498072
rect 153334 498130 153394 498204
rect 419582 498133 419642 498204
rect 154481 498130 154547 498133
rect 153334 498128 154547 498130
rect 153334 498072 154486 498128
rect 154542 498072 154547 498128
rect 153334 498070 154547 498072
rect 419582 498128 419691 498133
rect 419582 498072 419630 498128
rect 419686 498072 419691 498128
rect 419582 498070 419691 498072
rect 150985 498067 151051 498068
rect 154481 498067 154547 498070
rect 419625 498067 419691 498070
rect 433517 498130 433583 498133
rect 434478 498130 434484 498132
rect 433517 498128 434484 498130
rect 433517 498072 433522 498128
rect 433578 498072 434484 498128
rect 433517 498070 434484 498072
rect 433517 498067 433583 498070
rect 434478 498068 434484 498070
rect 434548 498068 434554 498132
rect 440233 498130 440299 498133
rect 441102 498130 441108 498132
rect 440233 498128 441108 498130
rect 440233 498072 440238 498128
rect 440294 498072 441108 498128
rect 440233 498070 441108 498072
rect 440233 498067 440299 498070
rect 441102 498068 441108 498070
rect 441172 498068 441178 498132
rect 454677 498130 454743 498133
rect 455646 498130 455706 498204
rect 454677 498128 455706 498130
rect 454677 498072 454682 498128
rect 454738 498072 455706 498128
rect 454677 498070 455706 498072
rect 455781 498130 455847 498133
rect 456190 498130 456196 498132
rect 455781 498128 456196 498130
rect 455781 498072 455786 498128
rect 455842 498072 456196 498128
rect 455781 498070 456196 498072
rect 454677 498067 454743 498070
rect 455781 498067 455847 498070
rect 456190 498068 456196 498070
rect 456260 498068 456266 498132
rect 462313 498130 462379 498133
rect 463558 498130 463618 498204
rect 462313 498128 463618 498130
rect 462313 498072 462318 498128
rect 462374 498072 463618 498128
rect 462313 498070 463618 498072
rect 462313 498067 462379 498070
rect 96337 497860 96403 497861
rect 96286 497858 96292 497860
rect 96246 497798 96292 497858
rect 96356 497856 96403 497860
rect 96398 497800 96403 497856
rect 583520 497844 584960 498084
rect 96286 497796 96292 497798
rect 96356 497796 96403 497800
rect 96337 497795 96403 497796
rect 71814 497388 71820 497452
rect 71884 497450 71890 497452
rect 73061 497450 73127 497453
rect 71884 497448 73127 497450
rect 71884 497392 73066 497448
rect 73122 497392 73127 497448
rect 71884 497390 73127 497392
rect 71884 497388 71890 497390
rect 73061 497387 73127 497390
rect 456793 497314 456859 497317
rect 458030 497314 458036 497316
rect 456793 497312 458036 497314
rect 456793 497256 456798 497312
rect 456854 497256 458036 497312
rect 456793 497254 458036 497256
rect 456793 497251 456859 497254
rect 458030 497252 458036 497254
rect 458100 497252 458106 497316
rect 432137 497178 432203 497181
rect 432270 497178 432276 497180
rect 432137 497176 432276 497178
rect 432137 497120 432142 497176
rect 432198 497120 432276 497176
rect 432137 497118 432276 497120
rect 432137 497115 432203 497118
rect 432270 497116 432276 497118
rect 432340 497116 432346 497180
rect 80830 496980 80836 497044
rect 80900 497042 80906 497044
rect 81157 497042 81223 497045
rect 80900 497040 81223 497042
rect 80900 496984 81162 497040
rect 81218 496984 81223 497040
rect 80900 496982 81223 496984
rect 80900 496980 80906 496982
rect 81157 496979 81223 496982
rect 83406 496980 83412 497044
rect 83476 497042 83482 497044
rect 84009 497042 84075 497045
rect 83476 497040 84075 497042
rect 83476 496984 84014 497040
rect 84070 496984 84075 497040
rect 83476 496982 84075 496984
rect 83476 496980 83482 496982
rect 84009 496979 84075 496982
rect 87086 496980 87092 497044
rect 87156 497042 87162 497044
rect 88149 497042 88215 497045
rect 87156 497040 88215 497042
rect 87156 496984 88154 497040
rect 88210 496984 88215 497040
rect 87156 496982 88215 496984
rect 87156 496980 87162 496982
rect 88149 496979 88215 496982
rect 92790 496980 92796 497044
rect 92860 497042 92866 497044
rect 93669 497042 93735 497045
rect 92860 497040 93735 497042
rect 92860 496984 93674 497040
rect 93730 496984 93735 497040
rect 92860 496982 93735 496984
rect 92860 496980 92866 496982
rect 93669 496979 93735 496982
rect 95182 496980 95188 497044
rect 95252 497042 95258 497044
rect 96429 497042 96495 497045
rect 95252 497040 96495 497042
rect 95252 496984 96434 497040
rect 96490 496984 96495 497040
rect 95252 496982 96495 496984
rect 95252 496980 95258 496982
rect 96429 496979 96495 496982
rect 98310 496980 98316 497044
rect 98380 497042 98386 497044
rect 99281 497042 99347 497045
rect 98380 497040 99347 497042
rect 98380 496984 99286 497040
rect 99342 496984 99347 497040
rect 98380 496982 99347 496984
rect 98380 496980 98386 496982
rect 99281 496979 99347 496982
rect 100886 496980 100892 497044
rect 100956 497042 100962 497044
rect 101949 497042 102015 497045
rect 106089 497044 106155 497045
rect 106038 497042 106044 497044
rect 100956 497040 102015 497042
rect 100956 496984 101954 497040
rect 102010 496984 102015 497040
rect 100956 496982 102015 496984
rect 105998 496982 106044 497042
rect 106108 497040 106155 497044
rect 106150 496984 106155 497040
rect 100956 496980 100962 496982
rect 101949 496979 102015 496982
rect 106038 496980 106044 496982
rect 106108 496980 106155 496984
rect 108062 496980 108068 497044
rect 108132 497042 108138 497044
rect 108849 497042 108915 497045
rect 108132 497040 108915 497042
rect 108132 496984 108854 497040
rect 108910 496984 108915 497040
rect 108132 496982 108915 496984
rect 108132 496980 108138 496982
rect 106089 496979 106155 496980
rect 108849 496979 108915 496982
rect 426433 497042 426499 497045
rect 426566 497042 426572 497044
rect 426433 497040 426572 497042
rect 426433 496984 426438 497040
rect 426494 496984 426572 497040
rect 426433 496982 426572 496984
rect 426433 496979 426499 496982
rect 426566 496980 426572 496982
rect 426636 496980 426642 497044
rect 427905 497042 427971 497045
rect 428222 497042 428228 497044
rect 427905 497040 428228 497042
rect 427905 496984 427910 497040
rect 427966 496984 428228 497040
rect 427905 496982 428228 496984
rect 427905 496979 427971 496982
rect 428222 496980 428228 496982
rect 428292 496980 428298 497044
rect 430573 497042 430639 497045
rect 431166 497042 431172 497044
rect 430573 497040 431172 497042
rect 430573 496984 430578 497040
rect 430634 496984 431172 497040
rect 430573 496982 431172 496984
rect 430573 496979 430639 496982
rect 431166 496980 431172 496982
rect 431236 496980 431242 497044
rect 433425 497042 433491 497045
rect 433558 497042 433564 497044
rect 433425 497040 433564 497042
rect 433425 496984 433430 497040
rect 433486 496984 433564 497040
rect 433425 496982 433564 496984
rect 433425 496979 433491 496982
rect 433558 496980 433564 496982
rect 433628 496980 433634 497044
rect 434713 497042 434779 497045
rect 435950 497042 435956 497044
rect 434713 497040 435956 497042
rect 434713 496984 434718 497040
rect 434774 496984 435956 497040
rect 434713 496982 435956 496984
rect 434713 496979 434779 496982
rect 435950 496980 435956 496982
rect 436020 496980 436026 497044
rect 437473 497042 437539 497045
rect 438526 497042 438532 497044
rect 437473 497040 438532 497042
rect 437473 496984 437478 497040
rect 437534 496984 438532 497040
rect 437473 496982 438532 496984
rect 437473 496979 437539 496982
rect 438526 496980 438532 496982
rect 438596 496980 438602 497044
rect 441613 497042 441679 497045
rect 442758 497042 442764 497044
rect 441613 497040 442764 497042
rect 441613 496984 441618 497040
rect 441674 496984 442764 497040
rect 441613 496982 442764 496984
rect 441613 496979 441679 496982
rect 442758 496980 442764 496982
rect 442828 496980 442834 497044
rect 443085 497042 443151 497045
rect 443862 497042 443868 497044
rect 443085 497040 443868 497042
rect 443085 496984 443090 497040
rect 443146 496984 443868 497040
rect 443085 496982 443868 496984
rect 443085 496979 443151 496982
rect 443862 496980 443868 496982
rect 443932 496980 443938 497044
rect 445845 497042 445911 497045
rect 446254 497042 446260 497044
rect 445845 497040 446260 497042
rect 445845 496984 445850 497040
rect 445906 496984 446260 497040
rect 445845 496982 446260 496984
rect 445845 496979 445911 496982
rect 446254 496980 446260 496982
rect 446324 496980 446330 497044
rect 447133 497042 447199 497045
rect 448278 497042 448284 497044
rect 447133 497040 448284 497042
rect 447133 496984 447138 497040
rect 447194 496984 448284 497040
rect 447133 496982 448284 496984
rect 447133 496979 447199 496982
rect 448278 496980 448284 496982
rect 448348 496980 448354 497044
rect 448605 497042 448671 497045
rect 449750 497042 449756 497044
rect 448605 497040 449756 497042
rect 448605 496984 448610 497040
rect 448666 496984 449756 497040
rect 448605 496982 449756 496984
rect 448605 496979 448671 496982
rect 449750 496980 449756 496982
rect 449820 496980 449826 497044
rect 449985 497042 450051 497045
rect 451038 497042 451044 497044
rect 449985 497040 451044 497042
rect 449985 496984 449990 497040
rect 450046 496984 451044 497040
rect 449985 496982 451044 496984
rect 449985 496979 450051 496982
rect 451038 496980 451044 496982
rect 451108 496980 451114 497044
rect 452653 497042 452719 497045
rect 453614 497042 453620 497044
rect 452653 497040 453620 497042
rect 452653 496984 452658 497040
rect 452714 496984 453620 497040
rect 452653 496982 453620 496984
rect 452653 496979 452719 496982
rect 453614 496980 453620 496982
rect 453684 496980 453690 497044
rect 458265 497042 458331 497045
rect 458950 497042 458956 497044
rect 458265 497040 458956 497042
rect 458265 496984 458270 497040
rect 458326 496984 458956 497040
rect 458265 496982 458956 496984
rect 458265 496979 458331 496982
rect 458950 496980 458956 496982
rect 459020 496980 459026 497044
rect 498193 497042 498259 497045
rect 498510 497042 498516 497044
rect 498193 497040 498516 497042
rect 498193 496984 498198 497040
rect 498254 496984 498516 497040
rect 498193 496982 498516 496984
rect 498193 496979 498259 496982
rect 498510 496980 498516 496982
rect 498580 496980 498586 497044
rect 66161 496908 66227 496909
rect 66110 496906 66116 496908
rect 66070 496846 66116 496906
rect 66180 496904 66227 496908
rect 66222 496848 66227 496904
rect 66110 496844 66116 496846
rect 66180 496844 66227 496848
rect 68318 496844 68324 496908
rect 68388 496906 68394 496908
rect 68921 496906 68987 496909
rect 68388 496904 68987 496906
rect 68388 496848 68926 496904
rect 68982 496848 68987 496904
rect 68388 496846 68987 496848
rect 68388 496844 68394 496846
rect 66161 496843 66227 496844
rect 68921 496843 68987 496846
rect 69606 496844 69612 496908
rect 69676 496906 69682 496908
rect 70301 496906 70367 496909
rect 69676 496904 70367 496906
rect 69676 496848 70306 496904
rect 70362 496848 70367 496904
rect 69676 496846 70367 496848
rect 69676 496844 69682 496846
rect 70301 496843 70367 496846
rect 70526 496844 70532 496908
rect 70596 496906 70602 496908
rect 71681 496906 71747 496909
rect 70596 496904 71747 496906
rect 70596 496848 71686 496904
rect 71742 496848 71747 496904
rect 70596 496846 71747 496848
rect 70596 496844 70602 496846
rect 71681 496843 71747 496846
rect 75494 496844 75500 496908
rect 75564 496906 75570 496908
rect 75821 496906 75887 496909
rect 75564 496904 75887 496906
rect 75564 496848 75826 496904
rect 75882 496848 75887 496904
rect 75564 496846 75887 496848
rect 75564 496844 75570 496846
rect 75821 496843 75887 496846
rect 76598 496844 76604 496908
rect 76668 496906 76674 496908
rect 77201 496906 77267 496909
rect 78305 496908 78371 496909
rect 78254 496906 78260 496908
rect 76668 496904 77267 496906
rect 76668 496848 77206 496904
rect 77262 496848 77267 496904
rect 76668 496846 77267 496848
rect 78214 496846 78260 496906
rect 78324 496904 78371 496908
rect 78366 496848 78371 496904
rect 76668 496844 76674 496846
rect 77201 496843 77267 496846
rect 78254 496844 78260 496846
rect 78324 496844 78371 496848
rect 81014 496844 81020 496908
rect 81084 496906 81090 496908
rect 81249 496906 81315 496909
rect 81084 496904 81315 496906
rect 81084 496848 81254 496904
rect 81310 496848 81315 496904
rect 81084 496846 81315 496848
rect 81084 496844 81090 496846
rect 78305 496843 78371 496844
rect 81249 496843 81315 496846
rect 82486 496844 82492 496908
rect 82556 496906 82562 496908
rect 82721 496906 82787 496909
rect 82556 496904 82787 496906
rect 82556 496848 82726 496904
rect 82782 496848 82787 496904
rect 82556 496846 82787 496848
rect 82556 496844 82562 496846
rect 82721 496843 82787 496846
rect 83590 496844 83596 496908
rect 83660 496906 83666 496908
rect 84101 496906 84167 496909
rect 83660 496904 84167 496906
rect 83660 496848 84106 496904
rect 84162 496848 84167 496904
rect 83660 496846 84167 496848
rect 83660 496844 83666 496846
rect 84101 496843 84167 496846
rect 84510 496844 84516 496908
rect 84580 496906 84586 496908
rect 85481 496906 85547 496909
rect 88241 496908 88307 496909
rect 88190 496906 88196 496908
rect 84580 496904 85547 496906
rect 84580 496848 85486 496904
rect 85542 496848 85547 496904
rect 84580 496846 85547 496848
rect 88150 496846 88196 496906
rect 88260 496904 88307 496908
rect 88302 496848 88307 496904
rect 84580 496844 84586 496846
rect 85481 496843 85547 496846
rect 88190 496844 88196 496846
rect 88260 496844 88307 496848
rect 88558 496844 88564 496908
rect 88628 496906 88634 496908
rect 89161 496906 89227 496909
rect 88628 496904 89227 496906
rect 88628 496848 89166 496904
rect 89222 496848 89227 496904
rect 88628 496846 89227 496848
rect 88628 496844 88634 496846
rect 88241 496843 88307 496844
rect 89161 496843 89227 496846
rect 90766 496844 90772 496908
rect 90836 496906 90842 496908
rect 91001 496906 91067 496909
rect 91185 496908 91251 496909
rect 90836 496904 91067 496906
rect 90836 496848 91006 496904
rect 91062 496848 91067 496904
rect 90836 496846 91067 496848
rect 90836 496844 90842 496846
rect 91001 496843 91067 496846
rect 91134 496844 91140 496908
rect 91204 496906 91251 496908
rect 91204 496904 91296 496906
rect 91246 496848 91296 496904
rect 91204 496846 91296 496848
rect 91204 496844 91251 496846
rect 93526 496844 93532 496908
rect 93596 496906 93602 496908
rect 93761 496906 93827 496909
rect 93596 496904 93827 496906
rect 93596 496848 93766 496904
rect 93822 496848 93827 496904
rect 93596 496846 93827 496848
rect 93596 496844 93602 496846
rect 91185 496843 91251 496844
rect 93761 496843 93827 496846
rect 93894 496844 93900 496908
rect 93964 496906 93970 496908
rect 95141 496906 95207 496909
rect 93964 496904 95207 496906
rect 93964 496848 95146 496904
rect 95202 496848 95207 496904
rect 93964 496846 95207 496848
rect 93964 496844 93970 496846
rect 95141 496843 95207 496846
rect 97574 496844 97580 496908
rect 97644 496906 97650 496908
rect 97901 496906 97967 496909
rect 97644 496904 97967 496906
rect 97644 496848 97906 496904
rect 97962 496848 97967 496904
rect 97644 496846 97967 496848
rect 97644 496844 97650 496846
rect 97901 496843 97967 496846
rect 98678 496844 98684 496908
rect 98748 496906 98754 496908
rect 99189 496906 99255 496909
rect 98748 496904 99255 496906
rect 98748 496848 99194 496904
rect 99250 496848 99255 496904
rect 98748 496846 99255 496848
rect 98748 496844 98754 496846
rect 99189 496843 99255 496846
rect 99966 496844 99972 496908
rect 100036 496906 100042 496908
rect 100661 496906 100727 496909
rect 100036 496904 100727 496906
rect 100036 496848 100666 496904
rect 100722 496848 100727 496904
rect 100036 496846 100727 496848
rect 100036 496844 100042 496846
rect 100661 496843 100727 496846
rect 101254 496844 101260 496908
rect 101324 496906 101330 496908
rect 102041 496906 102107 496909
rect 101324 496904 102107 496906
rect 101324 496848 102046 496904
rect 102102 496848 102107 496904
rect 101324 496846 102107 496848
rect 101324 496844 101330 496846
rect 102041 496843 102107 496846
rect 102174 496844 102180 496908
rect 102244 496906 102250 496908
rect 103329 496906 103395 496909
rect 102244 496904 103395 496906
rect 102244 496848 103334 496904
rect 103390 496848 103395 496904
rect 102244 496846 103395 496848
rect 102244 496844 102250 496846
rect 103329 496843 103395 496846
rect 104382 496844 104388 496908
rect 104452 496906 104458 496908
rect 104709 496906 104775 496909
rect 104452 496904 104775 496906
rect 104452 496848 104714 496904
rect 104770 496848 104775 496904
rect 104452 496846 104775 496848
rect 104452 496844 104458 496846
rect 104709 496843 104775 496846
rect 105854 496844 105860 496908
rect 105924 496906 105930 496908
rect 106181 496906 106247 496909
rect 105924 496904 106247 496906
rect 105924 496848 106186 496904
rect 106242 496848 106247 496904
rect 105924 496846 106247 496848
rect 105924 496844 105930 496846
rect 106181 496843 106247 496846
rect 106958 496844 106964 496908
rect 107028 496906 107034 496908
rect 107561 496906 107627 496909
rect 107028 496904 107627 496906
rect 107028 496848 107566 496904
rect 107622 496848 107627 496904
rect 107028 496846 107627 496848
rect 107028 496844 107034 496846
rect 107561 496843 107627 496846
rect 108430 496844 108436 496908
rect 108500 496906 108506 496908
rect 108941 496906 109007 496909
rect 108500 496904 109007 496906
rect 108500 496848 108946 496904
rect 109002 496848 109007 496904
rect 108500 496846 109007 496848
rect 108500 496844 108506 496846
rect 108941 496843 109007 496846
rect 109166 496844 109172 496908
rect 109236 496906 109242 496908
rect 110321 496906 110387 496909
rect 109236 496904 110387 496906
rect 109236 496848 110326 496904
rect 110382 496848 110387 496904
rect 109236 496846 110387 496848
rect 109236 496844 109242 496846
rect 110321 496843 110387 496846
rect 111006 496844 111012 496908
rect 111076 496906 111082 496908
rect 111701 496906 111767 496909
rect 111076 496904 111767 496906
rect 111076 496848 111706 496904
rect 111762 496848 111767 496904
rect 111076 496846 111767 496848
rect 111076 496844 111082 496846
rect 111701 496843 111767 496846
rect 123518 496844 123524 496908
rect 123588 496906 123594 496908
rect 124121 496906 124187 496909
rect 123588 496904 124187 496906
rect 123588 496848 124126 496904
rect 124182 496848 124187 496904
rect 123588 496846 124187 496848
rect 123588 496844 123594 496846
rect 124121 496843 124187 496846
rect 130878 496844 130884 496908
rect 130948 496906 130954 496908
rect 131021 496906 131087 496909
rect 130948 496904 131087 496906
rect 130948 496848 131026 496904
rect 131082 496848 131087 496904
rect 130948 496846 131087 496848
rect 130948 496844 130954 496846
rect 131021 496843 131087 496846
rect 133454 496844 133460 496908
rect 133524 496906 133530 496908
rect 133781 496906 133847 496909
rect 133524 496904 133847 496906
rect 133524 496848 133786 496904
rect 133842 496848 133847 496904
rect 133524 496846 133847 496848
rect 133524 496844 133530 496846
rect 133781 496843 133847 496846
rect 136030 496844 136036 496908
rect 136100 496906 136106 496908
rect 136541 496906 136607 496909
rect 136100 496904 136607 496906
rect 136100 496848 136546 496904
rect 136602 496848 136607 496904
rect 136100 496846 136607 496848
rect 136100 496844 136106 496846
rect 136541 496843 136607 496846
rect 138606 496844 138612 496908
rect 138676 496906 138682 496908
rect 139301 496906 139367 496909
rect 138676 496904 139367 496906
rect 138676 496848 139306 496904
rect 139362 496848 139367 496904
rect 138676 496846 139367 496848
rect 138676 496844 138682 496846
rect 139301 496843 139367 496846
rect 140998 496844 141004 496908
rect 141068 496906 141074 496908
rect 142061 496906 142127 496909
rect 143441 496908 143507 496909
rect 143390 496906 143396 496908
rect 141068 496904 142127 496906
rect 141068 496848 142066 496904
rect 142122 496848 142127 496904
rect 141068 496846 142127 496848
rect 143350 496846 143396 496906
rect 143460 496904 143507 496908
rect 143502 496848 143507 496904
rect 141068 496844 141074 496846
rect 142061 496843 142127 496846
rect 143390 496844 143396 496846
rect 143460 496844 143507 496848
rect 148542 496844 148548 496908
rect 148612 496906 148618 496908
rect 148961 496906 149027 496909
rect 148612 496904 149027 496906
rect 148612 496848 148966 496904
rect 149022 496848 149027 496904
rect 148612 496846 149027 496848
rect 148612 496844 148618 496846
rect 143441 496843 143507 496844
rect 148961 496843 149027 496846
rect 155902 496844 155908 496908
rect 155972 496906 155978 496908
rect 157241 496906 157307 496909
rect 155972 496904 157307 496906
rect 155972 496848 157246 496904
rect 157302 496848 157307 496904
rect 155972 496846 157307 496848
rect 155972 496844 155978 496846
rect 157241 496843 157307 496846
rect 415393 496906 415459 496909
rect 415526 496906 415532 496908
rect 415393 496904 415532 496906
rect 415393 496848 415398 496904
rect 415454 496848 415532 496904
rect 415393 496846 415532 496848
rect 415393 496843 415459 496846
rect 415526 496844 415532 496846
rect 415596 496844 415602 496908
rect 416773 496906 416839 496909
rect 417182 496906 417188 496908
rect 416773 496904 417188 496906
rect 416773 496848 416778 496904
rect 416834 496848 417188 496904
rect 416773 496846 417188 496848
rect 416773 496843 416839 496846
rect 417182 496844 417188 496846
rect 417252 496844 417258 496908
rect 418153 496906 418219 496909
rect 418286 496906 418292 496908
rect 418153 496904 418292 496906
rect 418153 496848 418158 496904
rect 418214 496848 418292 496904
rect 418153 496846 418292 496848
rect 418153 496843 418219 496846
rect 418286 496844 418292 496846
rect 418356 496844 418362 496908
rect 419533 496906 419599 496909
rect 420494 496906 420500 496908
rect 419533 496904 420500 496906
rect 419533 496848 419538 496904
rect 419594 496848 420500 496904
rect 419533 496846 420500 496848
rect 419533 496843 419599 496846
rect 420494 496844 420500 496846
rect 420564 496844 420570 496908
rect 420913 496906 420979 496909
rect 421782 496906 421788 496908
rect 420913 496904 421788 496906
rect 420913 496848 420918 496904
rect 420974 496848 421788 496904
rect 420913 496846 421788 496848
rect 420913 496843 420979 496846
rect 421782 496844 421788 496846
rect 421852 496844 421858 496908
rect 422293 496906 422359 496909
rect 423070 496906 423076 496908
rect 422293 496904 423076 496906
rect 422293 496848 422298 496904
rect 422354 496848 423076 496904
rect 422293 496846 423076 496848
rect 422293 496843 422359 496846
rect 423070 496844 423076 496846
rect 423140 496844 423146 496908
rect 423673 496906 423739 496909
rect 424174 496906 424180 496908
rect 423673 496904 424180 496906
rect 423673 496848 423678 496904
rect 423734 496848 424180 496904
rect 423673 496846 424180 496848
rect 423673 496843 423739 496846
rect 424174 496844 424180 496846
rect 424244 496844 424250 496908
rect 425053 496906 425119 496909
rect 425462 496906 425468 496908
rect 425053 496904 425468 496906
rect 425053 496848 425058 496904
rect 425114 496848 425468 496904
rect 425053 496846 425468 496848
rect 425053 496843 425119 496846
rect 425462 496844 425468 496846
rect 425532 496844 425538 496908
rect 426525 496906 426591 496909
rect 427670 496906 427676 496908
rect 426525 496904 427676 496906
rect 426525 496848 426530 496904
rect 426586 496848 427676 496904
rect 426525 496846 427676 496848
rect 426525 496843 426591 496846
rect 427670 496844 427676 496846
rect 427740 496844 427746 496908
rect 427813 496906 427879 496909
rect 428590 496906 428596 496908
rect 427813 496904 428596 496906
rect 427813 496848 427818 496904
rect 427874 496848 428596 496904
rect 427813 496846 428596 496848
rect 427813 496843 427879 496846
rect 428590 496844 428596 496846
rect 428660 496844 428666 496908
rect 429193 496906 429259 496909
rect 430062 496906 430068 496908
rect 429193 496904 430068 496906
rect 429193 496848 429198 496904
rect 429254 496848 430068 496904
rect 429193 496846 430068 496848
rect 429193 496843 429259 496846
rect 430062 496844 430068 496846
rect 430132 496844 430138 496908
rect 430665 496906 430731 496909
rect 433333 496908 433399 496909
rect 430798 496906 430804 496908
rect 430665 496904 430804 496906
rect 430665 496848 430670 496904
rect 430726 496848 430804 496904
rect 430665 496846 430804 496848
rect 430665 496843 430731 496846
rect 430798 496844 430804 496846
rect 430868 496844 430874 496908
rect 433333 496906 433380 496908
rect 433288 496904 433380 496906
rect 433288 496848 433338 496904
rect 433288 496846 433380 496848
rect 433333 496844 433380 496846
rect 433444 496844 433450 496908
rect 434805 496906 434871 496909
rect 435766 496906 435772 496908
rect 434805 496904 435772 496906
rect 434805 496848 434810 496904
rect 434866 496848 435772 496904
rect 434805 496846 435772 496848
rect 433333 496843 433399 496844
rect 434805 496843 434871 496846
rect 435766 496844 435772 496846
rect 435836 496844 435842 496908
rect 436093 496906 436159 496909
rect 436870 496906 436876 496908
rect 436093 496904 436876 496906
rect 436093 496848 436098 496904
rect 436154 496848 436876 496904
rect 436093 496846 436876 496848
rect 436093 496843 436159 496846
rect 436870 496844 436876 496846
rect 436940 496844 436946 496908
rect 437565 496906 437631 496909
rect 438342 496906 438348 496908
rect 437565 496904 438348 496906
rect 437565 496848 437570 496904
rect 437626 496848 438348 496904
rect 437565 496846 438348 496848
rect 437565 496843 437631 496846
rect 438342 496844 438348 496846
rect 438412 496844 438418 496908
rect 438853 496906 438919 496909
rect 439446 496906 439452 496908
rect 438853 496904 439452 496906
rect 438853 496848 438858 496904
rect 438914 496848 439452 496904
rect 438853 496846 439452 496848
rect 438853 496843 438919 496846
rect 439446 496844 439452 496846
rect 439516 496844 439522 496908
rect 440325 496906 440391 496909
rect 440550 496906 440556 496908
rect 440325 496904 440556 496906
rect 440325 496848 440330 496904
rect 440386 496848 440556 496904
rect 440325 496846 440556 496848
rect 440325 496843 440391 496846
rect 440550 496844 440556 496846
rect 440620 496844 440626 496908
rect 441705 496906 441771 496909
rect 442022 496906 442028 496908
rect 441705 496904 442028 496906
rect 441705 496848 441710 496904
rect 441766 496848 442028 496904
rect 441705 496846 442028 496848
rect 441705 496843 441771 496846
rect 442022 496844 442028 496846
rect 442092 496844 442098 496908
rect 442993 496906 443059 496909
rect 443494 496906 443500 496908
rect 442993 496904 443500 496906
rect 442993 496848 442998 496904
rect 443054 496848 443500 496904
rect 442993 496846 443500 496848
rect 442993 496843 443059 496846
rect 443494 496844 443500 496846
rect 443564 496844 443570 496908
rect 444373 496906 444439 496909
rect 445937 496908 446003 496909
rect 444782 496906 444788 496908
rect 444373 496904 444788 496906
rect 444373 496848 444378 496904
rect 444434 496848 444788 496904
rect 444373 496846 444788 496848
rect 444373 496843 444439 496846
rect 444782 496844 444788 496846
rect 444852 496844 444858 496908
rect 445886 496844 445892 496908
rect 445956 496906 446003 496908
rect 447225 496906 447291 496909
rect 447542 496906 447548 496908
rect 445956 496904 446048 496906
rect 445998 496848 446048 496904
rect 445956 496846 446048 496848
rect 447225 496904 447548 496906
rect 447225 496848 447230 496904
rect 447286 496848 447548 496904
rect 447225 496846 447548 496848
rect 445956 496844 446003 496846
rect 445937 496843 446003 496844
rect 447225 496843 447291 496846
rect 447542 496844 447548 496846
rect 447612 496844 447618 496908
rect 448513 496906 448579 496909
rect 448646 496906 448652 496908
rect 448513 496904 448652 496906
rect 448513 496848 448518 496904
rect 448574 496848 448652 496904
rect 448513 496846 448652 496848
rect 448513 496843 448579 496846
rect 448646 496844 448652 496846
rect 448716 496844 448722 496908
rect 449893 496906 449959 496909
rect 450854 496906 450860 496908
rect 449893 496904 450860 496906
rect 449893 496848 449898 496904
rect 449954 496848 450860 496904
rect 449893 496846 450860 496848
rect 449893 496843 449959 496846
rect 450854 496844 450860 496846
rect 450924 496844 450930 496908
rect 451273 496906 451339 496909
rect 452510 496906 452516 496908
rect 451273 496904 452516 496906
rect 451273 496848 451278 496904
rect 451334 496848 452516 496904
rect 451273 496846 452516 496848
rect 451273 496843 451339 496846
rect 452510 496844 452516 496846
rect 452580 496844 452586 496908
rect 452745 496906 452811 496909
rect 453246 496906 453252 496908
rect 452745 496904 453252 496906
rect 452745 496848 452750 496904
rect 452806 496848 453252 496904
rect 452745 496846 453252 496848
rect 452745 496843 452811 496846
rect 453246 496844 453252 496846
rect 453316 496844 453322 496908
rect 454033 496906 454099 496909
rect 456885 496908 456951 496909
rect 454350 496906 454356 496908
rect 454033 496904 454356 496906
rect 454033 496848 454038 496904
rect 454094 496848 454356 496904
rect 454033 496846 454356 496848
rect 454033 496843 454099 496846
rect 454350 496844 454356 496846
rect 454420 496844 454426 496908
rect 456885 496906 456932 496908
rect 456840 496904 456932 496906
rect 456840 496848 456890 496904
rect 456840 496846 456932 496848
rect 456885 496844 456932 496846
rect 456996 496844 457002 496908
rect 458173 496906 458239 496909
rect 460933 496908 460999 496909
rect 458398 496906 458404 496908
rect 458173 496904 458404 496906
rect 458173 496848 458178 496904
rect 458234 496848 458404 496904
rect 458173 496846 458404 496848
rect 456885 496843 456951 496844
rect 458173 496843 458239 496846
rect 458398 496844 458404 496846
rect 458468 496844 458474 496908
rect 460933 496904 460980 496908
rect 461044 496906 461050 496908
rect 465073 496906 465139 496909
rect 465942 496906 465948 496908
rect 460933 496848 460938 496904
rect 460933 496844 460980 496848
rect 461044 496846 461090 496906
rect 465073 496904 465948 496906
rect 465073 496848 465078 496904
rect 465134 496848 465948 496904
rect 465073 496846 465948 496848
rect 461044 496844 461050 496846
rect 460933 496843 460999 496844
rect 465073 496843 465139 496846
rect 465942 496844 465948 496846
rect 466012 496844 466018 496908
rect 467833 496906 467899 496909
rect 468150 496906 468156 496908
rect 467833 496904 468156 496906
rect 467833 496848 467838 496904
rect 467894 496848 468156 496904
rect 467833 496846 468156 496848
rect 467833 496843 467899 496846
rect 468150 496844 468156 496846
rect 468220 496844 468226 496908
rect 470593 496906 470659 496909
rect 473353 496908 473419 496909
rect 470910 496906 470916 496908
rect 470593 496904 470916 496906
rect 470593 496848 470598 496904
rect 470654 496848 470916 496904
rect 470593 496846 470916 496848
rect 470593 496843 470659 496846
rect 470910 496844 470916 496846
rect 470980 496844 470986 496908
rect 473302 496844 473308 496908
rect 473372 496906 473419 496908
rect 474733 496906 474799 496909
rect 475878 496906 475884 496908
rect 473372 496904 473464 496906
rect 473414 496848 473464 496904
rect 473372 496846 473464 496848
rect 474733 496904 475884 496906
rect 474733 496848 474738 496904
rect 474794 496848 475884 496904
rect 474733 496846 475884 496848
rect 473372 496844 473419 496846
rect 473353 496843 473419 496844
rect 474733 496843 474799 496846
rect 475878 496844 475884 496846
rect 475948 496844 475954 496908
rect 477493 496906 477559 496909
rect 478454 496906 478460 496908
rect 477493 496904 478460 496906
rect 477493 496848 477498 496904
rect 477554 496848 478460 496904
rect 477493 496846 478460 496848
rect 477493 496843 477559 496846
rect 478454 496844 478460 496846
rect 478524 496844 478530 496908
rect 480253 496906 480319 496909
rect 480662 496906 480668 496908
rect 480253 496904 480668 496906
rect 480253 496848 480258 496904
rect 480314 496848 480668 496904
rect 480253 496846 480668 496848
rect 480253 496843 480319 496846
rect 480662 496844 480668 496846
rect 480732 496844 480738 496908
rect 483013 496906 483079 496909
rect 483422 496906 483428 496908
rect 483013 496904 483428 496906
rect 483013 496848 483018 496904
rect 483074 496848 483428 496904
rect 483013 496846 483428 496848
rect 483013 496843 483079 496846
rect 483422 496844 483428 496846
rect 483492 496844 483498 496908
rect 485773 496906 485839 496909
rect 488533 496908 488599 496909
rect 485998 496906 486004 496908
rect 485773 496904 486004 496906
rect 485773 496848 485778 496904
rect 485834 496848 486004 496904
rect 485773 496846 486004 496848
rect 485773 496843 485839 496846
rect 485998 496844 486004 496846
rect 486068 496844 486074 496908
rect 488533 496906 488580 496908
rect 488488 496904 488580 496906
rect 488488 496848 488538 496904
rect 488488 496846 488580 496848
rect 488533 496844 488580 496846
rect 488644 496844 488650 496908
rect 489913 496906 489979 496909
rect 490966 496906 490972 496908
rect 489913 496904 490972 496906
rect 489913 496848 489918 496904
rect 489974 496848 490972 496904
rect 489913 496846 490972 496848
rect 488533 496843 488599 496844
rect 489913 496843 489979 496846
rect 490966 496844 490972 496846
rect 491036 496844 491042 496908
rect 492673 496906 492739 496909
rect 493358 496906 493364 496908
rect 492673 496904 493364 496906
rect 492673 496848 492678 496904
rect 492734 496848 493364 496904
rect 492673 496846 493364 496848
rect 492673 496843 492739 496846
rect 493358 496844 493364 496846
rect 493428 496844 493434 496908
rect 495433 496906 495499 496909
rect 500953 496908 501019 496909
rect 495934 496906 495940 496908
rect 495433 496904 495940 496906
rect 495433 496848 495438 496904
rect 495494 496848 495940 496904
rect 495433 496846 495940 496848
rect 495433 496843 495499 496846
rect 495934 496844 495940 496846
rect 496004 496844 496010 496908
rect 500902 496906 500908 496908
rect 500862 496846 500908 496906
rect 500972 496904 501019 496908
rect 501014 496848 501019 496904
rect 500902 496844 500908 496846
rect 500972 496844 501019 496848
rect 500953 496843 501019 496844
rect 502333 496906 502399 496909
rect 503294 496906 503300 496908
rect 502333 496904 503300 496906
rect 502333 496848 502338 496904
rect 502394 496848 503300 496904
rect 502333 496846 503300 496848
rect 502333 496843 502399 496846
rect 503294 496844 503300 496846
rect 503364 496844 503370 496908
rect 505093 496906 505159 496909
rect 505502 496906 505508 496908
rect 505093 496904 505508 496906
rect 505093 496848 505098 496904
rect 505154 496848 505508 496904
rect 505093 496846 505508 496848
rect 505093 496843 505159 496846
rect 505502 496844 505508 496846
rect 505572 496844 505578 496908
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect -960 423452 480 423692
rect 370865 422378 370931 422381
rect 412766 422378 412772 422380
rect 370865 422376 412772 422378
rect 370865 422320 370870 422376
rect 370926 422320 412772 422376
rect 370865 422318 412772 422320
rect 370865 422315 370931 422318
rect 412766 422316 412772 422318
rect 412836 422316 412842 422380
rect 169150 420956 169156 421020
rect 169220 421018 169226 421020
rect 380893 421018 380959 421021
rect 169220 421016 380959 421018
rect 169220 420960 380898 421016
rect 380954 420960 380959 421016
rect 169220 420958 380959 420960
rect 169220 420956 169226 420958
rect 380893 420955 380959 420958
rect 400673 421018 400739 421021
rect 414606 421018 414612 421020
rect 400673 421016 414612 421018
rect 400673 420960 400678 421016
rect 400734 420960 414612 421016
rect 400673 420958 414612 420960
rect 400673 420955 400739 420958
rect 414606 420956 414612 420958
rect 414676 420956 414682 421020
rect 351085 420202 351151 420205
rect 408534 420202 408540 420204
rect 351085 420200 408540 420202
rect 351085 420144 351090 420200
rect 351146 420144 408540 420200
rect 351085 420142 408540 420144
rect 351085 420139 351151 420142
rect 408534 420140 408540 420142
rect 408604 420140 408610 420204
rect 190729 420066 190795 420069
rect 190686 420064 190795 420066
rect 190686 420008 190734 420064
rect 190790 420008 190795 420064
rect 190686 420003 190795 420008
rect 190686 419492 190746 420003
rect 412081 418978 412147 418981
rect 409860 418976 412147 418978
rect 409860 418920 412086 418976
rect 412142 418920 412147 418976
rect 409860 418918 412147 418920
rect 412081 418915 412147 418918
rect 186313 418434 186379 418437
rect 186313 418432 190164 418434
rect 186313 418376 186318 418432
rect 186374 418376 190164 418432
rect 186313 418374 190164 418376
rect 186313 418371 186379 418374
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect 190361 417890 190427 417893
rect 190318 417888 190427 417890
rect 190318 417832 190366 417888
rect 190422 417832 190427 417888
rect 190318 417827 190427 417832
rect 190318 417316 190378 417827
rect 412081 416938 412147 416941
rect 409860 416936 412147 416938
rect 409860 416880 412086 416936
rect 412142 416880 412147 416936
rect 409860 416878 412147 416880
rect 412081 416875 412147 416878
rect 187601 416394 187667 416397
rect 187601 416392 190164 416394
rect 187601 416336 187606 416392
rect 187662 416336 190164 416392
rect 187601 416334 190164 416336
rect 187601 416331 187667 416334
rect 186313 415306 186379 415309
rect 186313 415304 190164 415306
rect 186313 415248 186318 415304
rect 186374 415248 190164 415304
rect 186313 415246 190164 415248
rect 186313 415243 186379 415246
rect 410701 414898 410767 414901
rect 409860 414896 410767 414898
rect 409860 414840 410706 414896
rect 410762 414840 410767 414896
rect 409860 414838 410767 414840
rect 410701 414835 410767 414838
rect 187509 414218 187575 414221
rect 187509 414216 190164 414218
rect 187509 414160 187514 414216
rect 187570 414160 190164 414216
rect 187509 414158 190164 414160
rect 187509 414155 187575 414158
rect 186865 413130 186931 413133
rect 409321 413130 409387 413133
rect 186865 413128 190164 413130
rect 186865 413072 186870 413128
rect 186926 413072 190164 413128
rect 186865 413070 190164 413072
rect 409278 413128 409387 413130
rect 409278 413072 409326 413128
rect 409382 413072 409387 413128
rect 186865 413067 186931 413070
rect 409278 413067 409387 413072
rect 409278 412828 409338 413067
rect 186313 412178 186379 412181
rect 186313 412176 190164 412178
rect 186313 412120 186318 412176
rect 186374 412120 190164 412176
rect 186313 412118 190164 412120
rect 186313 412115 186379 412118
rect 186313 411090 186379 411093
rect 186313 411088 190164 411090
rect 186313 411032 186318 411088
rect 186374 411032 190164 411088
rect 186313 411030 190164 411032
rect 186313 411027 186379 411030
rect -960 410396 480 410636
rect 409278 410277 409338 410788
rect 409278 410272 409387 410277
rect 409278 410216 409326 410272
rect 409382 410216 409387 410272
rect 409278 410214 409387 410216
rect 409321 410211 409387 410214
rect 186405 410002 186471 410005
rect 186405 410000 190164 410002
rect 186405 409944 186410 410000
rect 186466 409944 190164 410000
rect 186405 409942 190164 409944
rect 186405 409939 186471 409942
rect 437473 409186 437539 409189
rect 437473 409184 440036 409186
rect 437473 409128 437478 409184
rect 437534 409128 440036 409184
rect 437473 409126 440036 409128
rect 437473 409123 437539 409126
rect 189165 408914 189231 408917
rect 189165 408912 190164 408914
rect 189165 408856 189170 408912
rect 189226 408856 190164 408912
rect 189165 408854 190164 408856
rect 189165 408851 189231 408854
rect 409822 408852 409828 408916
rect 409892 408852 409898 408916
rect 409830 408748 409890 408852
rect 187509 407962 187575 407965
rect 187509 407960 190164 407962
rect 187509 407904 187514 407960
rect 187570 407904 190164 407960
rect 187509 407902 190164 407904
rect 187509 407899 187575 407902
rect 437473 407554 437539 407557
rect 437473 407552 440036 407554
rect 437473 407496 437478 407552
rect 437534 407496 440036 407552
rect 437473 407494 440036 407496
rect 437473 407491 437539 407494
rect 186313 406874 186379 406877
rect 186313 406872 190164 406874
rect 186313 406816 186318 406872
rect 186374 406816 190164 406872
rect 186313 406814 190164 406816
rect 186313 406811 186379 406814
rect 412950 406738 412956 406740
rect 409860 406678 412956 406738
rect 412950 406676 412956 406678
rect 413020 406676 413026 406740
rect 437473 405922 437539 405925
rect 437473 405920 440036 405922
rect 437473 405864 437478 405920
rect 437534 405864 440036 405920
rect 437473 405862 440036 405864
rect 437473 405859 437539 405862
rect 188797 405786 188863 405789
rect 188797 405784 190164 405786
rect 188797 405728 188802 405784
rect 188858 405728 190164 405784
rect 188797 405726 190164 405728
rect 188797 405723 188863 405726
rect 583520 404820 584960 405060
rect 188705 404698 188771 404701
rect 188705 404696 190164 404698
rect 188705 404640 188710 404696
rect 188766 404640 190164 404696
rect 188705 404638 190164 404640
rect 188705 404635 188771 404638
rect 409321 404426 409387 404429
rect 409462 404426 409522 404668
rect 409321 404424 409522 404426
rect 409321 404368 409326 404424
rect 409382 404368 409522 404424
rect 409321 404366 409522 404368
rect 409321 404363 409387 404366
rect 437473 404290 437539 404293
rect 437473 404288 440036 404290
rect 437473 404232 437478 404288
rect 437534 404232 440036 404288
rect 437473 404230 440036 404232
rect 437473 404227 437539 404230
rect 186313 403746 186379 403749
rect 186313 403744 190164 403746
rect 186313 403688 186318 403744
rect 186374 403688 190164 403744
rect 186313 403686 190164 403688
rect 186313 403683 186379 403686
rect 550633 403066 550699 403069
rect 549884 403064 550699 403066
rect 549884 403008 550638 403064
rect 550694 403008 550699 403064
rect 549884 403006 550699 403008
rect 550633 403003 550699 403006
rect 187049 402658 187115 402661
rect 437473 402658 437539 402661
rect 187049 402656 190164 402658
rect 187049 402600 187054 402656
rect 187110 402600 190164 402656
rect 187049 402598 190164 402600
rect 437473 402656 440036 402658
rect 437473 402600 437478 402656
rect 437534 402600 440036 402656
rect 437473 402598 440036 402600
rect 187049 402595 187115 402598
rect 437473 402595 437539 402598
rect 409830 401978 409890 402492
rect 412398 401978 412404 401980
rect 409830 401918 412404 401978
rect 412398 401916 412404 401918
rect 412468 401916 412474 401980
rect 186313 401570 186379 401573
rect 186313 401568 190164 401570
rect 186313 401512 186318 401568
rect 186374 401512 190164 401568
rect 186313 401510 190164 401512
rect 186313 401507 186379 401510
rect 437473 401026 437539 401029
rect 437473 401024 440036 401026
rect 437473 400968 437478 401024
rect 437534 400968 440036 401024
rect 437473 400966 440036 400968
rect 437473 400963 437539 400966
rect 187509 400482 187575 400485
rect 410609 400482 410675 400485
rect 187509 400480 190164 400482
rect 187509 400424 187514 400480
rect 187570 400424 190164 400480
rect 187509 400422 190164 400424
rect 409860 400480 410675 400482
rect 409860 400424 410614 400480
rect 410670 400424 410675 400480
rect 409860 400422 410675 400424
rect 187509 400419 187575 400422
rect 410609 400419 410675 400422
rect 131941 400210 132007 400213
rect 129782 400208 132007 400210
rect 129782 400152 131946 400208
rect 132002 400152 132007 400208
rect 129782 400150 132007 400152
rect 129782 399636 129842 400150
rect 131941 400147 132007 400150
rect 189257 399530 189323 399533
rect 189257 399528 190164 399530
rect 189257 399472 189262 399528
rect 189318 399472 190164 399528
rect 189257 399470 190164 399472
rect 189257 399467 189323 399470
rect 437473 399394 437539 399397
rect 437473 399392 440036 399394
rect 437473 399336 437478 399392
rect 437534 399336 440036 399392
rect 437473 399334 440036 399336
rect 437473 399331 437539 399334
rect 131205 399122 131271 399125
rect 129968 399120 131271 399122
rect 129968 399064 131210 399120
rect 131266 399064 131271 399120
rect 129968 399062 131271 399064
rect 131205 399059 131271 399062
rect 409413 398850 409479 398853
rect 409413 398848 409522 398850
rect 409413 398792 409418 398848
rect 409474 398792 409522 398848
rect 409413 398787 409522 398792
rect 131205 398578 131271 398581
rect 129968 398576 131271 398578
rect 129968 398520 131210 398576
rect 131266 398520 131271 398576
rect 129968 398518 131271 398520
rect 131205 398515 131271 398518
rect 189349 398442 189415 398445
rect 189349 398440 190164 398442
rect 189349 398384 189354 398440
rect 189410 398384 190164 398440
rect 409462 398412 409522 398787
rect 189349 398382 190164 398384
rect 189349 398379 189415 398382
rect 131941 397898 132007 397901
rect 129968 397896 132007 397898
rect 129968 397840 131946 397896
rect 132002 397840 132007 397896
rect 129968 397838 132007 397840
rect 131941 397835 132007 397838
rect 437565 397762 437631 397765
rect 437565 397760 440036 397762
rect 437565 397704 437570 397760
rect 437626 397704 440036 397760
rect 437565 397702 440036 397704
rect 437565 397699 437631 397702
rect -960 397340 480 397580
rect 131481 397354 131547 397357
rect 129968 397352 131547 397354
rect 129968 397296 131486 397352
rect 131542 397296 131547 397352
rect 129968 397294 131547 397296
rect 131481 397291 131547 397294
rect 188981 397354 189047 397357
rect 188981 397352 190164 397354
rect 188981 397296 188986 397352
rect 189042 397296 190164 397352
rect 188981 397294 190164 397296
rect 188981 397291 189047 397294
rect 131297 396810 131363 396813
rect 129968 396808 131363 396810
rect 129968 396752 131302 396808
rect 131358 396752 131363 396808
rect 129968 396750 131363 396752
rect 131297 396747 131363 396750
rect 411989 396402 412055 396405
rect 409860 396400 412055 396402
rect 409860 396344 411994 396400
rect 412050 396344 412055 396400
rect 409860 396342 412055 396344
rect 411989 396339 412055 396342
rect 131205 396266 131271 396269
rect 129968 396264 131271 396266
rect 129968 396208 131210 396264
rect 131266 396208 131271 396264
rect 129968 396206 131271 396208
rect 131205 396203 131271 396206
rect 187325 396266 187391 396269
rect 187325 396264 190164 396266
rect 187325 396208 187330 396264
rect 187386 396208 190164 396264
rect 187325 396206 190164 396208
rect 187325 396203 187391 396206
rect 436737 396130 436803 396133
rect 436737 396128 440036 396130
rect 436737 396072 436742 396128
rect 436798 396072 440036 396128
rect 436737 396070 440036 396072
rect 436737 396067 436803 396070
rect 131205 395586 131271 395589
rect 129968 395584 131271 395586
rect 129968 395528 131210 395584
rect 131266 395528 131271 395584
rect 129968 395526 131271 395528
rect 131205 395523 131271 395526
rect 186313 395314 186379 395317
rect 186313 395312 190164 395314
rect 186313 395256 186318 395312
rect 186374 395256 190164 395312
rect 186313 395254 190164 395256
rect 186313 395251 186379 395254
rect 131297 395042 131363 395045
rect 129968 395040 131363 395042
rect 129968 394984 131302 395040
rect 131358 394984 131363 395040
rect 129968 394982 131363 394984
rect 131297 394979 131363 394982
rect 131205 394498 131271 394501
rect 129968 394496 131271 394498
rect 129968 394440 131210 394496
rect 131266 394440 131271 394496
rect 129968 394438 131271 394440
rect 131205 394435 131271 394438
rect 437565 394498 437631 394501
rect 437565 394496 440036 394498
rect 437565 394440 437570 394496
rect 437626 394440 440036 394496
rect 437565 394438 440036 394440
rect 437565 394435 437631 394438
rect 410425 394362 410491 394365
rect 409860 394360 410491 394362
rect 409860 394304 410430 394360
rect 410486 394304 410491 394360
rect 409860 394302 410491 394304
rect 410425 394299 410491 394302
rect 187141 394226 187207 394229
rect 187141 394224 190164 394226
rect 187141 394168 187146 394224
rect 187202 394168 190164 394224
rect 187141 394166 190164 394168
rect 187141 394163 187207 394166
rect 132033 393818 132099 393821
rect 129968 393816 132099 393818
rect 129968 393760 132038 393816
rect 132094 393760 132099 393816
rect 129968 393758 132099 393760
rect 132033 393755 132099 393758
rect 131205 393274 131271 393277
rect 129968 393272 131271 393274
rect 129968 393216 131210 393272
rect 131266 393216 131271 393272
rect 129968 393214 131271 393216
rect 131205 393211 131271 393214
rect 186313 393138 186379 393141
rect 186313 393136 190164 393138
rect 186313 393080 186318 393136
rect 186374 393080 190164 393136
rect 186313 393078 190164 393080
rect 186313 393075 186379 393078
rect 437473 392866 437539 392869
rect 437473 392864 440036 392866
rect 437473 392808 437478 392864
rect 437534 392808 440036 392864
rect 437473 392806 440036 392808
rect 437473 392803 437539 392806
rect 132033 392730 132099 392733
rect 129968 392728 132099 392730
rect 129968 392672 132038 392728
rect 132094 392672 132099 392728
rect 129968 392670 132099 392672
rect 132033 392667 132099 392670
rect 410425 392322 410491 392325
rect 409860 392320 410491 392322
rect 409860 392264 410430 392320
rect 410486 392264 410491 392320
rect 409860 392262 410491 392264
rect 410425 392259 410491 392262
rect 131297 392186 131363 392189
rect 129968 392184 131363 392186
rect 129968 392128 131302 392184
rect 131358 392128 131363 392184
rect 129968 392126 131363 392128
rect 131297 392123 131363 392126
rect 189073 392050 189139 392053
rect 189073 392048 190164 392050
rect 189073 391992 189078 392048
rect 189134 391992 190164 392048
rect 189073 391990 190164 391992
rect 189073 391987 189139 391990
rect 583520 391628 584960 391868
rect 131205 391506 131271 391509
rect 129968 391504 131271 391506
rect 129968 391448 131210 391504
rect 131266 391448 131271 391504
rect 129968 391446 131271 391448
rect 131205 391443 131271 391446
rect 437473 391234 437539 391237
rect 437473 391232 440036 391234
rect 437473 391176 437478 391232
rect 437534 391176 440036 391232
rect 437473 391174 440036 391176
rect 437473 391171 437539 391174
rect 186313 391098 186379 391101
rect 186313 391096 190164 391098
rect 186313 391040 186318 391096
rect 186374 391040 190164 391096
rect 186313 391038 190164 391040
rect 186313 391035 186379 391038
rect 131481 390962 131547 390965
rect 129968 390960 131547 390962
rect 129968 390904 131486 390960
rect 131542 390904 131547 390960
rect 129968 390902 131547 390904
rect 131481 390899 131547 390902
rect 131113 390418 131179 390421
rect 129968 390416 131179 390418
rect 129968 390360 131118 390416
rect 131174 390360 131179 390416
rect 129968 390358 131179 390360
rect 131113 390355 131179 390358
rect 411989 390282 412055 390285
rect 409860 390280 412055 390282
rect 409860 390224 411994 390280
rect 412050 390224 412055 390280
rect 409860 390222 412055 390224
rect 411989 390219 412055 390222
rect 187233 390010 187299 390013
rect 187233 390008 190164 390010
rect 187233 389952 187238 390008
rect 187294 389952 190164 390008
rect 187233 389950 190164 389952
rect 187233 389947 187299 389950
rect 131481 389874 131547 389877
rect 129968 389872 131547 389874
rect 129968 389816 131486 389872
rect 131542 389816 131547 389872
rect 129968 389814 131547 389816
rect 131481 389811 131547 389814
rect 437749 389602 437815 389605
rect 437749 389600 440036 389602
rect 437749 389544 437754 389600
rect 437810 389544 440036 389600
rect 437749 389542 440036 389544
rect 437749 389539 437815 389542
rect 552289 389330 552355 389333
rect 549884 389328 552355 389330
rect 549884 389272 552294 389328
rect 552350 389272 552355 389328
rect 549884 389270 552355 389272
rect 552289 389267 552355 389270
rect 131205 389194 131271 389197
rect 129968 389192 131271 389194
rect 129968 389136 131210 389192
rect 131266 389136 131271 389192
rect 129968 389134 131271 389136
rect 131205 389131 131271 389134
rect 186313 388922 186379 388925
rect 186313 388920 190164 388922
rect 186313 388864 186318 388920
rect 186374 388864 190164 388920
rect 186313 388862 190164 388864
rect 186313 388859 186379 388862
rect 131297 388650 131363 388653
rect 129968 388648 131363 388650
rect 129968 388592 131302 388648
rect 131358 388592 131363 388648
rect 129968 388590 131363 388592
rect 131297 388587 131363 388590
rect 411897 388242 411963 388245
rect 409860 388240 411963 388242
rect 409860 388184 411902 388240
rect 411958 388184 411963 388240
rect 409860 388182 411963 388184
rect 411897 388179 411963 388182
rect 131205 388106 131271 388109
rect 129968 388104 131271 388106
rect 129968 388048 131210 388104
rect 131266 388048 131271 388104
rect 129968 388046 131271 388048
rect 131205 388043 131271 388046
rect 186405 387970 186471 387973
rect 186405 387968 190164 387970
rect 186405 387912 186410 387968
rect 186466 387912 190164 387968
rect 186405 387910 190164 387912
rect 186405 387907 186471 387910
rect 438301 387834 438367 387837
rect 438301 387832 440036 387834
rect 438301 387776 438306 387832
rect 438362 387776 440036 387832
rect 438301 387774 440036 387776
rect 438301 387771 438367 387774
rect 131113 387426 131179 387429
rect 129968 387424 131179 387426
rect 129968 387368 131118 387424
rect 131174 387368 131179 387424
rect 129968 387366 131179 387368
rect 131113 387363 131179 387366
rect 131205 386882 131271 386885
rect 129968 386880 131271 386882
rect 129968 386824 131210 386880
rect 131266 386824 131271 386880
rect 129968 386822 131271 386824
rect 131205 386819 131271 386822
rect 187325 386882 187391 386885
rect 187325 386880 190164 386882
rect 187325 386824 187330 386880
rect 187386 386824 190164 386880
rect 187325 386822 190164 386824
rect 187325 386819 187391 386822
rect 131297 386338 131363 386341
rect 129968 386336 131363 386338
rect 129968 386280 131302 386336
rect 131358 386280 131363 386336
rect 129968 386278 131363 386280
rect 131297 386275 131363 386278
rect 438393 386202 438459 386205
rect 438393 386200 440036 386202
rect 438393 386144 438398 386200
rect 438454 386144 440036 386200
rect 438393 386142 440036 386144
rect 438393 386139 438459 386142
rect 411805 386066 411871 386069
rect 409860 386064 411871 386066
rect 409860 386008 411810 386064
rect 411866 386008 411871 386064
rect 409860 386006 411871 386008
rect 411805 386003 411871 386006
rect 131113 385794 131179 385797
rect 129968 385792 131179 385794
rect 129968 385736 131118 385792
rect 131174 385736 131179 385792
rect 129968 385734 131179 385736
rect 131113 385731 131179 385734
rect 186313 385794 186379 385797
rect 186313 385792 190164 385794
rect 186313 385736 186318 385792
rect 186374 385736 190164 385792
rect 186313 385734 190164 385736
rect 186313 385731 186379 385734
rect 131205 385114 131271 385117
rect 129968 385112 131271 385114
rect 129968 385056 131210 385112
rect 131266 385056 131271 385112
rect 129968 385054 131271 385056
rect 131205 385051 131271 385054
rect 187417 384706 187483 384709
rect 187417 384704 190164 384706
rect 187417 384648 187422 384704
rect 187478 384648 190164 384704
rect 187417 384646 190164 384648
rect 187417 384643 187483 384646
rect 131113 384570 131179 384573
rect 129968 384568 131179 384570
rect -960 384284 480 384524
rect 129968 384512 131118 384568
rect 131174 384512 131179 384568
rect 129968 384510 131179 384512
rect 131113 384507 131179 384510
rect 437473 384570 437539 384573
rect 437473 384568 440036 384570
rect 437473 384512 437478 384568
rect 437534 384512 440036 384568
rect 437473 384510 440036 384512
rect 437473 384507 437539 384510
rect 131205 384026 131271 384029
rect 411805 384026 411871 384029
rect 129968 384024 131271 384026
rect 129968 383968 131210 384024
rect 131266 383968 131271 384024
rect 129968 383966 131271 383968
rect 409860 384024 411871 384026
rect 409860 383968 411810 384024
rect 411866 383968 411871 384024
rect 409860 383966 411871 383968
rect 131205 383963 131271 383966
rect 411805 383963 411871 383966
rect 131113 383482 131179 383485
rect 129968 383480 131179 383482
rect 129968 383424 131118 383480
rect 131174 383424 131179 383480
rect 129968 383422 131179 383424
rect 131113 383419 131179 383422
rect 437933 382938 437999 382941
rect 437933 382936 440036 382938
rect 437933 382880 437938 382936
rect 437994 382880 440036 382936
rect 437933 382878 440036 382880
rect 437933 382875 437999 382878
rect 131205 382802 131271 382805
rect 129968 382800 131271 382802
rect 129968 382744 131210 382800
rect 131266 382744 131271 382800
rect 129968 382742 131271 382744
rect 131205 382739 131271 382742
rect 189073 382666 189139 382669
rect 189073 382664 190164 382666
rect 189073 382608 189078 382664
rect 189134 382608 190164 382664
rect 189073 382606 190164 382608
rect 189073 382603 189139 382606
rect 131481 382258 131547 382261
rect 129968 382256 131547 382258
rect 129968 382200 131486 382256
rect 131542 382200 131547 382256
rect 129968 382198 131547 382200
rect 131481 382195 131547 382198
rect 411713 381986 411779 381989
rect 409860 381984 411779 381986
rect 409860 381928 411718 381984
rect 411774 381928 411779 381984
rect 409860 381926 411779 381928
rect 411713 381923 411779 381926
rect 132217 381714 132283 381717
rect 129968 381712 132283 381714
rect 129968 381656 132222 381712
rect 132278 381656 132283 381712
rect 129968 381654 132283 381656
rect 132217 381651 132283 381654
rect 187233 381578 187299 381581
rect 187233 381576 190164 381578
rect 187233 381520 187238 381576
rect 187294 381520 190164 381576
rect 187233 381518 190164 381520
rect 187233 381515 187299 381518
rect 437473 381306 437539 381309
rect 437473 381304 440036 381306
rect 437473 381248 437478 381304
rect 437534 381248 440036 381304
rect 437473 381246 440036 381248
rect 437473 381243 437539 381246
rect 131205 381034 131271 381037
rect 129968 381032 131271 381034
rect 129968 380976 131210 381032
rect 131266 380976 131271 381032
rect 129968 380974 131271 380976
rect 131205 380971 131271 380974
rect 131205 380490 131271 380493
rect 129968 380488 131271 380490
rect 129968 380432 131210 380488
rect 131266 380432 131271 380488
rect 129968 380430 131271 380432
rect 131205 380427 131271 380430
rect 187141 380490 187207 380493
rect 187141 380488 190164 380490
rect 187141 380432 187146 380488
rect 187202 380432 190164 380488
rect 187141 380430 190164 380432
rect 187141 380427 187207 380430
rect 131481 379946 131547 379949
rect 412173 379946 412239 379949
rect 129968 379944 131547 379946
rect 129968 379888 131486 379944
rect 131542 379888 131547 379944
rect 129968 379886 131547 379888
rect 409860 379944 412239 379946
rect 409860 379888 412178 379944
rect 412234 379888 412239 379944
rect 409860 379886 412239 379888
rect 131481 379883 131547 379886
rect 412173 379883 412239 379886
rect 437473 379674 437539 379677
rect 437473 379672 440036 379674
rect 437473 379616 437478 379672
rect 437534 379616 440036 379672
rect 437473 379614 440036 379616
rect 437473 379611 437539 379614
rect 186405 379538 186471 379541
rect 186405 379536 190164 379538
rect 186405 379480 186410 379536
rect 186466 379480 190164 379536
rect 186405 379478 190164 379480
rect 186405 379475 186471 379478
rect 131113 379402 131179 379405
rect 129968 379400 131179 379402
rect 129968 379344 131118 379400
rect 131174 379344 131179 379400
rect 129968 379342 131179 379344
rect 131113 379339 131179 379342
rect 131297 378722 131363 378725
rect 129968 378720 131363 378722
rect 129968 378664 131302 378720
rect 131358 378664 131363 378720
rect 129968 378662 131363 378664
rect 131297 378659 131363 378662
rect 186313 378450 186379 378453
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 186313 378448 190164 378450
rect 186313 378392 186318 378448
rect 186374 378392 190164 378448
rect 186313 378390 190164 378392
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 186313 378387 186379 378390
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 131205 378178 131271 378181
rect 129968 378176 131271 378178
rect 129968 378120 131210 378176
rect 131266 378120 131271 378176
rect 129968 378118 131271 378120
rect 131205 378115 131271 378118
rect 437473 378042 437539 378045
rect 437473 378040 440036 378042
rect 437473 377984 437478 378040
rect 437534 377984 440036 378040
rect 437473 377982 440036 377984
rect 437473 377979 437539 377982
rect 131113 377634 131179 377637
rect 129968 377632 131179 377634
rect 129968 377576 131118 377632
rect 131174 377576 131179 377632
rect 129968 377574 131179 377576
rect 131113 377571 131179 377574
rect 186313 377362 186379 377365
rect 409830 377362 409890 377876
rect 410006 377362 410012 377364
rect 186313 377360 190164 377362
rect 186313 377304 186318 377360
rect 186374 377304 190164 377360
rect 186313 377302 190164 377304
rect 409830 377302 410012 377362
rect 186313 377299 186379 377302
rect 410006 377300 410012 377302
rect 410076 377300 410082 377364
rect 131205 377090 131271 377093
rect 129968 377088 131271 377090
rect 129968 377032 131210 377088
rect 131266 377032 131271 377088
rect 129968 377030 131271 377032
rect 131205 377027 131271 377030
rect 131205 376410 131271 376413
rect 129968 376408 131271 376410
rect 129968 376352 131210 376408
rect 131266 376352 131271 376408
rect 129968 376350 131271 376352
rect 131205 376347 131271 376350
rect 437473 376410 437539 376413
rect 437473 376408 440036 376410
rect 437473 376352 437478 376408
rect 437534 376352 440036 376408
rect 437473 376350 440036 376352
rect 437473 376347 437539 376350
rect 186313 376274 186379 376277
rect 186313 376272 190164 376274
rect 186313 376216 186318 376272
rect 186374 376216 190164 376272
rect 186313 376214 190164 376216
rect 186313 376211 186379 376214
rect 131481 375866 131547 375869
rect 411805 375866 411871 375869
rect 129968 375864 131547 375866
rect 129968 375808 131486 375864
rect 131542 375808 131547 375864
rect 129968 375806 131547 375808
rect 409860 375864 411871 375866
rect 409860 375808 411810 375864
rect 411866 375808 411871 375864
rect 409860 375806 411871 375808
rect 131481 375803 131547 375806
rect 411805 375803 411871 375806
rect 552197 375594 552263 375597
rect 549884 375592 552263 375594
rect 549884 375536 552202 375592
rect 552258 375536 552263 375592
rect 549884 375534 552263 375536
rect 552197 375531 552263 375534
rect 131205 375322 131271 375325
rect 129968 375320 131271 375322
rect 129968 375264 131210 375320
rect 131266 375264 131271 375320
rect 129968 375262 131271 375264
rect 131205 375259 131271 375262
rect 186405 375322 186471 375325
rect 186405 375320 190164 375322
rect 186405 375264 186410 375320
rect 186466 375264 190164 375320
rect 186405 375262 190164 375264
rect 186405 375259 186471 375262
rect 437473 374778 437539 374781
rect 437473 374776 440036 374778
rect 437473 374720 437478 374776
rect 437534 374720 440036 374776
rect 437473 374718 440036 374720
rect 437473 374715 437539 374718
rect 131113 374642 131179 374645
rect 129968 374640 131179 374642
rect 129968 374584 131118 374640
rect 131174 374584 131179 374640
rect 129968 374582 131179 374584
rect 131113 374579 131179 374582
rect 186313 374234 186379 374237
rect 186313 374232 190164 374234
rect 186313 374176 186318 374232
rect 186374 374176 190164 374232
rect 186313 374174 190164 374176
rect 186313 374171 186379 374174
rect 131205 374098 131271 374101
rect 129968 374096 131271 374098
rect 129968 374040 131210 374096
rect 131266 374040 131271 374096
rect 129968 374038 131271 374040
rect 131205 374035 131271 374038
rect 410517 373826 410583 373829
rect 409860 373824 410583 373826
rect 409860 373768 410522 373824
rect 410578 373768 410583 373824
rect 409860 373766 410583 373768
rect 410517 373763 410583 373766
rect 131205 373554 131271 373557
rect 129968 373552 131271 373554
rect 129968 373496 131210 373552
rect 131266 373496 131271 373552
rect 129968 373494 131271 373496
rect 131205 373491 131271 373494
rect 186313 373146 186379 373149
rect 437013 373146 437079 373149
rect 186313 373144 190164 373146
rect 186313 373088 186318 373144
rect 186374 373088 190164 373144
rect 186313 373086 190164 373088
rect 437013 373144 440036 373146
rect 437013 373088 437018 373144
rect 437074 373088 440036 373144
rect 437013 373086 440036 373088
rect 186313 373083 186379 373086
rect 437013 373083 437079 373086
rect 131481 373010 131547 373013
rect 129968 373008 131547 373010
rect 129968 372952 131486 373008
rect 131542 372952 131547 373008
rect 129968 372950 131547 372952
rect 131481 372947 131547 372950
rect 131113 372330 131179 372333
rect 129968 372328 131179 372330
rect 129968 372272 131118 372328
rect 131174 372272 131179 372328
rect 129968 372270 131179 372272
rect 131113 372267 131179 372270
rect 186313 372058 186379 372061
rect 186313 372056 190164 372058
rect 186313 372000 186318 372056
rect 186374 372000 190164 372056
rect 186313 371998 190164 372000
rect 186313 371995 186379 371998
rect 131205 371786 131271 371789
rect 411253 371786 411319 371789
rect 129968 371784 131271 371786
rect 129968 371728 131210 371784
rect 131266 371728 131271 371784
rect 129968 371726 131271 371728
rect 409860 371784 411319 371786
rect 409860 371728 411258 371784
rect 411314 371728 411319 371784
rect 409860 371726 411319 371728
rect 131205 371723 131271 371726
rect 411253 371723 411319 371726
rect 437473 371514 437539 371517
rect 437473 371512 440036 371514
rect -960 371228 480 371468
rect 437473 371456 437478 371512
rect 437534 371456 440036 371512
rect 437473 371454 440036 371456
rect 437473 371451 437539 371454
rect 131941 371242 132007 371245
rect 129968 371240 132007 371242
rect 129968 371184 131946 371240
rect 132002 371184 132007 371240
rect 129968 371182 132007 371184
rect 131941 371179 132007 371182
rect 186313 371106 186379 371109
rect 186313 371104 190164 371106
rect 186313 371048 186318 371104
rect 186374 371048 190164 371104
rect 186313 371046 190164 371048
rect 186313 371043 186379 371046
rect 131113 370698 131179 370701
rect 129968 370696 131179 370698
rect 129968 370640 131118 370696
rect 131174 370640 131179 370696
rect 129968 370638 131179 370640
rect 131113 370635 131179 370638
rect 131205 370018 131271 370021
rect 129968 370016 131271 370018
rect 129968 369960 131210 370016
rect 131266 369960 131271 370016
rect 129968 369958 131271 369960
rect 131205 369955 131271 369958
rect 186405 370018 186471 370021
rect 186405 370016 190164 370018
rect 186405 369960 186410 370016
rect 186466 369960 190164 370016
rect 186405 369958 190164 369960
rect 186405 369955 186471 369958
rect 437473 369882 437539 369885
rect 437473 369880 440036 369882
rect 437473 369824 437478 369880
rect 437534 369824 440036 369880
rect 437473 369822 440036 369824
rect 437473 369819 437539 369822
rect 410241 369610 410307 369613
rect 409860 369608 410307 369610
rect 409860 369552 410246 369608
rect 410302 369552 410307 369608
rect 409860 369550 410307 369552
rect 410241 369547 410307 369550
rect 131205 369474 131271 369477
rect 129968 369472 131271 369474
rect 129968 369416 131210 369472
rect 131266 369416 131271 369472
rect 129968 369414 131271 369416
rect 131205 369411 131271 369414
rect 131481 368930 131547 368933
rect 129968 368928 131547 368930
rect 129968 368872 131486 368928
rect 131542 368872 131547 368928
rect 129968 368870 131547 368872
rect 131481 368867 131547 368870
rect 186313 368930 186379 368933
rect 186313 368928 190164 368930
rect 186313 368872 186318 368928
rect 186374 368872 190164 368928
rect 186313 368870 190164 368872
rect 186313 368867 186379 368870
rect 131205 368250 131271 368253
rect 129968 368248 131271 368250
rect 129968 368192 131210 368248
rect 131266 368192 131271 368248
rect 129968 368190 131271 368192
rect 131205 368187 131271 368190
rect 437473 368250 437539 368253
rect 437473 368248 440036 368250
rect 437473 368192 437478 368248
rect 437534 368192 440036 368248
rect 437473 368190 440036 368192
rect 437473 368187 437539 368190
rect 186313 367842 186379 367845
rect 186313 367840 190164 367842
rect 186313 367784 186318 367840
rect 186374 367784 190164 367840
rect 186313 367782 190164 367784
rect 186313 367779 186379 367782
rect 131113 367706 131179 367709
rect 129968 367704 131179 367706
rect 129968 367648 131118 367704
rect 131174 367648 131179 367704
rect 129968 367646 131179 367648
rect 131113 367643 131179 367646
rect 412265 367570 412331 367573
rect 409860 367568 412331 367570
rect 409860 367512 412270 367568
rect 412326 367512 412331 367568
rect 409860 367510 412331 367512
rect 412265 367507 412331 367510
rect 131205 367162 131271 367165
rect 129968 367160 131271 367162
rect 129968 367104 131210 367160
rect 131266 367104 131271 367160
rect 129968 367102 131271 367104
rect 131205 367099 131271 367102
rect 186313 366890 186379 366893
rect 186313 366888 190164 366890
rect 186313 366832 186318 366888
rect 186374 366832 190164 366888
rect 186313 366830 190164 366832
rect 186313 366827 186379 366830
rect 132217 366618 132283 366621
rect 129968 366616 132283 366618
rect 129968 366560 132222 366616
rect 132278 366560 132283 366616
rect 129968 366558 132283 366560
rect 132217 366555 132283 366558
rect 437473 366482 437539 366485
rect 437473 366480 440036 366482
rect 437473 366424 437478 366480
rect 437534 366424 440036 366480
rect 437473 366422 440036 366424
rect 437473 366419 437539 366422
rect 131205 365938 131271 365941
rect 129968 365936 131271 365938
rect 129968 365880 131210 365936
rect 131266 365880 131271 365936
rect 129968 365878 131271 365880
rect 131205 365875 131271 365878
rect 186405 365802 186471 365805
rect 186405 365800 190164 365802
rect 186405 365744 186410 365800
rect 186466 365744 190164 365800
rect 186405 365742 190164 365744
rect 186405 365739 186471 365742
rect 411253 365530 411319 365533
rect 409860 365528 411319 365530
rect 409860 365472 411258 365528
rect 411314 365472 411319 365528
rect 409860 365470 411319 365472
rect 411253 365467 411319 365470
rect 131113 365394 131179 365397
rect 129968 365392 131179 365394
rect 129968 365336 131118 365392
rect 131174 365336 131179 365392
rect 129968 365334 131179 365336
rect 131113 365331 131179 365334
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect 131205 364850 131271 364853
rect 129968 364848 131271 364850
rect 129968 364792 131210 364848
rect 131266 364792 131271 364848
rect 129968 364790 131271 364792
rect 131205 364787 131271 364790
rect 437473 364850 437539 364853
rect 437473 364848 440036 364850
rect 437473 364792 437478 364848
rect 437534 364792 440036 364848
rect 437473 364790 440036 364792
rect 437473 364787 437539 364790
rect 186313 364714 186379 364717
rect 186313 364712 190164 364714
rect 186313 364656 186318 364712
rect 186374 364656 190164 364712
rect 186313 364654 190164 364656
rect 186313 364651 186379 364654
rect 131481 364306 131547 364309
rect 129968 364304 131547 364306
rect 129968 364248 131486 364304
rect 131542 364248 131547 364304
rect 129968 364246 131547 364248
rect 131481 364243 131547 364246
rect 131113 363626 131179 363629
rect 129968 363624 131179 363626
rect 129968 363568 131118 363624
rect 131174 363568 131179 363624
rect 129968 363566 131179 363568
rect 131113 363563 131179 363566
rect 186313 363626 186379 363629
rect 186313 363624 190164 363626
rect 186313 363568 186318 363624
rect 186374 363568 190164 363624
rect 186313 363566 190164 363568
rect 186313 363563 186379 363566
rect 410149 363490 410215 363493
rect 409860 363488 410215 363490
rect 409860 363432 410154 363488
rect 410210 363432 410215 363488
rect 409860 363430 410215 363432
rect 410149 363427 410215 363430
rect 437473 363218 437539 363221
rect 437473 363216 440036 363218
rect 437473 363160 437478 363216
rect 437534 363160 440036 363216
rect 437473 363158 440036 363160
rect 437473 363155 437539 363158
rect 131205 363082 131271 363085
rect 129968 363080 131271 363082
rect 129968 363024 131210 363080
rect 131266 363024 131271 363080
rect 129968 363022 131271 363024
rect 131205 363019 131271 363022
rect 186313 362674 186379 362677
rect 186313 362672 190164 362674
rect 186313 362616 186318 362672
rect 186374 362616 190164 362672
rect 186313 362614 190164 362616
rect 186313 362611 186379 362614
rect 131113 362538 131179 362541
rect 129968 362536 131179 362538
rect 129968 362480 131118 362536
rect 131174 362480 131179 362536
rect 129968 362478 131179 362480
rect 131113 362475 131179 362478
rect 131205 361858 131271 361861
rect 552013 361858 552079 361861
rect 129968 361856 131271 361858
rect 129968 361800 131210 361856
rect 131266 361800 131271 361856
rect 129968 361798 131271 361800
rect 549884 361856 552079 361858
rect 549884 361800 552018 361856
rect 552074 361800 552079 361856
rect 549884 361798 552079 361800
rect 131205 361795 131271 361798
rect 552013 361795 552079 361798
rect 186313 361586 186379 361589
rect 437473 361586 437539 361589
rect 186313 361584 190164 361586
rect 186313 361528 186318 361584
rect 186374 361528 190164 361584
rect 186313 361526 190164 361528
rect 437473 361584 440036 361586
rect 437473 361528 437478 361584
rect 437534 361528 440036 361584
rect 437473 361526 440036 361528
rect 186313 361523 186379 361526
rect 437473 361523 437539 361526
rect 412541 361450 412607 361453
rect 409860 361448 412607 361450
rect 409860 361392 412546 361448
rect 412602 361392 412607 361448
rect 409860 361390 412607 361392
rect 412541 361387 412607 361390
rect 131113 361314 131179 361317
rect 129968 361312 131179 361314
rect 129968 361256 131118 361312
rect 131174 361256 131179 361312
rect 129968 361254 131179 361256
rect 131113 361251 131179 361254
rect 132125 360770 132191 360773
rect 129968 360768 132191 360770
rect 129968 360712 132130 360768
rect 132186 360712 132191 360768
rect 129968 360710 132191 360712
rect 132125 360707 132191 360710
rect 186405 360498 186471 360501
rect 186405 360496 190164 360498
rect 186405 360440 186410 360496
rect 186466 360440 190164 360496
rect 186405 360438 190164 360440
rect 186405 360435 186471 360438
rect 131205 360226 131271 360229
rect 129968 360224 131271 360226
rect 129968 360168 131210 360224
rect 131266 360168 131271 360224
rect 129968 360166 131271 360168
rect 131205 360163 131271 360166
rect 436921 359954 436987 359957
rect 436921 359952 440036 359954
rect 436921 359896 436926 359952
rect 436982 359896 440036 359952
rect 436921 359894 440036 359896
rect 436921 359891 436987 359894
rect 132033 359546 132099 359549
rect 129968 359544 132099 359546
rect 129968 359488 132038 359544
rect 132094 359488 132099 359544
rect 129968 359486 132099 359488
rect 132033 359483 132099 359486
rect 186313 359410 186379 359413
rect 411253 359410 411319 359413
rect 186313 359408 190164 359410
rect 186313 359352 186318 359408
rect 186374 359352 190164 359408
rect 186313 359350 190164 359352
rect 409860 359408 411319 359410
rect 409860 359352 411258 359408
rect 411314 359352 411319 359408
rect 409860 359350 411319 359352
rect 186313 359347 186379 359350
rect 411253 359347 411319 359350
rect 131205 359002 131271 359005
rect 129968 359000 131271 359002
rect 129968 358944 131210 359000
rect 131266 358944 131271 359000
rect 129968 358942 131271 358944
rect 131205 358939 131271 358942
rect -960 358308 480 358548
rect 131113 358458 131179 358461
rect 129968 358456 131179 358458
rect 129968 358400 131118 358456
rect 131174 358400 131179 358456
rect 129968 358398 131179 358400
rect 131113 358395 131179 358398
rect 187417 358458 187483 358461
rect 187417 358456 190164 358458
rect 187417 358400 187422 358456
rect 187478 358400 190164 358456
rect 187417 358398 190164 358400
rect 187417 358395 187483 358398
rect 437473 358322 437539 358325
rect 437473 358320 440036 358322
rect 437473 358264 437478 358320
rect 437534 358264 440036 358320
rect 437473 358262 440036 358264
rect 437473 358259 437539 358262
rect 131205 357914 131271 357917
rect 129968 357912 131271 357914
rect 129968 357856 131210 357912
rect 131266 357856 131271 357912
rect 129968 357854 131271 357856
rect 131205 357851 131271 357854
rect 186313 357370 186379 357373
rect 411345 357370 411411 357373
rect 186313 357368 190164 357370
rect 186313 357312 186318 357368
rect 186374 357312 190164 357368
rect 186313 357310 190164 357312
rect 409860 357368 411411 357370
rect 409860 357312 411350 357368
rect 411406 357312 411411 357368
rect 409860 357310 411411 357312
rect 186313 357307 186379 357310
rect 411345 357307 411411 357310
rect 131297 357234 131363 357237
rect 129968 357232 131363 357234
rect 129968 357176 131302 357232
rect 131358 357176 131363 357232
rect 129968 357174 131363 357176
rect 131297 357171 131363 357174
rect 131113 356690 131179 356693
rect 129968 356688 131179 356690
rect 129968 356632 131118 356688
rect 131174 356632 131179 356688
rect 129968 356630 131179 356632
rect 131113 356627 131179 356630
rect 437473 356690 437539 356693
rect 437473 356688 440036 356690
rect 437473 356632 437478 356688
rect 437534 356632 440036 356688
rect 437473 356630 440036 356632
rect 437473 356627 437539 356630
rect 186405 356282 186471 356285
rect 186405 356280 190164 356282
rect 186405 356224 186410 356280
rect 186466 356224 190164 356280
rect 186405 356222 190164 356224
rect 186405 356219 186471 356222
rect 131205 356146 131271 356149
rect 129968 356144 131271 356146
rect 129968 356088 131210 356144
rect 131266 356088 131271 356144
rect 129968 356086 131271 356088
rect 131205 356083 131271 356086
rect 409873 355874 409939 355877
rect 409830 355872 409939 355874
rect 409830 355816 409878 355872
rect 409934 355816 409939 355872
rect 409830 355811 409939 355816
rect 131297 355466 131363 355469
rect 129968 355464 131363 355466
rect 129968 355408 131302 355464
rect 131358 355408 131363 355464
rect 129968 355406 131363 355408
rect 131297 355403 131363 355406
rect 186313 355330 186379 355333
rect 186313 355328 190164 355330
rect 186313 355272 186318 355328
rect 186374 355272 190164 355328
rect 409830 355300 409890 355811
rect 186313 355270 190164 355272
rect 186313 355267 186379 355270
rect 437473 355058 437539 355061
rect 437473 355056 440036 355058
rect 437473 355000 437478 355056
rect 437534 355000 440036 355056
rect 437473 354998 440036 355000
rect 437473 354995 437539 354998
rect 131205 354922 131271 354925
rect 129968 354920 131271 354922
rect 129968 354864 131210 354920
rect 131266 354864 131271 354920
rect 129968 354862 131271 354864
rect 131205 354859 131271 354862
rect 131113 354378 131179 354381
rect 129968 354376 131179 354378
rect 129968 354320 131118 354376
rect 131174 354320 131179 354376
rect 129968 354318 131179 354320
rect 131113 354315 131179 354318
rect 186313 354242 186379 354245
rect 186313 354240 190164 354242
rect 186313 354184 186318 354240
rect 186374 354184 190164 354240
rect 186313 354182 190164 354184
rect 186313 354179 186379 354182
rect 131205 353834 131271 353837
rect 129968 353832 131271 353834
rect 129968 353776 131210 353832
rect 131266 353776 131271 353832
rect 129968 353774 131271 353776
rect 131205 353771 131271 353774
rect 437473 353426 437539 353429
rect 437473 353424 440036 353426
rect 437473 353368 437478 353424
rect 437534 353368 440036 353424
rect 437473 353366 440036 353368
rect 437473 353363 437539 353366
rect 131205 353154 131271 353157
rect 129968 353152 131271 353154
rect 129968 353096 131210 353152
rect 131266 353096 131271 353152
rect 129968 353094 131271 353096
rect 131205 353091 131271 353094
rect 186405 353154 186471 353157
rect 411253 353154 411319 353157
rect 186405 353152 190164 353154
rect 186405 353096 186410 353152
rect 186466 353096 190164 353152
rect 186405 353094 190164 353096
rect 409860 353152 411319 353154
rect 409860 353096 411258 353152
rect 411314 353096 411319 353152
rect 409860 353094 411319 353096
rect 186405 353091 186471 353094
rect 411253 353091 411319 353094
rect 131113 352610 131179 352613
rect 129968 352608 131179 352610
rect 129968 352552 131118 352608
rect 131174 352552 131179 352608
rect 129968 352550 131179 352552
rect 131113 352547 131179 352550
rect 131481 352066 131547 352069
rect 129968 352064 131547 352066
rect 129968 352008 131486 352064
rect 131542 352008 131547 352064
rect 129968 352006 131547 352008
rect 131481 352003 131547 352006
rect 186313 352066 186379 352069
rect 186313 352064 190164 352066
rect 186313 352008 186318 352064
rect 186374 352008 190164 352064
rect 186313 352006 190164 352008
rect 186313 352003 186379 352006
rect 437473 351794 437539 351797
rect 437473 351792 440036 351794
rect 437473 351736 437478 351792
rect 437534 351736 440036 351792
rect 583520 351780 584960 352020
rect 437473 351734 440036 351736
rect 437473 351731 437539 351734
rect 131113 351522 131179 351525
rect 129968 351520 131179 351522
rect 129968 351464 131118 351520
rect 131174 351464 131179 351520
rect 129968 351462 131179 351464
rect 131113 351459 131179 351462
rect 186313 351114 186379 351117
rect 411621 351114 411687 351117
rect 186313 351112 190164 351114
rect 186313 351056 186318 351112
rect 186374 351056 190164 351112
rect 186313 351054 190164 351056
rect 409860 351112 411687 351114
rect 409860 351056 411626 351112
rect 411682 351056 411687 351112
rect 409860 351054 411687 351056
rect 186313 351051 186379 351054
rect 411621 351051 411687 351054
rect 131205 350842 131271 350845
rect 129968 350840 131271 350842
rect 129968 350784 131210 350840
rect 131266 350784 131271 350840
rect 129968 350782 131271 350784
rect 131205 350779 131271 350782
rect 131113 350298 131179 350301
rect 129968 350296 131179 350298
rect 129968 350240 131118 350296
rect 131174 350240 131179 350296
rect 129968 350238 131179 350240
rect 131113 350235 131179 350238
rect 437473 350162 437539 350165
rect 437473 350160 440036 350162
rect 437473 350104 437478 350160
rect 437534 350104 440036 350160
rect 437473 350102 440036 350104
rect 437473 350099 437539 350102
rect 28901 350026 28967 350029
rect 186313 350026 186379 350029
rect 28901 350024 30084 350026
rect 28901 349968 28906 350024
rect 28962 349968 30084 350024
rect 28901 349966 30084 349968
rect 186313 350024 190164 350026
rect 186313 349968 186318 350024
rect 186374 349968 190164 350024
rect 186313 349966 190164 349968
rect 28901 349963 28967 349966
rect 186313 349963 186379 349966
rect 131205 349754 131271 349757
rect 129968 349752 131271 349754
rect 129968 349696 131210 349752
rect 131266 349696 131271 349752
rect 129968 349694 131271 349696
rect 131205 349691 131271 349694
rect 131205 349074 131271 349077
rect 410609 349074 410675 349077
rect 129968 349072 131271 349074
rect 129968 349016 131210 349072
rect 131266 349016 131271 349072
rect 129968 349014 131271 349016
rect 409860 349072 410675 349074
rect 409860 349016 410614 349072
rect 410670 349016 410675 349072
rect 409860 349014 410675 349016
rect 131205 349011 131271 349014
rect 410609 349011 410675 349014
rect 186405 348938 186471 348941
rect 186405 348936 190164 348938
rect 186405 348880 186410 348936
rect 186466 348880 190164 348936
rect 186405 348878 190164 348880
rect 186405 348875 186471 348878
rect 131297 348530 131363 348533
rect 129968 348528 131363 348530
rect 129968 348472 131302 348528
rect 131358 348472 131363 348528
rect 129968 348470 131363 348472
rect 131297 348467 131363 348470
rect 437473 348530 437539 348533
rect 437473 348528 440036 348530
rect 437473 348472 437478 348528
rect 437534 348472 440036 348528
rect 437473 348470 440036 348472
rect 437473 348467 437539 348470
rect 552197 348122 552263 348125
rect 549884 348120 552263 348122
rect 549884 348064 552202 348120
rect 552258 348064 552263 348120
rect 549884 348062 552263 348064
rect 552197 348059 552263 348062
rect 131481 347986 131547 347989
rect 129968 347984 131547 347986
rect 129968 347928 131486 347984
rect 131542 347928 131547 347984
rect 129968 347926 131547 347928
rect 131481 347923 131547 347926
rect 186313 347850 186379 347853
rect 186313 347848 190164 347850
rect 186313 347792 186318 347848
rect 186374 347792 190164 347848
rect 186313 347790 190164 347792
rect 186313 347787 186379 347790
rect 131113 347442 131179 347445
rect 129968 347440 131179 347442
rect 129968 347384 131118 347440
rect 131174 347384 131179 347440
rect 129968 347382 131179 347384
rect 131113 347379 131179 347382
rect 411437 347034 411503 347037
rect 409860 347032 411503 347034
rect 409860 346976 411442 347032
rect 411498 346976 411503 347032
rect 409860 346974 411503 346976
rect 411437 346971 411503 346974
rect 186313 346898 186379 346901
rect 437473 346898 437539 346901
rect 186313 346896 190164 346898
rect 186313 346840 186318 346896
rect 186374 346840 190164 346896
rect 186313 346838 190164 346840
rect 437473 346896 440036 346898
rect 437473 346840 437478 346896
rect 437534 346840 440036 346896
rect 437473 346838 440036 346840
rect 186313 346835 186379 346838
rect 437473 346835 437539 346838
rect 131205 346762 131271 346765
rect 129968 346760 131271 346762
rect 129968 346704 131210 346760
rect 131266 346704 131271 346760
rect 129968 346702 131271 346704
rect 131205 346699 131271 346702
rect 131205 346218 131271 346221
rect 129968 346216 131271 346218
rect 129968 346160 131210 346216
rect 131266 346160 131271 346216
rect 129968 346158 131271 346160
rect 131205 346155 131271 346158
rect 186313 345810 186379 345813
rect 186313 345808 190164 345810
rect 186313 345752 186318 345808
rect 186374 345752 190164 345808
rect 186313 345750 190164 345752
rect 186313 345747 186379 345750
rect 131113 345674 131179 345677
rect 129968 345672 131179 345674
rect 129968 345616 131118 345672
rect 131174 345616 131179 345672
rect 129968 345614 131179 345616
rect 131113 345611 131179 345614
rect -960 345252 480 345492
rect 437473 345266 437539 345269
rect 437473 345264 440036 345266
rect 437473 345208 437478 345264
rect 437534 345208 440036 345264
rect 437473 345206 440036 345208
rect 437473 345203 437539 345206
rect 131205 345130 131271 345133
rect 129968 345128 131271 345130
rect 129968 345072 131210 345128
rect 131266 345072 131271 345128
rect 129968 345070 131271 345072
rect 131205 345067 131271 345070
rect 411253 344994 411319 344997
rect 409860 344992 411319 344994
rect 409860 344936 411258 344992
rect 411314 344936 411319 344992
rect 409860 344934 411319 344936
rect 411253 344931 411319 344934
rect 186313 344722 186379 344725
rect 186313 344720 190164 344722
rect 186313 344664 186318 344720
rect 186374 344664 190164 344720
rect 186313 344662 190164 344664
rect 186313 344659 186379 344662
rect 131297 344450 131363 344453
rect 129968 344448 131363 344450
rect 129968 344392 131302 344448
rect 131358 344392 131363 344448
rect 129968 344390 131363 344392
rect 131297 344387 131363 344390
rect 131205 343906 131271 343909
rect 129968 343904 131271 343906
rect 129968 343848 131210 343904
rect 131266 343848 131271 343904
rect 129968 343846 131271 343848
rect 131205 343843 131271 343846
rect 186313 343634 186379 343637
rect 186313 343632 190164 343634
rect 186313 343576 186318 343632
rect 186374 343576 190164 343632
rect 186313 343574 190164 343576
rect 186313 343571 186379 343574
rect 437473 343498 437539 343501
rect 437473 343496 440036 343498
rect 437473 343440 437478 343496
rect 437534 343440 440036 343496
rect 437473 343438 440036 343440
rect 437473 343435 437539 343438
rect 131205 343362 131271 343365
rect 129968 343360 131271 343362
rect 129968 343304 131210 343360
rect 131266 343304 131271 343360
rect 129968 343302 131271 343304
rect 131205 343299 131271 343302
rect 411253 342954 411319 342957
rect 409860 342952 411319 342954
rect 409860 342896 411258 342952
rect 411314 342896 411319 342952
rect 409860 342894 411319 342896
rect 411253 342891 411319 342894
rect 131481 342682 131547 342685
rect 129968 342680 131547 342682
rect 129968 342624 131486 342680
rect 131542 342624 131547 342680
rect 129968 342622 131547 342624
rect 131481 342619 131547 342622
rect 186405 342682 186471 342685
rect 186405 342680 190164 342682
rect 186405 342624 186410 342680
rect 186466 342624 190164 342680
rect 186405 342622 190164 342624
rect 186405 342619 186471 342622
rect 131113 342138 131179 342141
rect 129968 342136 131179 342138
rect 129968 342080 131118 342136
rect 131174 342080 131179 342136
rect 129968 342078 131179 342080
rect 131113 342075 131179 342078
rect 438485 341866 438551 341869
rect 438485 341864 440036 341866
rect 438485 341808 438490 341864
rect 438546 341808 440036 341864
rect 438485 341806 440036 341808
rect 438485 341803 438551 341806
rect 131297 341594 131363 341597
rect 129968 341592 131363 341594
rect 129968 341536 131302 341592
rect 131358 341536 131363 341592
rect 129968 341534 131363 341536
rect 131297 341531 131363 341534
rect 186313 341594 186379 341597
rect 186313 341592 190164 341594
rect 186313 341536 186318 341592
rect 186374 341536 190164 341592
rect 186313 341534 190164 341536
rect 186313 341531 186379 341534
rect 131205 341050 131271 341053
rect 129968 341048 131271 341050
rect 129968 340992 131210 341048
rect 131266 340992 131271 341048
rect 129968 340990 131271 340992
rect 131205 340987 131271 340990
rect 411437 340914 411503 340917
rect 409860 340912 411503 340914
rect 409860 340856 411442 340912
rect 411498 340856 411503 340912
rect 409860 340854 411503 340856
rect 411437 340851 411503 340854
rect 186313 340506 186379 340509
rect 186313 340504 190164 340506
rect 186313 340448 186318 340504
rect 186374 340448 190164 340504
rect 186313 340446 190164 340448
rect 186313 340443 186379 340446
rect 131297 340370 131363 340373
rect 129968 340368 131363 340370
rect 129968 340312 131302 340368
rect 131358 340312 131363 340368
rect 129968 340310 131363 340312
rect 131297 340307 131363 340310
rect 437841 340234 437907 340237
rect 437841 340232 440036 340234
rect 437841 340176 437846 340232
rect 437902 340176 440036 340232
rect 437841 340174 440036 340176
rect 437841 340171 437907 340174
rect 131205 339826 131271 339829
rect 129968 339824 131271 339826
rect 129968 339768 131210 339824
rect 131266 339768 131271 339824
rect 129968 339766 131271 339768
rect 131205 339763 131271 339766
rect 186313 339418 186379 339421
rect 186313 339416 190164 339418
rect 186313 339360 186318 339416
rect 186374 339360 190164 339416
rect 186313 339358 190164 339360
rect 186313 339355 186379 339358
rect 131113 339282 131179 339285
rect 129968 339280 131179 339282
rect 129968 339224 131118 339280
rect 131174 339224 131179 339280
rect 129968 339222 131179 339224
rect 131113 339219 131179 339222
rect 410701 338874 410767 338877
rect 409860 338872 410767 338874
rect 409860 338816 410706 338872
rect 410762 338816 410767 338872
rect 409860 338814 410767 338816
rect 410701 338811 410767 338814
rect 131205 338738 131271 338741
rect 129968 338736 131271 338738
rect 129968 338680 131210 338736
rect 131266 338680 131271 338736
rect 129968 338678 131271 338680
rect 131205 338675 131271 338678
rect 437473 338602 437539 338605
rect 437473 338600 440036 338602
rect 437473 338544 437478 338600
rect 437534 338544 440036 338600
rect 437473 338542 440036 338544
rect 437473 338539 437539 338542
rect 186405 338466 186471 338469
rect 186405 338464 190164 338466
rect 186405 338408 186410 338464
rect 186466 338408 190164 338464
rect 583520 338452 584960 338692
rect 186405 338406 190164 338408
rect 186405 338403 186471 338406
rect 131481 338058 131547 338061
rect 129968 338056 131547 338058
rect 129968 338000 131486 338056
rect 131542 338000 131547 338056
rect 129968 337998 131547 338000
rect 131481 337995 131547 337998
rect 132033 337514 132099 337517
rect 129968 337512 132099 337514
rect 129968 337456 132038 337512
rect 132094 337456 132099 337512
rect 129968 337454 132099 337456
rect 132033 337451 132099 337454
rect 186313 337378 186379 337381
rect 186313 337376 190164 337378
rect 186313 337320 186318 337376
rect 186374 337320 190164 337376
rect 186313 337318 190164 337320
rect 186313 337315 186379 337318
rect 131205 336970 131271 336973
rect 129968 336968 131271 336970
rect 129968 336912 131210 336968
rect 131266 336912 131271 336968
rect 129968 336910 131271 336912
rect 131205 336907 131271 336910
rect 437473 336970 437539 336973
rect 437473 336968 440036 336970
rect 437473 336912 437478 336968
rect 437534 336912 440036 336968
rect 437473 336910 440036 336912
rect 437473 336907 437539 336910
rect 411253 336834 411319 336837
rect 409860 336832 411319 336834
rect 409860 336776 411258 336832
rect 411314 336776 411319 336832
rect 409860 336774 411319 336776
rect 411253 336771 411319 336774
rect 131113 336290 131179 336293
rect 129968 336288 131179 336290
rect 129968 336232 131118 336288
rect 131174 336232 131179 336288
rect 129968 336230 131179 336232
rect 131113 336227 131179 336230
rect 186313 336290 186379 336293
rect 186313 336288 190164 336290
rect 186313 336232 186318 336288
rect 186374 336232 190164 336288
rect 186313 336230 190164 336232
rect 186313 336227 186379 336230
rect 131205 335746 131271 335749
rect 129968 335744 131271 335746
rect 129968 335688 131210 335744
rect 131266 335688 131271 335744
rect 129968 335686 131271 335688
rect 131205 335683 131271 335686
rect 437565 335338 437631 335341
rect 437565 335336 440036 335338
rect 437565 335280 437570 335336
rect 437626 335280 440036 335336
rect 437565 335278 440036 335280
rect 437565 335275 437631 335278
rect 131205 335202 131271 335205
rect 129968 335200 131271 335202
rect 129968 335144 131210 335200
rect 131266 335144 131271 335200
rect 129968 335142 131271 335144
rect 131205 335139 131271 335142
rect 186313 335202 186379 335205
rect 186313 335200 190164 335202
rect 186313 335144 186318 335200
rect 186374 335144 190164 335200
rect 186313 335142 190164 335144
rect 186313 335139 186379 335142
rect 132217 334658 132283 334661
rect 412817 334658 412883 334661
rect 129968 334656 132283 334658
rect 129968 334600 132222 334656
rect 132278 334600 132283 334656
rect 129968 334598 132283 334600
rect 409860 334656 412883 334658
rect 409860 334600 412822 334656
rect 412878 334600 412883 334656
rect 409860 334598 412883 334600
rect 132217 334595 132283 334598
rect 412817 334595 412883 334598
rect 552013 334386 552079 334389
rect 549884 334384 552079 334386
rect 549884 334328 552018 334384
rect 552074 334328 552079 334384
rect 549884 334326 552079 334328
rect 552013 334323 552079 334326
rect 186405 334250 186471 334253
rect 186405 334248 190164 334250
rect 186405 334192 186410 334248
rect 186466 334192 190164 334248
rect 186405 334190 190164 334192
rect 186405 334187 186471 334190
rect 131113 333978 131179 333981
rect 129968 333976 131179 333978
rect 129968 333920 131118 333976
rect 131174 333920 131179 333976
rect 129968 333918 131179 333920
rect 131113 333915 131179 333918
rect 437473 333706 437539 333709
rect 437473 333704 440036 333706
rect 437473 333648 437478 333704
rect 437534 333648 440036 333704
rect 437473 333646 440036 333648
rect 437473 333643 437539 333646
rect 131297 333434 131363 333437
rect 129968 333432 131363 333434
rect 129968 333376 131302 333432
rect 131358 333376 131363 333432
rect 129968 333374 131363 333376
rect 131297 333371 131363 333374
rect 186313 333162 186379 333165
rect 410057 333162 410123 333165
rect 186313 333160 190164 333162
rect 186313 333104 186318 333160
rect 186374 333104 190164 333160
rect 186313 333102 190164 333104
rect 409830 333160 410123 333162
rect 409830 333104 410062 333160
rect 410118 333104 410123 333160
rect 409830 333102 410123 333104
rect 186313 333099 186379 333102
rect 131205 332890 131271 332893
rect 129968 332888 131271 332890
rect 129968 332832 131210 332888
rect 131266 332832 131271 332888
rect 129968 332830 131271 332832
rect 131205 332827 131271 332830
rect 409830 332588 409890 333102
rect 410057 333099 410123 333102
rect -960 332196 480 332436
rect 132217 332346 132283 332349
rect 129968 332344 132283 332346
rect 129968 332288 132222 332344
rect 132278 332288 132283 332344
rect 129968 332286 132283 332288
rect 132217 332283 132283 332286
rect 186313 332074 186379 332077
rect 437473 332074 437539 332077
rect 186313 332072 190164 332074
rect 186313 332016 186318 332072
rect 186374 332016 190164 332072
rect 186313 332014 190164 332016
rect 437473 332072 440036 332074
rect 437473 332016 437478 332072
rect 437534 332016 440036 332072
rect 437473 332014 440036 332016
rect 186313 332011 186379 332014
rect 437473 332011 437539 332014
rect 131481 331666 131547 331669
rect 129968 331664 131547 331666
rect 129968 331608 131486 331664
rect 131542 331608 131547 331664
rect 129968 331606 131547 331608
rect 131481 331603 131547 331606
rect 131113 331122 131179 331125
rect 129968 331120 131179 331122
rect 129968 331064 131118 331120
rect 131174 331064 131179 331120
rect 129968 331062 131179 331064
rect 131113 331059 131179 331062
rect 186313 330986 186379 330989
rect 186313 330984 190164 330986
rect 186313 330928 186318 330984
rect 186374 330928 190164 330984
rect 186313 330926 190164 330928
rect 186313 330923 186379 330926
rect 132217 330578 132283 330581
rect 411253 330578 411319 330581
rect 129968 330576 132283 330578
rect 129968 330520 132222 330576
rect 132278 330520 132283 330576
rect 129968 330518 132283 330520
rect 409860 330576 411319 330578
rect 409860 330520 411258 330576
rect 411314 330520 411319 330576
rect 409860 330518 411319 330520
rect 132217 330515 132283 330518
rect 411253 330515 411319 330518
rect 437473 330442 437539 330445
rect 437473 330440 440036 330442
rect 437473 330384 437478 330440
rect 437534 330384 440036 330440
rect 437473 330382 440036 330384
rect 437473 330379 437539 330382
rect 186405 330034 186471 330037
rect 186405 330032 190164 330034
rect 186405 329976 186410 330032
rect 186466 329976 190164 330032
rect 186405 329974 190164 329976
rect 186405 329971 186471 329974
rect 131205 329898 131271 329901
rect 129968 329896 131271 329898
rect 129968 329840 131210 329896
rect 131266 329840 131271 329896
rect 129968 329838 131271 329840
rect 131205 329835 131271 329838
rect 131205 329354 131271 329357
rect 129968 329352 131271 329354
rect 129968 329296 131210 329352
rect 131266 329296 131271 329352
rect 129968 329294 131271 329296
rect 131205 329291 131271 329294
rect 186313 328946 186379 328949
rect 186313 328944 190164 328946
rect 186313 328888 186318 328944
rect 186374 328888 190164 328944
rect 186313 328886 190164 328888
rect 186313 328883 186379 328886
rect 131297 328810 131363 328813
rect 129968 328808 131363 328810
rect 129968 328752 131302 328808
rect 131358 328752 131363 328808
rect 129968 328750 131363 328752
rect 131297 328747 131363 328750
rect 437473 328810 437539 328813
rect 437473 328808 440036 328810
rect 437473 328752 437478 328808
rect 437534 328752 440036 328808
rect 437473 328750 440036 328752
rect 437473 328747 437539 328750
rect 131113 328266 131179 328269
rect 129968 328264 131179 328266
rect 129968 328208 131118 328264
rect 131174 328208 131179 328264
rect 129968 328206 131179 328208
rect 131113 328203 131179 328206
rect 186313 327858 186379 327861
rect 186313 327856 190164 327858
rect 186313 327800 186318 327856
rect 186374 327800 190164 327856
rect 186313 327798 190164 327800
rect 186313 327795 186379 327798
rect 131205 327586 131271 327589
rect 129968 327584 131271 327586
rect 129968 327528 131210 327584
rect 131266 327528 131271 327584
rect 129968 327526 131271 327528
rect 131205 327523 131271 327526
rect 437473 327178 437539 327181
rect 437473 327176 440036 327178
rect 437473 327120 437478 327176
rect 437534 327120 440036 327176
rect 437473 327118 440036 327120
rect 437473 327115 437539 327118
rect 132217 327042 132283 327045
rect 129968 327040 132283 327042
rect 129968 326984 132222 327040
rect 132278 326984 132283 327040
rect 129968 326982 132283 326984
rect 132217 326979 132283 326982
rect 186313 326770 186379 326773
rect 186313 326768 190164 326770
rect 186313 326712 186318 326768
rect 186374 326712 190164 326768
rect 186313 326710 190164 326712
rect 186313 326707 186379 326710
rect 131297 326498 131363 326501
rect 411253 326498 411319 326501
rect 129968 326496 131363 326498
rect 129968 326440 131302 326496
rect 131358 326440 131363 326496
rect 129968 326438 131363 326440
rect 409860 326496 411319 326498
rect 409860 326440 411258 326496
rect 411314 326440 411319 326496
rect 409860 326438 411319 326440
rect 131297 326435 131363 326438
rect 411253 326435 411319 326438
rect 131205 325954 131271 325957
rect 129968 325952 131271 325954
rect 129968 325896 131210 325952
rect 131266 325896 131271 325952
rect 129968 325894 131271 325896
rect 131205 325891 131271 325894
rect 186405 325818 186471 325821
rect 186405 325816 190164 325818
rect 186405 325760 186410 325816
rect 186466 325760 190164 325816
rect 186405 325758 190164 325760
rect 186405 325755 186471 325758
rect 438761 325546 438827 325549
rect 438761 325544 440036 325546
rect 438761 325488 438766 325544
rect 438822 325488 440036 325544
rect 438761 325486 440036 325488
rect 438761 325483 438827 325486
rect 131205 325274 131271 325277
rect 129968 325272 131271 325274
rect 129968 325216 131210 325272
rect 131266 325216 131271 325272
rect 129968 325214 131271 325216
rect 131205 325211 131271 325214
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 131481 324730 131547 324733
rect 129968 324728 131547 324730
rect 129968 324672 131486 324728
rect 131542 324672 131547 324728
rect 129968 324670 131547 324672
rect 131481 324667 131547 324670
rect 186313 324730 186379 324733
rect 186313 324728 190164 324730
rect 186313 324672 186318 324728
rect 186374 324672 190164 324728
rect 186313 324670 190164 324672
rect 186313 324667 186379 324670
rect 411253 324458 411319 324461
rect 409860 324456 411319 324458
rect 409860 324400 411258 324456
rect 411314 324400 411319 324456
rect 409860 324398 411319 324400
rect 411253 324395 411319 324398
rect 131113 324186 131179 324189
rect 129968 324184 131179 324186
rect 129968 324128 131118 324184
rect 131174 324128 131179 324184
rect 129968 324126 131179 324128
rect 131113 324123 131179 324126
rect 438577 323914 438643 323917
rect 438577 323912 440036 323914
rect 438577 323856 438582 323912
rect 438638 323856 440036 323912
rect 438577 323854 440036 323856
rect 438577 323851 438643 323854
rect 186313 323642 186379 323645
rect 186313 323640 190164 323642
rect 186313 323584 186318 323640
rect 186374 323584 190164 323640
rect 186313 323582 190164 323584
rect 186313 323579 186379 323582
rect 131481 323506 131547 323509
rect 129968 323504 131547 323506
rect 129968 323448 131486 323504
rect 131542 323448 131547 323504
rect 129968 323446 131547 323448
rect 131481 323443 131547 323446
rect 131205 322962 131271 322965
rect 129968 322960 131271 322962
rect 129968 322904 131210 322960
rect 131266 322904 131271 322960
rect 129968 322902 131271 322904
rect 131205 322899 131271 322902
rect 186313 322690 186379 322693
rect 186313 322688 190164 322690
rect 186313 322632 186318 322688
rect 186374 322632 190164 322688
rect 186313 322630 190164 322632
rect 186313 322627 186379 322630
rect 131113 322418 131179 322421
rect 411529 322418 411595 322421
rect 129968 322416 131179 322418
rect 129968 322360 131118 322416
rect 131174 322360 131179 322416
rect 129968 322358 131179 322360
rect 409860 322416 411595 322418
rect 409860 322360 411534 322416
rect 411590 322360 411595 322416
rect 409860 322358 411595 322360
rect 131113 322355 131179 322358
rect 411529 322355 411595 322358
rect 438485 322146 438551 322149
rect 438485 322144 440036 322146
rect 438485 322088 438490 322144
rect 438546 322088 440036 322144
rect 438485 322086 440036 322088
rect 438485 322083 438551 322086
rect 131205 321874 131271 321877
rect 129968 321872 131271 321874
rect 129968 321816 131210 321872
rect 131266 321816 131271 321872
rect 129968 321814 131271 321816
rect 131205 321811 131271 321814
rect 186405 321602 186471 321605
rect 186405 321600 190164 321602
rect 186405 321544 186410 321600
rect 186466 321544 190164 321600
rect 186405 321542 190164 321544
rect 186405 321539 186471 321542
rect 131113 321194 131179 321197
rect 129968 321192 131179 321194
rect 129968 321136 131118 321192
rect 131174 321136 131179 321192
rect 129968 321134 131179 321136
rect 131113 321131 131179 321134
rect 409965 320922 410031 320925
rect 409830 320920 410031 320922
rect 409830 320864 409970 320920
rect 410026 320864 410031 320920
rect 409830 320862 410031 320864
rect 131205 320650 131271 320653
rect 129968 320648 131271 320650
rect 129968 320592 131210 320648
rect 131266 320592 131271 320648
rect 129968 320590 131271 320592
rect 131205 320587 131271 320590
rect 186313 320514 186379 320517
rect 186313 320512 190164 320514
rect 186313 320456 186318 320512
rect 186374 320456 190164 320512
rect 186313 320454 190164 320456
rect 186313 320451 186379 320454
rect 409830 320348 409890 320862
rect 409965 320859 410031 320862
rect 552105 320650 552171 320653
rect 549884 320648 552171 320650
rect 549884 320592 552110 320648
rect 552166 320592 552171 320648
rect 549884 320590 552171 320592
rect 552105 320587 552171 320590
rect 438393 320514 438459 320517
rect 438393 320512 440036 320514
rect 438393 320456 438398 320512
rect 438454 320456 440036 320512
rect 438393 320454 440036 320456
rect 438393 320451 438459 320454
rect 131941 320106 132007 320109
rect 129968 320104 132007 320106
rect 129968 320048 131946 320104
rect 132002 320048 132007 320104
rect 129968 320046 132007 320048
rect 131941 320043 132007 320046
rect 132217 319562 132283 319565
rect 129968 319560 132283 319562
rect 129968 319504 132222 319560
rect 132278 319504 132283 319560
rect 129968 319502 132283 319504
rect 132217 319499 132283 319502
rect 186313 319426 186379 319429
rect 186313 319424 190164 319426
rect -960 319140 480 319380
rect 186313 319368 186318 319424
rect 186374 319368 190164 319424
rect 186313 319366 190164 319368
rect 186313 319363 186379 319366
rect 131205 318882 131271 318885
rect 129968 318880 131271 318882
rect 129968 318824 131210 318880
rect 131266 318824 131271 318880
rect 129968 318822 131271 318824
rect 131205 318819 131271 318822
rect 437473 318882 437539 318885
rect 437473 318880 440036 318882
rect 437473 318824 437478 318880
rect 437534 318824 440036 318880
rect 437473 318822 440036 318824
rect 437473 318819 437539 318822
rect 186313 318474 186379 318477
rect 186313 318472 190164 318474
rect 186313 318416 186318 318472
rect 186374 318416 190164 318472
rect 186313 318414 190164 318416
rect 186313 318411 186379 318414
rect 132125 318338 132191 318341
rect 129968 318336 132191 318338
rect 129968 318280 132130 318336
rect 132186 318280 132191 318336
rect 129968 318278 132191 318280
rect 132125 318275 132191 318278
rect 411253 318202 411319 318205
rect 409860 318200 411319 318202
rect 409860 318144 411258 318200
rect 411314 318144 411319 318200
rect 409860 318142 411319 318144
rect 411253 318139 411319 318142
rect 131481 317794 131547 317797
rect 129968 317792 131547 317794
rect 129968 317736 131486 317792
rect 131542 317736 131547 317792
rect 129968 317734 131547 317736
rect 131481 317731 131547 317734
rect 186405 317386 186471 317389
rect 186405 317384 190164 317386
rect 186405 317328 186410 317384
rect 186466 317328 190164 317384
rect 186405 317326 190164 317328
rect 186405 317323 186471 317326
rect 438669 317250 438735 317253
rect 438669 317248 440036 317250
rect 438669 317192 438674 317248
rect 438730 317192 440036 317248
rect 438669 317190 440036 317192
rect 438669 317187 438735 317190
rect 132217 317114 132283 317117
rect 129968 317112 132283 317114
rect 129968 317056 132222 317112
rect 132278 317056 132283 317112
rect 129968 317054 132283 317056
rect 132217 317051 132283 317054
rect 131205 316570 131271 316573
rect 129968 316568 131271 316570
rect 129968 316512 131210 316568
rect 131266 316512 131271 316568
rect 129968 316510 131271 316512
rect 131205 316507 131271 316510
rect 186313 316298 186379 316301
rect 186313 316296 190164 316298
rect 186313 316240 186318 316296
rect 186374 316240 190164 316296
rect 186313 316238 190164 316240
rect 186313 316235 186379 316238
rect 411253 316162 411319 316165
rect 409860 316160 411319 316162
rect 409860 316104 411258 316160
rect 411314 316104 411319 316160
rect 409860 316102 411319 316104
rect 411253 316099 411319 316102
rect 131481 316026 131547 316029
rect 129968 316024 131547 316026
rect 129968 315968 131486 316024
rect 131542 315968 131547 316024
rect 129968 315966 131547 315968
rect 131481 315963 131547 315966
rect 437473 315618 437539 315621
rect 437473 315616 440036 315618
rect 437473 315560 437478 315616
rect 437534 315560 440036 315616
rect 437473 315558 440036 315560
rect 437473 315555 437539 315558
rect 131205 315482 131271 315485
rect 129968 315480 131271 315482
rect 129968 315424 131210 315480
rect 131266 315424 131271 315480
rect 129968 315422 131271 315424
rect 131205 315419 131271 315422
rect 186313 315210 186379 315213
rect 186313 315208 190164 315210
rect 186313 315152 186318 315208
rect 186374 315152 190164 315208
rect 186313 315150 190164 315152
rect 186313 315147 186379 315150
rect 131297 314802 131363 314805
rect 129968 314800 131363 314802
rect 129968 314744 131302 314800
rect 131358 314744 131363 314800
rect 129968 314742 131363 314744
rect 131297 314739 131363 314742
rect 131113 314258 131179 314261
rect 129968 314256 131179 314258
rect 129968 314200 131118 314256
rect 131174 314200 131179 314256
rect 129968 314198 131179 314200
rect 131113 314195 131179 314198
rect 186313 314258 186379 314261
rect 186313 314256 190164 314258
rect 186313 314200 186318 314256
rect 186374 314200 190164 314256
rect 186313 314198 190164 314200
rect 186313 314195 186379 314198
rect 411253 314122 411319 314125
rect 409860 314120 411319 314122
rect 409860 314064 411258 314120
rect 411314 314064 411319 314120
rect 409860 314062 411319 314064
rect 411253 314059 411319 314062
rect 437473 313986 437539 313989
rect 437473 313984 440036 313986
rect 437473 313928 437478 313984
rect 437534 313928 440036 313984
rect 437473 313926 440036 313928
rect 437473 313923 437539 313926
rect 131205 313714 131271 313717
rect 129968 313712 131271 313714
rect 129968 313656 131210 313712
rect 131266 313656 131271 313712
rect 129968 313654 131271 313656
rect 131205 313651 131271 313654
rect 131297 313170 131363 313173
rect 129968 313168 131363 313170
rect 129968 313112 131302 313168
rect 131358 313112 131363 313168
rect 129968 313110 131363 313112
rect 131297 313107 131363 313110
rect 186313 313170 186379 313173
rect 186313 313168 190164 313170
rect 186313 313112 186318 313168
rect 186374 313112 190164 313168
rect 186313 313110 190164 313112
rect 186313 313107 186379 313110
rect 131113 312490 131179 312493
rect 129968 312488 131179 312490
rect 129968 312432 131118 312488
rect 131174 312432 131179 312488
rect 129968 312430 131179 312432
rect 131113 312427 131179 312430
rect 438025 312354 438091 312357
rect 438025 312352 440036 312354
rect 438025 312296 438030 312352
rect 438086 312296 440036 312352
rect 438025 312294 440036 312296
rect 438025 312291 438091 312294
rect 186405 312082 186471 312085
rect 411253 312082 411319 312085
rect 186405 312080 190164 312082
rect 186405 312024 186410 312080
rect 186466 312024 190164 312080
rect 186405 312022 190164 312024
rect 409860 312080 411319 312082
rect 409860 312024 411258 312080
rect 411314 312024 411319 312080
rect 409860 312022 411319 312024
rect 186405 312019 186471 312022
rect 411253 312019 411319 312022
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 131205 311946 131271 311949
rect 129968 311944 131271 311946
rect 129968 311888 131210 311944
rect 131266 311888 131271 311944
rect 583520 311932 584960 312022
rect 129968 311886 131271 311888
rect 131205 311883 131271 311886
rect 131205 311402 131271 311405
rect 129968 311400 131271 311402
rect 129968 311344 131210 311400
rect 131266 311344 131271 311400
rect 129968 311342 131271 311344
rect 131205 311339 131271 311342
rect 186313 310994 186379 310997
rect 186313 310992 190164 310994
rect 186313 310936 186318 310992
rect 186374 310936 190164 310992
rect 186313 310934 190164 310936
rect 186313 310931 186379 310934
rect 131481 310722 131547 310725
rect 129968 310720 131547 310722
rect 129968 310664 131486 310720
rect 131542 310664 131547 310720
rect 129968 310662 131547 310664
rect 131481 310659 131547 310662
rect 437473 310722 437539 310725
rect 437473 310720 440036 310722
rect 437473 310664 437478 310720
rect 437534 310664 440036 310720
rect 437473 310662 440036 310664
rect 437473 310659 437539 310662
rect 131113 310178 131179 310181
rect 129968 310176 131179 310178
rect 129968 310120 131118 310176
rect 131174 310120 131179 310176
rect 129968 310118 131179 310120
rect 131113 310115 131179 310118
rect 186313 310042 186379 310045
rect 411253 310042 411319 310045
rect 186313 310040 190164 310042
rect 186313 309984 186318 310040
rect 186374 309984 190164 310040
rect 186313 309982 190164 309984
rect 409860 310040 411319 310042
rect 409860 309984 411258 310040
rect 411314 309984 411319 310040
rect 409860 309982 411319 309984
rect 186313 309979 186379 309982
rect 411253 309979 411319 309982
rect 131205 309634 131271 309637
rect 129968 309632 131271 309634
rect 129968 309576 131210 309632
rect 131266 309576 131271 309632
rect 129968 309574 131271 309576
rect 131205 309571 131271 309574
rect 131113 309090 131179 309093
rect 129968 309088 131179 309090
rect 129968 309032 131118 309088
rect 131174 309032 131179 309088
rect 129968 309030 131179 309032
rect 131113 309027 131179 309030
rect 437473 309090 437539 309093
rect 437473 309088 440036 309090
rect 437473 309032 437478 309088
rect 437534 309032 440036 309088
rect 437473 309030 440036 309032
rect 437473 309027 437539 309030
rect 186313 308954 186379 308957
rect 186313 308952 190164 308954
rect 186313 308896 186318 308952
rect 186374 308896 190164 308952
rect 186313 308894 190164 308896
rect 186313 308891 186379 308894
rect 131481 308410 131547 308413
rect 129968 308408 131547 308410
rect 129968 308352 131486 308408
rect 131542 308352 131547 308408
rect 129968 308350 131547 308352
rect 131481 308347 131547 308350
rect 410517 308002 410583 308005
rect 409860 308000 410583 308002
rect 409860 307972 410522 308000
rect 409830 307944 410522 307972
rect 410578 307944 410583 308000
rect 409830 307942 410583 307944
rect 131205 307866 131271 307869
rect 129968 307864 131271 307866
rect 129968 307808 131210 307864
rect 131266 307808 131271 307864
rect 129968 307806 131271 307808
rect 131205 307803 131271 307806
rect 186405 307866 186471 307869
rect 186405 307864 190164 307866
rect 186405 307808 186410 307864
rect 186466 307808 190164 307864
rect 186405 307806 190164 307808
rect 186405 307803 186471 307806
rect 409830 307733 409890 307942
rect 410517 307939 410583 307942
rect 409830 307728 409939 307733
rect 409830 307672 409878 307728
rect 409934 307672 409939 307728
rect 409830 307670 409939 307672
rect 409873 307667 409939 307670
rect 437565 307458 437631 307461
rect 437565 307456 440036 307458
rect 437565 307400 437570 307456
rect 437626 307400 440036 307456
rect 437565 307398 440036 307400
rect 437565 307395 437631 307398
rect 131113 307322 131179 307325
rect 129968 307320 131179 307322
rect 129968 307264 131118 307320
rect 131174 307264 131179 307320
rect 129968 307262 131179 307264
rect 131113 307259 131179 307262
rect 131205 306778 131271 306781
rect 129968 306776 131271 306778
rect 129968 306720 131210 306776
rect 131266 306720 131271 306776
rect 129968 306718 131271 306720
rect 131205 306715 131271 306718
rect 186313 306778 186379 306781
rect 186313 306776 190164 306778
rect 186313 306720 186318 306776
rect 186374 306720 190164 306776
rect 186313 306718 190164 306720
rect 186313 306715 186379 306718
rect 549854 306506 549914 306884
rect 550541 306506 550607 306509
rect 549854 306504 550607 306506
rect 549854 306448 550546 306504
rect 550602 306448 550607 306504
rect 549854 306446 550607 306448
rect 550541 306443 550607 306446
rect -960 306084 480 306324
rect 131113 306098 131179 306101
rect 129968 306096 131179 306098
rect 129968 306040 131118 306096
rect 131174 306040 131179 306096
rect 129968 306038 131179 306040
rect 131113 306035 131179 306038
rect 186313 305826 186379 305829
rect 186313 305824 190164 305826
rect 186313 305768 186318 305824
rect 186374 305768 190164 305824
rect 186313 305766 190164 305768
rect 186313 305763 186379 305766
rect 131481 305554 131547 305557
rect 129968 305552 131547 305554
rect 129968 305496 131486 305552
rect 131542 305496 131547 305552
rect 129968 305494 131547 305496
rect 131481 305491 131547 305494
rect 409830 305418 409890 305932
rect 437473 305826 437539 305829
rect 437473 305824 440036 305826
rect 437473 305768 437478 305824
rect 437534 305768 440036 305824
rect 437473 305766 440036 305768
rect 437473 305763 437539 305766
rect 409965 305418 410031 305421
rect 409830 305416 410031 305418
rect 409830 305360 409970 305416
rect 410026 305360 410031 305416
rect 409830 305358 410031 305360
rect 409965 305355 410031 305358
rect 131205 305010 131271 305013
rect 129968 305008 131271 305010
rect 129968 304952 131210 305008
rect 131266 304952 131271 305008
rect 129968 304950 131271 304952
rect 131205 304947 131271 304950
rect 186681 304738 186747 304741
rect 186681 304736 190164 304738
rect 186681 304680 186686 304736
rect 186742 304680 190164 304736
rect 186681 304678 190164 304680
rect 186681 304675 186747 304678
rect 131297 304330 131363 304333
rect 129968 304328 131363 304330
rect 129968 304272 131302 304328
rect 131358 304272 131363 304328
rect 129968 304270 131363 304272
rect 131297 304267 131363 304270
rect 436829 304194 436895 304197
rect 436829 304192 440036 304194
rect 436829 304136 436834 304192
rect 436890 304136 440036 304192
rect 436829 304134 440036 304136
rect 436829 304131 436895 304134
rect 411253 303922 411319 303925
rect 409860 303920 411319 303922
rect 409860 303864 411258 303920
rect 411314 303864 411319 303920
rect 409860 303862 411319 303864
rect 411253 303859 411319 303862
rect 131205 303786 131271 303789
rect 129968 303784 131271 303786
rect 129968 303728 131210 303784
rect 131266 303728 131271 303784
rect 129968 303726 131271 303728
rect 131205 303723 131271 303726
rect 186405 303650 186471 303653
rect 186405 303648 190164 303650
rect 186405 303592 186410 303648
rect 186466 303592 190164 303648
rect 186405 303590 190164 303592
rect 186405 303587 186471 303590
rect 131113 303242 131179 303245
rect 129968 303240 131179 303242
rect 129968 303184 131118 303240
rect 131174 303184 131179 303240
rect 129968 303182 131179 303184
rect 131113 303179 131179 303182
rect 131205 302698 131271 302701
rect 129968 302696 131271 302698
rect 129968 302640 131210 302696
rect 131266 302640 131271 302696
rect 129968 302638 131271 302640
rect 131205 302635 131271 302638
rect 186313 302562 186379 302565
rect 438301 302562 438367 302565
rect 186313 302560 190164 302562
rect 186313 302504 186318 302560
rect 186374 302504 190164 302560
rect 186313 302502 190164 302504
rect 438301 302560 440036 302562
rect 438301 302504 438306 302560
rect 438362 302504 440036 302560
rect 438301 302502 440036 302504
rect 186313 302499 186379 302502
rect 438301 302499 438367 302502
rect 131481 302018 131547 302021
rect 129968 302016 131547 302018
rect 129968 301960 131486 302016
rect 131542 301960 131547 302016
rect 129968 301958 131547 301960
rect 131481 301955 131547 301958
rect 411294 301746 411300 301748
rect 409860 301686 411300 301746
rect 411294 301684 411300 301686
rect 411364 301746 411370 301748
rect 411529 301746 411595 301749
rect 411364 301744 411595 301746
rect 411364 301688 411534 301744
rect 411590 301688 411595 301744
rect 411364 301686 411595 301688
rect 411364 301684 411370 301686
rect 411529 301683 411595 301686
rect 186313 301610 186379 301613
rect 186313 301608 190164 301610
rect 186313 301552 186318 301608
rect 186374 301552 190164 301608
rect 186313 301550 190164 301552
rect 186313 301547 186379 301550
rect 132033 301474 132099 301477
rect 129968 301472 132099 301474
rect 129968 301416 132038 301472
rect 132094 301416 132099 301472
rect 129968 301414 132099 301416
rect 132033 301411 132099 301414
rect 131205 300930 131271 300933
rect 129968 300928 131271 300930
rect 129968 300872 131210 300928
rect 131266 300872 131271 300928
rect 129968 300870 131271 300872
rect 131205 300867 131271 300870
rect 438393 300930 438459 300933
rect 438393 300928 440036 300930
rect 438393 300872 438398 300928
rect 438454 300872 440036 300928
rect 438393 300870 440036 300872
rect 438393 300867 438459 300870
rect 186313 300522 186379 300525
rect 186313 300520 190164 300522
rect 186313 300464 186318 300520
rect 186374 300464 190164 300520
rect 186313 300462 190164 300464
rect 186313 300459 186379 300462
rect 129782 300114 129842 300356
rect 131113 300114 131179 300117
rect 129782 300112 131179 300114
rect 129782 300056 131118 300112
rect 131174 300056 131179 300112
rect 129782 300054 131179 300056
rect 131113 300051 131179 300054
rect 410149 299706 410215 299709
rect 410517 299706 410583 299709
rect 409860 299704 410583 299706
rect 409860 299648 410154 299704
rect 410210 299648 410522 299704
rect 410578 299648 410583 299704
rect 409860 299646 410583 299648
rect 410149 299643 410215 299646
rect 410517 299643 410583 299646
rect 186313 299434 186379 299437
rect 186313 299432 190164 299434
rect 186313 299376 186318 299432
rect 186374 299376 190164 299432
rect 186313 299374 190164 299376
rect 186313 299371 186379 299374
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 186405 298346 186471 298349
rect 186405 298344 190164 298346
rect 186405 298288 186410 298344
rect 186466 298288 190164 298344
rect 186405 298286 190164 298288
rect 186405 298283 186471 298286
rect 411253 297666 411319 297669
rect 411478 297666 411484 297668
rect 409860 297664 411484 297666
rect 409860 297608 411258 297664
rect 411314 297608 411484 297664
rect 409860 297606 411484 297608
rect 411253 297603 411319 297606
rect 411478 297604 411484 297606
rect 411548 297604 411554 297668
rect 186313 297394 186379 297397
rect 186313 297392 190164 297394
rect 186313 297336 186318 297392
rect 186374 297336 190164 297392
rect 186313 297334 190164 297336
rect 186313 297331 186379 297334
rect 186313 296306 186379 296309
rect 186313 296304 190164 296306
rect 186313 296248 186318 296304
rect 186374 296248 190164 296304
rect 186313 296246 190164 296248
rect 186313 296243 186379 296246
rect 410149 295626 410215 295629
rect 409860 295624 410215 295626
rect 409860 295568 410154 295624
rect 410210 295568 410215 295624
rect 409860 295566 410215 295568
rect 410149 295563 410215 295566
rect 186313 295218 186379 295221
rect 186313 295216 190164 295218
rect 186313 295160 186318 295216
rect 186374 295160 190164 295216
rect 186313 295158 190164 295160
rect 186313 295155 186379 295158
rect 186405 294266 186471 294269
rect 186405 294264 190164 294266
rect 186405 294208 186410 294264
rect 186466 294208 190164 294264
rect 186405 294206 190164 294208
rect 186405 294203 186471 294206
rect 411253 293586 411319 293589
rect 409860 293584 411319 293586
rect 409860 293528 411258 293584
rect 411314 293528 411319 293584
rect 409860 293526 411319 293528
rect 411253 293523 411319 293526
rect -960 293028 480 293268
rect 186313 293178 186379 293181
rect 186313 293176 190164 293178
rect 186313 293120 186318 293176
rect 186374 293120 190164 293176
rect 186313 293118 190164 293120
rect 186313 293115 186379 293118
rect 186313 292090 186379 292093
rect 186313 292088 190164 292090
rect 186313 292032 186318 292088
rect 186374 292032 190164 292088
rect 186313 292030 190164 292032
rect 186313 292027 186379 292030
rect 411253 291546 411319 291549
rect 409860 291544 411319 291546
rect 409860 291488 411258 291544
rect 411314 291488 411319 291544
rect 409860 291486 411319 291488
rect 411253 291483 411319 291486
rect 186313 291002 186379 291005
rect 186313 291000 190164 291002
rect 186313 290944 186318 291000
rect 186374 290944 190164 291000
rect 186313 290942 190164 290944
rect 186313 290939 186379 290942
rect 186405 290050 186471 290053
rect 186405 290048 190164 290050
rect 186405 289992 186410 290048
rect 186466 289992 190164 290048
rect 186405 289990 190164 289992
rect 186405 289987 186471 289990
rect 411253 289506 411319 289509
rect 409860 289504 411319 289506
rect 409860 289448 411258 289504
rect 411314 289448 411319 289504
rect 409860 289446 411319 289448
rect 411253 289443 411319 289446
rect 186313 288962 186379 288965
rect 186313 288960 190164 288962
rect 186313 288904 186318 288960
rect 186374 288904 190164 288960
rect 186313 288902 190164 288904
rect 186313 288899 186379 288902
rect 186313 287874 186379 287877
rect 186313 287872 190164 287874
rect 186313 287816 186318 287872
rect 186374 287816 190164 287872
rect 186313 287814 190164 287816
rect 186313 287811 186379 287814
rect 411253 287466 411319 287469
rect 409860 287464 411319 287466
rect 409860 287408 411258 287464
rect 411314 287408 411319 287464
rect 409860 287406 411319 287408
rect 411253 287403 411319 287406
rect 186313 286786 186379 286789
rect 186313 286784 190164 286786
rect 186313 286728 186318 286784
rect 186374 286728 190164 286784
rect 186313 286726 190164 286728
rect 186313 286723 186379 286726
rect 186405 285834 186471 285837
rect 186405 285832 190164 285834
rect 186405 285776 186410 285832
rect 186466 285776 190164 285832
rect 186405 285774 190164 285776
rect 186405 285771 186471 285774
rect 411253 285290 411319 285293
rect 409860 285288 411319 285290
rect 409860 285232 411258 285288
rect 411314 285232 411319 285288
rect 583520 285276 584960 285516
rect 409860 285230 411319 285232
rect 411253 285227 411319 285230
rect 186313 284746 186379 284749
rect 186313 284744 190164 284746
rect 186313 284688 186318 284744
rect 186374 284688 190164 284744
rect 186313 284686 190164 284688
rect 186313 284683 186379 284686
rect 186313 283658 186379 283661
rect 186313 283656 190164 283658
rect 186313 283600 186318 283656
rect 186374 283600 190164 283656
rect 186313 283598 190164 283600
rect 186313 283595 186379 283598
rect 411253 283250 411319 283253
rect 409860 283248 411319 283250
rect 409860 283192 411258 283248
rect 411314 283192 411319 283248
rect 409860 283190 411319 283192
rect 411253 283187 411319 283190
rect 186313 282570 186379 282573
rect 186313 282568 190164 282570
rect 186313 282512 186318 282568
rect 186374 282512 190164 282568
rect 186313 282510 190164 282512
rect 186313 282507 186379 282510
rect 186405 281618 186471 281621
rect 186405 281616 190164 281618
rect 186405 281560 186410 281616
rect 186466 281560 190164 281616
rect 186405 281558 190164 281560
rect 186405 281555 186471 281558
rect 411253 281210 411319 281213
rect 409860 281208 411319 281210
rect 409860 281152 411258 281208
rect 411314 281152 411319 281208
rect 409860 281150 411319 281152
rect 411253 281147 411319 281150
rect 186313 280530 186379 280533
rect 186313 280528 190164 280530
rect 186313 280472 186318 280528
rect 186374 280472 190164 280528
rect 186313 280470 190164 280472
rect 186313 280467 186379 280470
rect -960 279972 480 280212
rect 186313 279442 186379 279445
rect 186313 279440 190164 279442
rect 186313 279384 186318 279440
rect 186374 279384 190164 279440
rect 186313 279382 190164 279384
rect 186313 279379 186379 279382
rect 411253 279170 411319 279173
rect 409860 279168 411319 279170
rect 409860 279112 411258 279168
rect 411314 279112 411319 279168
rect 409860 279110 411319 279112
rect 411253 279107 411319 279110
rect 186313 278354 186379 278357
rect 186313 278352 190164 278354
rect 186313 278296 186318 278352
rect 186374 278296 190164 278352
rect 186313 278294 190164 278296
rect 186313 278291 186379 278294
rect 186313 277402 186379 277405
rect 186313 277400 190164 277402
rect 186313 277344 186318 277400
rect 186374 277344 190164 277400
rect 186313 277342 190164 277344
rect 186313 277339 186379 277342
rect 411253 277130 411319 277133
rect 409860 277128 411319 277130
rect 409860 277072 411258 277128
rect 411314 277072 411319 277128
rect 409860 277070 411319 277072
rect 411253 277067 411319 277070
rect 186405 276314 186471 276317
rect 186405 276312 190164 276314
rect 186405 276256 186410 276312
rect 186466 276256 190164 276312
rect 186405 276254 190164 276256
rect 186405 276251 186471 276254
rect 186313 275226 186379 275229
rect 186313 275224 190164 275226
rect 186313 275168 186318 275224
rect 186374 275168 190164 275224
rect 186313 275166 190164 275168
rect 186313 275163 186379 275166
rect 411253 275090 411319 275093
rect 409860 275088 411319 275090
rect 409860 275032 411258 275088
rect 411314 275032 411319 275088
rect 409860 275030 411319 275032
rect 411253 275027 411319 275030
rect 186313 274138 186379 274141
rect 186313 274136 190164 274138
rect 186313 274080 186318 274136
rect 186374 274080 190164 274136
rect 186313 274078 190164 274080
rect 186313 274075 186379 274078
rect 186313 273186 186379 273189
rect 186313 273184 190164 273186
rect 186313 273128 186318 273184
rect 186374 273128 190164 273184
rect 186313 273126 190164 273128
rect 186313 273123 186379 273126
rect 411253 273050 411319 273053
rect 409860 273048 411319 273050
rect 409860 272992 411258 273048
rect 411314 272992 411319 273048
rect 409860 272990 411319 272992
rect 411253 272987 411319 272990
rect 579797 272234 579863 272237
rect 583520 272234 584960 272324
rect 579797 272232 584960 272234
rect 579797 272176 579802 272232
rect 579858 272176 584960 272232
rect 579797 272174 584960 272176
rect 579797 272171 579863 272174
rect 186405 272098 186471 272101
rect 186405 272096 190164 272098
rect 186405 272040 186410 272096
rect 186466 272040 190164 272096
rect 583520 272084 584960 272174
rect 186405 272038 190164 272040
rect 186405 272035 186471 272038
rect 186313 271010 186379 271013
rect 411253 271010 411319 271013
rect 186313 271008 190164 271010
rect 186313 270952 186318 271008
rect 186374 270952 190164 271008
rect 186313 270950 190164 270952
rect 409860 271008 411319 271010
rect 409860 270952 411258 271008
rect 411314 270952 411319 271008
rect 409860 270950 411319 270952
rect 186313 270947 186379 270950
rect 411253 270947 411319 270950
rect 186313 269922 186379 269925
rect 186313 269920 190164 269922
rect 186313 269864 186318 269920
rect 186374 269864 190164 269920
rect 186313 269862 190164 269864
rect 186313 269859 186379 269862
rect 186405 268970 186471 268973
rect 411253 268970 411319 268973
rect 186405 268968 190164 268970
rect 186405 268912 186410 268968
rect 186466 268912 190164 268968
rect 186405 268910 190164 268912
rect 409860 268968 411319 268970
rect 409860 268912 411258 268968
rect 411314 268912 411319 268968
rect 409860 268910 411319 268912
rect 186405 268907 186471 268910
rect 411253 268907 411319 268910
rect 186313 267882 186379 267885
rect 186313 267880 190164 267882
rect 186313 267824 186318 267880
rect 186374 267824 190164 267880
rect 186313 267822 190164 267824
rect 186313 267819 186379 267822
rect -960 267052 480 267292
rect 186313 266794 186379 266797
rect 411253 266794 411319 266797
rect 186313 266792 190164 266794
rect 186313 266736 186318 266792
rect 186374 266736 190164 266792
rect 186313 266734 190164 266736
rect 409860 266792 411319 266794
rect 409860 266736 411258 266792
rect 411314 266736 411319 266792
rect 409860 266734 411319 266736
rect 186313 266731 186379 266734
rect 411253 266731 411319 266734
rect 186313 265706 186379 265709
rect 186313 265704 190164 265706
rect 186313 265648 186318 265704
rect 186374 265648 190164 265704
rect 186313 265646 190164 265648
rect 186313 265643 186379 265646
rect 186313 264754 186379 264757
rect 411253 264754 411319 264757
rect 186313 264752 190164 264754
rect 186313 264696 186318 264752
rect 186374 264696 190164 264752
rect 186313 264694 190164 264696
rect 409860 264752 411319 264754
rect 409860 264696 411258 264752
rect 411314 264696 411319 264752
rect 409860 264694 411319 264696
rect 186313 264691 186379 264694
rect 411253 264691 411319 264694
rect 186405 263666 186471 263669
rect 186405 263664 190164 263666
rect 186405 263608 186410 263664
rect 186466 263608 190164 263664
rect 186405 263606 190164 263608
rect 186405 263603 186471 263606
rect 411253 262714 411319 262717
rect 409860 262712 411319 262714
rect 409860 262656 411258 262712
rect 411314 262656 411319 262712
rect 409860 262654 411319 262656
rect 411253 262651 411319 262654
rect 186313 262578 186379 262581
rect 186313 262576 190164 262578
rect 186313 262520 186318 262576
rect 186374 262520 190164 262576
rect 186313 262518 190164 262520
rect 186313 262515 186379 262518
rect 186313 261626 186379 261629
rect 186313 261624 190164 261626
rect 186313 261568 186318 261624
rect 186374 261568 190164 261624
rect 186313 261566 190164 261568
rect 186313 261563 186379 261566
rect 411253 260674 411319 260677
rect 409860 260672 411319 260674
rect 409860 260616 411258 260672
rect 411314 260616 411319 260672
rect 409860 260614 411319 260616
rect 411253 260611 411319 260614
rect 186313 260538 186379 260541
rect 186313 260536 190164 260538
rect 186313 260480 186318 260536
rect 186374 260480 190164 260536
rect 186313 260478 190164 260480
rect 186313 260475 186379 260478
rect 186405 259450 186471 259453
rect 186405 259448 190164 259450
rect 186405 259392 186410 259448
rect 186466 259392 190164 259448
rect 186405 259390 190164 259392
rect 186405 259387 186471 259390
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect 411253 258634 411319 258637
rect 409860 258632 411319 258634
rect 409860 258576 411258 258632
rect 411314 258576 411319 258632
rect 409860 258574 411319 258576
rect 411253 258571 411319 258574
rect 186313 258362 186379 258365
rect 186313 258360 190164 258362
rect 186313 258304 186318 258360
rect 186374 258304 190164 258360
rect 186313 258302 190164 258304
rect 186313 258299 186379 258302
rect 186313 257410 186379 257413
rect 186313 257408 190164 257410
rect 186313 257352 186318 257408
rect 186374 257352 190164 257408
rect 186313 257350 190164 257352
rect 186313 257347 186379 257350
rect 411253 256594 411319 256597
rect 409860 256592 411319 256594
rect 409860 256536 411258 256592
rect 411314 256536 411319 256592
rect 409860 256534 411319 256536
rect 411253 256531 411319 256534
rect 186313 256322 186379 256325
rect 186313 256320 190164 256322
rect 186313 256264 186318 256320
rect 186374 256264 190164 256320
rect 186313 256262 190164 256264
rect 186313 256259 186379 256262
rect 186313 255234 186379 255237
rect 186313 255232 190164 255234
rect 186313 255176 186318 255232
rect 186374 255176 190164 255232
rect 186313 255174 190164 255176
rect 186313 255171 186379 255174
rect 411253 254554 411319 254557
rect 409860 254552 411319 254554
rect 409860 254496 411258 254552
rect 411314 254496 411319 254552
rect 409860 254494 411319 254496
rect 411253 254491 411319 254494
rect -960 253996 480 254236
rect 186405 254146 186471 254149
rect 186405 254144 190164 254146
rect 186405 254088 186410 254144
rect 186466 254088 190164 254144
rect 186405 254086 190164 254088
rect 186405 254083 186471 254086
rect 186313 253194 186379 253197
rect 186313 253192 190164 253194
rect 186313 253136 186318 253192
rect 186374 253136 190164 253192
rect 186313 253134 190164 253136
rect 186313 253131 186379 253134
rect 410241 252514 410307 252517
rect 410793 252514 410859 252517
rect 409860 252512 410859 252514
rect 409860 252456 410246 252512
rect 410302 252456 410798 252512
rect 410854 252456 410859 252512
rect 409860 252454 410859 252456
rect 410241 252451 410307 252454
rect 410793 252451 410859 252454
rect 186313 252106 186379 252109
rect 186313 252104 190164 252106
rect 186313 252048 186318 252104
rect 186374 252048 190164 252104
rect 186313 252046 190164 252048
rect 186313 252043 186379 252046
rect 186313 251018 186379 251021
rect 186313 251016 190164 251018
rect 186313 250960 186318 251016
rect 186374 250960 190164 251016
rect 186313 250958 190164 250960
rect 186313 250955 186379 250958
rect 411253 250338 411319 250341
rect 409860 250336 411319 250338
rect 409860 250280 411258 250336
rect 411314 250280 411319 250336
rect 409860 250278 411319 250280
rect 411253 250275 411319 250278
rect 186405 249930 186471 249933
rect 186405 249928 190164 249930
rect 186405 249872 186410 249928
rect 186466 249872 190164 249928
rect 186405 249870 190164 249872
rect 186405 249867 186471 249870
rect 186313 248978 186379 248981
rect 186313 248976 190164 248978
rect 186313 248920 186318 248976
rect 186374 248920 190164 248976
rect 186313 248918 190164 248920
rect 186313 248915 186379 248918
rect 411805 248298 411871 248301
rect 409860 248296 411871 248298
rect 409860 248240 411810 248296
rect 411866 248240 411871 248296
rect 409860 248238 411871 248240
rect 411805 248235 411871 248238
rect 186313 247890 186379 247893
rect 186313 247888 190164 247890
rect 186313 247832 186318 247888
rect 186374 247832 190164 247888
rect 186313 247830 190164 247832
rect 186313 247827 186379 247830
rect 186313 246802 186379 246805
rect 186313 246800 190164 246802
rect 186313 246744 186318 246800
rect 186374 246744 190164 246800
rect 186313 246742 190164 246744
rect 186313 246739 186379 246742
rect 411253 246258 411319 246261
rect 409860 246256 411319 246258
rect 409860 246200 411258 246256
rect 411314 246200 411319 246256
rect 409860 246198 411319 246200
rect 411253 246195 411319 246198
rect 186405 245714 186471 245717
rect 186405 245712 190164 245714
rect 186405 245656 186410 245712
rect 186466 245656 190164 245712
rect 186405 245654 190164 245656
rect 186405 245651 186471 245654
rect 579797 245578 579863 245581
rect 583520 245578 584960 245668
rect 579797 245576 584960 245578
rect 579797 245520 579802 245576
rect 579858 245520 584960 245576
rect 579797 245518 584960 245520
rect 579797 245515 579863 245518
rect 583520 245428 584960 245518
rect 186313 244762 186379 244765
rect 186313 244760 190164 244762
rect 186313 244704 186318 244760
rect 186374 244704 190164 244760
rect 186313 244702 190164 244704
rect 186313 244699 186379 244702
rect 410517 244218 410583 244221
rect 410793 244218 410859 244221
rect 409860 244216 410859 244218
rect 409860 244160 410522 244216
rect 410578 244160 410798 244216
rect 410854 244160 410859 244216
rect 409860 244158 410859 244160
rect 410517 244155 410583 244158
rect 410793 244155 410859 244158
rect 186313 243674 186379 243677
rect 186313 243672 190164 243674
rect 186313 243616 186318 243672
rect 186374 243616 190164 243672
rect 186313 243614 190164 243616
rect 186313 243611 186379 243614
rect 186313 242586 186379 242589
rect 186313 242584 190164 242586
rect 186313 242528 186318 242584
rect 186374 242528 190164 242584
rect 186313 242526 190164 242528
rect 186313 242523 186379 242526
rect 411253 242178 411319 242181
rect 409860 242176 411319 242178
rect 409860 242120 411258 242176
rect 411314 242120 411319 242176
rect 409860 242118 411319 242120
rect 411253 242115 411319 242118
rect 186313 241498 186379 241501
rect 186313 241496 190164 241498
rect 186313 241440 186318 241496
rect 186374 241440 190164 241496
rect 186313 241438 190164 241440
rect 186313 241435 186379 241438
rect -960 240940 480 241180
rect 186405 240546 186471 240549
rect 186405 240544 190164 240546
rect 186405 240488 186410 240544
rect 186466 240488 190164 240544
rect 186405 240486 190164 240488
rect 186405 240483 186471 240486
rect 411253 240138 411319 240141
rect 411662 240138 411668 240140
rect 409860 240136 411668 240138
rect 409860 240080 411258 240136
rect 411314 240080 411668 240136
rect 409860 240078 411668 240080
rect 411253 240075 411319 240078
rect 411662 240076 411668 240078
rect 411732 240076 411738 240140
rect 186313 239458 186379 239461
rect 186313 239456 190164 239458
rect 186313 239400 186318 239456
rect 186374 239400 190164 239456
rect 186313 239398 190164 239400
rect 186313 239395 186379 239398
rect 186313 238370 186379 238373
rect 186313 238368 190164 238370
rect 186313 238312 186318 238368
rect 186374 238312 190164 238368
rect 186313 238310 190164 238312
rect 186313 238307 186379 238310
rect 411253 238098 411319 238101
rect 409860 238096 411319 238098
rect 409860 238040 411258 238096
rect 411314 238040 411319 238096
rect 409860 238038 411319 238040
rect 411253 238035 411319 238038
rect 186313 237282 186379 237285
rect 186313 237280 190164 237282
rect 186313 237224 186318 237280
rect 186374 237224 190164 237280
rect 186313 237222 190164 237224
rect 186313 237219 186379 237222
rect 186405 236330 186471 236333
rect 186405 236328 190164 236330
rect 186405 236272 186410 236328
rect 186466 236272 190164 236328
rect 186405 236270 190164 236272
rect 186405 236267 186471 236270
rect 409413 236194 409479 236197
rect 409413 236192 409522 236194
rect 409413 236136 409418 236192
rect 409474 236136 409522 236192
rect 409413 236131 409522 236136
rect 409462 236028 409522 236131
rect 186313 235242 186379 235245
rect 186313 235240 190164 235242
rect 186313 235184 186318 235240
rect 186374 235184 190164 235240
rect 186313 235182 190164 235184
rect 186313 235179 186379 235182
rect 186313 234154 186379 234157
rect 186313 234152 190164 234154
rect 186313 234096 186318 234152
rect 186374 234096 190164 234152
rect 186313 234094 190164 234096
rect 186313 234091 186379 234094
rect 411253 233882 411319 233885
rect 409860 233880 411319 233882
rect 409860 233824 411258 233880
rect 411314 233824 411319 233880
rect 409860 233822 411319 233824
rect 411253 233819 411319 233822
rect 186313 233066 186379 233069
rect 186313 233064 190164 233066
rect 186313 233008 186318 233064
rect 186374 233008 190164 233064
rect 186313 233006 190164 233008
rect 186313 233003 186379 233006
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect 186405 232114 186471 232117
rect 186405 232112 190164 232114
rect 186405 232056 186410 232112
rect 186466 232056 190164 232112
rect 186405 232054 190164 232056
rect 186405 232051 186471 232054
rect 411345 231842 411411 231845
rect 409860 231840 411411 231842
rect 409860 231784 411350 231840
rect 411406 231784 411411 231840
rect 409860 231782 411411 231784
rect 411345 231779 411411 231782
rect 186313 231026 186379 231029
rect 186313 231024 190164 231026
rect 186313 230968 186318 231024
rect 186374 230968 190164 231024
rect 186313 230966 190164 230968
rect 186313 230963 186379 230966
rect 186313 229938 186379 229941
rect 186313 229936 190164 229938
rect 186313 229880 186318 229936
rect 186374 229880 190164 229936
rect 186313 229878 190164 229880
rect 186313 229875 186379 229878
rect 411253 229802 411319 229805
rect 409860 229800 411319 229802
rect 409860 229744 411258 229800
rect 411314 229744 411319 229800
rect 409860 229742 411319 229744
rect 411253 229739 411319 229742
rect 186313 228986 186379 228989
rect 186313 228984 190164 228986
rect 186313 228928 186318 228984
rect 186374 228928 190164 228984
rect 186313 228926 190164 228928
rect 186313 228923 186379 228926
rect -960 227884 480 228124
rect 186405 227898 186471 227901
rect 409505 227898 409571 227901
rect 186405 227896 190164 227898
rect 186405 227840 186410 227896
rect 186466 227840 190164 227896
rect 186405 227838 190164 227840
rect 409462 227896 409571 227898
rect 409462 227840 409510 227896
rect 409566 227840 409571 227896
rect 186405 227835 186471 227838
rect 409462 227835 409571 227840
rect 409462 227732 409522 227835
rect 186313 226810 186379 226813
rect 186313 226808 190164 226810
rect 186313 226752 186318 226808
rect 186374 226752 190164 226808
rect 186313 226750 190164 226752
rect 186313 226747 186379 226750
rect 186313 225722 186379 225725
rect 411529 225722 411595 225725
rect 186313 225720 190164 225722
rect 186313 225664 186318 225720
rect 186374 225664 190164 225720
rect 186313 225662 190164 225664
rect 409860 225720 411595 225722
rect 409860 225664 411534 225720
rect 411590 225664 411595 225720
rect 409860 225662 411595 225664
rect 186313 225659 186379 225662
rect 411529 225659 411595 225662
rect 409454 224980 409460 225044
rect 409524 225042 409530 225044
rect 410333 225042 410399 225045
rect 409524 225040 410399 225042
rect 409524 224984 410338 225040
rect 410394 224984 410399 225040
rect 409524 224982 410399 224984
rect 409524 224980 409530 224982
rect 410333 224979 410399 224982
rect 186313 224770 186379 224773
rect 186313 224768 190164 224770
rect 186313 224712 186318 224768
rect 186374 224712 190164 224768
rect 186313 224710 190164 224712
rect 186313 224707 186379 224710
rect 186405 223682 186471 223685
rect 411253 223682 411319 223685
rect 186405 223680 190164 223682
rect 186405 223624 186410 223680
rect 186466 223624 190164 223680
rect 186405 223622 190164 223624
rect 409860 223680 411319 223682
rect 409860 223624 411258 223680
rect 411314 223624 411319 223680
rect 409860 223622 411319 223624
rect 186405 223619 186471 223622
rect 411253 223619 411319 223622
rect 186313 222594 186379 222597
rect 186313 222592 190164 222594
rect 186313 222536 186318 222592
rect 186374 222536 190164 222592
rect 186313 222534 190164 222536
rect 186313 222531 186379 222534
rect 410333 221642 410399 221645
rect 410793 221642 410859 221645
rect 409860 221640 410859 221642
rect 409860 221584 410338 221640
rect 410394 221584 410798 221640
rect 410854 221584 410859 221640
rect 409860 221582 410859 221584
rect 410333 221579 410399 221582
rect 410793 221579 410859 221582
rect 186313 221506 186379 221509
rect 186313 221504 190164 221506
rect 186313 221448 186318 221504
rect 186374 221448 190164 221504
rect 186313 221446 190164 221448
rect 186313 221443 186379 221446
rect 186497 220554 186563 220557
rect 186497 220552 190164 220554
rect 186497 220496 186502 220552
rect 186558 220496 190164 220552
rect 186497 220494 190164 220496
rect 186497 220491 186563 220494
rect 411989 219602 412055 219605
rect 409860 219600 412055 219602
rect 409860 219544 411994 219600
rect 412050 219544 412055 219600
rect 409860 219542 412055 219544
rect 411989 219539 412055 219542
rect 186405 219466 186471 219469
rect 186405 219464 190164 219466
rect 186405 219408 186410 219464
rect 186466 219408 190164 219464
rect 186405 219406 190164 219408
rect 186405 219403 186471 219406
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 186313 218378 186379 218381
rect 186313 218376 190164 218378
rect 186313 218320 186318 218376
rect 186374 218320 190164 218376
rect 186313 218318 190164 218320
rect 186313 218315 186379 218318
rect 411253 217426 411319 217429
rect 409860 217424 411319 217426
rect 409860 217368 411258 217424
rect 411314 217368 411319 217424
rect 409860 217366 411319 217368
rect 411253 217363 411319 217366
rect 186313 217290 186379 217293
rect 186313 217288 190164 217290
rect 186313 217232 186318 217288
rect 186374 217232 190164 217288
rect 186313 217230 190164 217232
rect 186313 217227 186379 217230
rect 186313 216338 186379 216341
rect 186313 216336 190164 216338
rect 186313 216280 186318 216336
rect 186374 216280 190164 216336
rect 186313 216278 190164 216280
rect 186313 216275 186379 216278
rect 411846 215386 411852 215388
rect 409860 215326 411852 215386
rect 411846 215324 411852 215326
rect 411916 215386 411922 215388
rect 412081 215386 412147 215389
rect 411916 215384 412147 215386
rect 411916 215328 412086 215384
rect 412142 215328 412147 215384
rect 411916 215326 412147 215328
rect 411916 215324 411922 215326
rect 412081 215323 412147 215326
rect 186313 215250 186379 215253
rect 186313 215248 190164 215250
rect 186313 215192 186318 215248
rect 186374 215192 190164 215248
rect 186313 215190 190164 215192
rect 186313 215187 186379 215190
rect -960 214828 480 215068
rect 186405 214162 186471 214165
rect 186405 214160 190164 214162
rect 186405 214104 186410 214160
rect 186466 214104 190164 214160
rect 186405 214102 190164 214104
rect 186405 214099 186471 214102
rect 411253 213346 411319 213349
rect 409860 213344 411319 213346
rect 409860 213288 411258 213344
rect 411314 213288 411319 213344
rect 409860 213286 411319 213288
rect 411253 213283 411319 213286
rect 186313 213074 186379 213077
rect 186313 213072 190164 213074
rect 186313 213016 186318 213072
rect 186374 213016 190164 213072
rect 186313 213014 190164 213016
rect 186313 213011 186379 213014
rect 186313 212122 186379 212125
rect 186313 212120 190164 212122
rect 186313 212064 186318 212120
rect 186374 212064 190164 212120
rect 186313 212062 190164 212064
rect 186313 212059 186379 212062
rect 411253 211306 411319 211309
rect 409860 211304 411319 211306
rect 409860 211248 411258 211304
rect 411314 211248 411319 211304
rect 409860 211246 411319 211248
rect 411253 211243 411319 211246
rect 186313 211034 186379 211037
rect 186313 211032 190164 211034
rect 186313 210976 186318 211032
rect 186374 210976 190164 211032
rect 186313 210974 190164 210976
rect 186313 210971 186379 210974
rect 186405 209946 186471 209949
rect 186405 209944 190164 209946
rect 186405 209888 186410 209944
rect 186466 209888 190164 209944
rect 186405 209886 190164 209888
rect 186405 209883 186471 209886
rect 411621 209266 411687 209269
rect 409860 209264 411687 209266
rect 409860 209208 411626 209264
rect 411682 209208 411687 209264
rect 409860 209206 411687 209208
rect 411621 209203 411687 209206
rect 186313 208858 186379 208861
rect 186313 208856 190164 208858
rect 186313 208800 186318 208856
rect 186374 208800 190164 208856
rect 186313 208798 190164 208800
rect 186313 208795 186379 208798
rect 186313 207906 186379 207909
rect 186313 207904 190164 207906
rect 186313 207848 186318 207904
rect 186374 207848 190164 207904
rect 186313 207846 190164 207848
rect 186313 207843 186379 207846
rect 411345 207226 411411 207229
rect 409860 207224 411411 207226
rect 409860 207168 411350 207224
rect 411406 207168 411411 207224
rect 409860 207166 411411 207168
rect 411345 207163 411411 207166
rect 186405 206818 186471 206821
rect 186405 206816 190164 206818
rect 186405 206760 186410 206816
rect 186466 206760 190164 206816
rect 186405 206758 190164 206760
rect 186405 206755 186471 206758
rect 186313 205730 186379 205733
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 186313 205728 190164 205730
rect 186313 205672 186318 205728
rect 186374 205672 190164 205728
rect 186313 205670 190164 205672
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 186313 205667 186379 205670
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 411253 205186 411319 205189
rect 409860 205184 411319 205186
rect 409860 205128 411258 205184
rect 411314 205128 411319 205184
rect 409860 205126 411319 205128
rect 411253 205123 411319 205126
rect 186313 204642 186379 204645
rect 186313 204640 190164 204642
rect 186313 204584 186318 204640
rect 186374 204584 190164 204640
rect 186313 204582 190164 204584
rect 186313 204579 186379 204582
rect 186313 203690 186379 203693
rect 186313 203688 190164 203690
rect 186313 203632 186318 203688
rect 186374 203632 190164 203688
rect 186313 203630 190164 203632
rect 186313 203627 186379 203630
rect 411253 203146 411319 203149
rect 409860 203144 411319 203146
rect 409860 203088 411258 203144
rect 411314 203088 411319 203144
rect 409860 203086 411319 203088
rect 411253 203083 411319 203086
rect 186313 202602 186379 202605
rect 186313 202600 190164 202602
rect 186313 202544 186318 202600
rect 186374 202544 190164 202600
rect 186313 202542 190164 202544
rect 186313 202539 186379 202542
rect -960 201772 480 202012
rect 186405 201514 186471 201517
rect 186405 201512 190164 201514
rect 186405 201456 186410 201512
rect 186466 201456 190164 201512
rect 186405 201454 190164 201456
rect 186405 201451 186471 201454
rect 411253 201106 411319 201109
rect 409860 201104 411319 201106
rect 409860 201048 411258 201104
rect 411314 201048 411319 201104
rect 409860 201046 411319 201048
rect 411253 201043 411319 201046
rect 186313 200562 186379 200565
rect 186313 200560 190164 200562
rect 186313 200504 186318 200560
rect 186374 200504 190164 200560
rect 186313 200502 190164 200504
rect 186313 200499 186379 200502
rect 399518 199548 399524 199612
rect 399588 199610 399594 199612
rect 409086 199610 409092 199612
rect 399588 199550 409092 199610
rect 399588 199548 399594 199550
rect 409086 199548 409092 199550
rect 409156 199548 409162 199612
rect 398925 199474 398991 199477
rect 411846 199474 411852 199476
rect 398925 199472 411852 199474
rect 398925 199416 398930 199472
rect 398986 199416 411852 199472
rect 398925 199414 411852 199416
rect 398925 199411 398991 199414
rect 411846 199412 411852 199414
rect 411916 199412 411922 199476
rect 399334 199276 399340 199340
rect 399404 199338 399410 199340
rect 412766 199338 412772 199340
rect 399404 199278 412772 199338
rect 399404 199276 399410 199278
rect 412766 199276 412772 199278
rect 412836 199276 412842 199340
rect 181437 198658 181503 198661
rect 403525 198658 403591 198661
rect 181437 198656 403591 198658
rect 181437 198600 181442 198656
rect 181498 198600 403530 198656
rect 403586 198600 403591 198656
rect 181437 198598 403591 198600
rect 181437 198595 181503 198598
rect 403525 198595 403591 198598
rect 180057 198522 180123 198525
rect 387793 198522 387859 198525
rect 180057 198520 387859 198522
rect 180057 198464 180062 198520
rect 180118 198464 387798 198520
rect 387854 198464 387859 198520
rect 180057 198462 387859 198464
rect 180057 198459 180123 198462
rect 387793 198459 387859 198462
rect 360101 198386 360167 198389
rect 417509 198386 417575 198389
rect 360101 198384 417575 198386
rect 360101 198328 360106 198384
rect 360162 198328 417514 198384
rect 417570 198328 417575 198384
rect 360101 198326 417575 198328
rect 360101 198323 360167 198326
rect 417509 198323 417575 198326
rect 292113 198114 292179 198117
rect 510797 198114 510863 198117
rect 292113 198112 510863 198114
rect 292113 198056 292118 198112
rect 292174 198056 510802 198112
rect 510858 198056 510863 198112
rect 292113 198054 510863 198056
rect 292113 198051 292179 198054
rect 510797 198051 510863 198054
rect 252185 197978 252251 197981
rect 510613 197978 510679 197981
rect 252185 197976 510679 197978
rect 252185 197920 252190 197976
rect 252246 197920 510618 197976
rect 510674 197920 510679 197976
rect 252185 197918 510679 197920
rect 252185 197915 252251 197918
rect 510613 197915 510679 197918
rect 398598 196556 398604 196620
rect 398668 196618 398674 196620
rect 409229 196618 409295 196621
rect 398668 196616 409295 196618
rect 398668 196560 409234 196616
rect 409290 196560 409295 196616
rect 398668 196558 409295 196560
rect 398668 196556 398674 196558
rect 409229 196555 409295 196558
rect 404353 196074 404419 196077
rect 408534 196074 408540 196076
rect 404353 196072 408540 196074
rect 404353 196016 404358 196072
rect 404414 196016 408540 196072
rect 404353 196014 408540 196016
rect 404353 196011 404419 196014
rect 408534 196012 408540 196014
rect 408604 196012 408610 196076
rect 395245 195530 395311 195533
rect 416957 195530 417023 195533
rect 395245 195528 417023 195530
rect 395245 195472 395250 195528
rect 395306 195472 416962 195528
rect 417018 195472 417023 195528
rect 395245 195470 417023 195472
rect 395245 195467 395311 195470
rect 416957 195467 417023 195470
rect 168281 195394 168347 195397
rect 409822 195394 409828 195396
rect 168281 195392 409828 195394
rect 168281 195336 168286 195392
rect 168342 195336 409828 195392
rect 168281 195334 409828 195336
rect 168281 195331 168347 195334
rect 409822 195332 409828 195334
rect 409892 195332 409898 195396
rect 167361 195258 167427 195261
rect 410006 195258 410012 195260
rect 167361 195256 410012 195258
rect 167361 195200 167366 195256
rect 167422 195200 410012 195256
rect 167361 195198 410012 195200
rect 167361 195195 167427 195198
rect 410006 195196 410012 195198
rect 410076 195196 410082 195260
rect 399702 194108 399708 194172
rect 399772 194170 399778 194172
rect 411478 194170 411484 194172
rect 399772 194110 411484 194170
rect 399772 194108 399778 194110
rect 411478 194108 411484 194110
rect 411548 194108 411554 194172
rect 168230 193972 168236 194036
rect 168300 194034 168306 194036
rect 410701 194034 410767 194037
rect 168300 194032 410767 194034
rect 168300 193976 410706 194032
rect 410762 193976 410767 194032
rect 168300 193974 410767 193976
rect 168300 193972 168306 193974
rect 410701 193971 410767 193974
rect 167310 193836 167316 193900
rect 167380 193898 167386 193900
rect 410609 193898 410675 193901
rect 167380 193896 410675 193898
rect 167380 193840 410614 193896
rect 410670 193840 410675 193896
rect 167380 193838 410675 193840
rect 167380 193836 167386 193838
rect 410609 193835 410675 193838
rect 260833 192538 260899 192541
rect 412950 192538 412956 192540
rect 260833 192536 412956 192538
rect 260833 192480 260838 192536
rect 260894 192480 412956 192536
rect 260833 192478 412956 192480
rect 260833 192475 260899 192478
rect 412950 192476 412956 192478
rect 413020 192476 413026 192540
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect -960 149684 480 149924
rect 168097 145618 168163 145621
rect 412398 145618 412404 145620
rect 168097 145616 412404 145618
rect 168097 145560 168102 145616
rect 168158 145560 412404 145616
rect 168097 145558 412404 145560
rect 168097 145555 168163 145558
rect 412398 145556 412404 145558
rect 412468 145556 412474 145620
rect 399477 144122 399543 144125
rect 411662 144122 411668 144124
rect 399477 144120 411668 144122
rect 399477 144064 399482 144120
rect 399538 144064 411668 144120
rect 399477 144062 411668 144064
rect 399477 144059 399543 144062
rect 411662 144060 411668 144062
rect 411732 144060 411738 144124
rect 400121 142762 400187 142765
rect 411294 142762 411300 142764
rect 400121 142760 411300 142762
rect 400121 142704 400126 142760
rect 400182 142704 411300 142760
rect 400121 142702 411300 142704
rect 400121 142699 400187 142702
rect 411294 142700 411300 142702
rect 411364 142700 411370 142764
rect 414606 142700 414612 142764
rect 414676 142762 414682 142764
rect 491293 142762 491359 142765
rect 414676 142760 491359 142762
rect 414676 142704 491298 142760
rect 491354 142704 491359 142760
rect 414676 142702 491359 142704
rect 414676 142700 414682 142702
rect 491293 142699 491359 142702
rect 169334 139980 169340 140044
rect 169404 140042 169410 140044
rect 392577 140042 392643 140045
rect 413829 140042 413895 140045
rect 169404 140040 392643 140042
rect 169404 139984 392582 140040
rect 392638 139984 392643 140040
rect 169404 139982 392643 139984
rect 169404 139980 169410 139982
rect 392577 139979 392643 139982
rect 402930 140040 413895 140042
rect 402930 139984 413834 140040
rect 413890 139984 413895 140040
rect 402930 139982 413895 139984
rect 168046 139844 168052 139908
rect 168116 139906 168122 139908
rect 168281 139906 168347 139909
rect 168116 139904 168347 139906
rect 168116 139848 168286 139904
rect 168342 139848 168347 139904
rect 168116 139846 168347 139848
rect 168116 139844 168122 139846
rect 168281 139843 168347 139846
rect 169518 139844 169524 139908
rect 169588 139906 169594 139908
rect 392761 139906 392827 139909
rect 402930 139906 402990 139982
rect 413829 139979 413895 139982
rect 169588 139904 392827 139906
rect 169588 139848 392766 139904
rect 392822 139848 392827 139904
rect 169588 139846 392827 139848
rect 169588 139844 169594 139846
rect 392761 139843 392827 139846
rect 400630 139846 402990 139906
rect 170305 139770 170371 139773
rect 395245 139770 395311 139773
rect 170305 139768 395311 139770
rect 170305 139712 170310 139768
rect 170366 139712 395250 139768
rect 395306 139712 395311 139768
rect 170305 139710 395311 139712
rect 170305 139707 170371 139710
rect 395245 139707 395311 139710
rect 167729 139634 167795 139637
rect 169477 139634 169543 139637
rect 167729 139632 168298 139634
rect 167729 139576 167734 139632
rect 167790 139576 168298 139632
rect 167729 139574 168298 139576
rect 167729 139571 167795 139574
rect 167678 139436 167684 139500
rect 167748 139498 167754 139500
rect 168097 139498 168163 139501
rect 167748 139496 168163 139498
rect 167748 139440 168102 139496
rect 168158 139440 168163 139496
rect 167748 139438 168163 139440
rect 168238 139498 168298 139574
rect 169477 139632 398850 139634
rect 169477 139576 169482 139632
rect 169538 139576 398850 139632
rect 169477 139574 398850 139576
rect 169477 139571 169543 139574
rect 397913 139498 397979 139501
rect 398790 139500 398850 139574
rect 398046 139498 398052 139500
rect 168238 139496 398052 139498
rect 168238 139440 397918 139496
rect 397974 139440 398052 139496
rect 168238 139438 398052 139440
rect 167748 139436 167754 139438
rect 168097 139435 168163 139438
rect 397913 139435 397979 139438
rect 398046 139436 398052 139438
rect 398116 139436 398122 139500
rect 398782 139436 398788 139500
rect 398852 139498 398858 139500
rect 399702 139498 399708 139500
rect 398852 139438 399708 139498
rect 398852 139436 398858 139438
rect 399702 139436 399708 139438
rect 399772 139436 399778 139500
rect 169845 139226 169911 139229
rect 169845 139224 170108 139226
rect 169845 139168 169850 139224
rect 169906 139168 170108 139224
rect 400630 139196 400690 139846
rect 580625 139362 580691 139365
rect 583520 139362 584960 139452
rect 580625 139360 584960 139362
rect 580625 139304 580630 139360
rect 580686 139304 584960 139360
rect 580625 139302 584960 139304
rect 580625 139299 580691 139302
rect 583520 139212 584960 139302
rect 169845 139166 170108 139168
rect 169845 139163 169911 139166
rect 168046 137532 168052 137596
rect 168116 137594 168122 137596
rect 168116 137534 170108 137594
rect 168116 137532 168122 137534
rect 398598 137532 398604 137596
rect 398668 137594 398674 137596
rect 398668 137534 400108 137594
rect 398668 137532 398674 137534
rect -960 136628 480 136868
rect 167361 136642 167427 136645
rect 167862 136642 167868 136644
rect 167361 136640 167868 136642
rect 167361 136584 167366 136640
rect 167422 136584 167868 136640
rect 167361 136582 167868 136584
rect 167361 136579 167427 136582
rect 167862 136580 167868 136582
rect 167932 136580 167938 136644
rect 167678 135900 167684 135964
rect 167748 135962 167754 135964
rect 397821 135962 397887 135965
rect 167748 135902 170108 135962
rect 397821 135960 400108 135962
rect 397821 135904 397826 135960
rect 397882 135904 400108 135960
rect 397821 135902 400108 135904
rect 167748 135900 167754 135902
rect 397821 135899 397887 135902
rect 167678 135628 167684 135692
rect 167748 135690 167754 135692
rect 170305 135690 170371 135693
rect 167748 135688 170371 135690
rect 167748 135632 170310 135688
rect 170366 135632 170371 135688
rect 167748 135630 170371 135632
rect 167748 135628 167754 135630
rect 170305 135627 170371 135630
rect 168189 134330 168255 134333
rect 397453 134330 397519 134333
rect 168189 134328 170108 134330
rect 168189 134272 168194 134328
rect 168250 134272 170108 134328
rect 168189 134270 170108 134272
rect 397453 134328 400108 134330
rect 397453 134272 397458 134328
rect 397514 134272 400108 134328
rect 397453 134270 400108 134272
rect 168189 134267 168255 134270
rect 397453 134267 397519 134270
rect 281533 133650 281599 133653
rect 512177 133650 512243 133653
rect 279926 133648 281599 133650
rect 279926 133592 281538 133648
rect 281594 133592 281599 133648
rect 279926 133590 281599 133592
rect 170213 133242 170279 133245
rect 170213 133240 170322 133242
rect 170213 133184 170218 133240
rect 170274 133184 170322 133240
rect 170213 133179 170322 133184
rect 170262 132668 170322 133179
rect 279926 133076 279986 133590
rect 281533 133587 281599 133590
rect 509926 133648 512243 133650
rect 509926 133592 512182 133648
rect 512238 133592 512243 133648
rect 509926 133590 512243 133592
rect 509926 133076 509986 133590
rect 512177 133587 512243 133590
rect 397453 132698 397519 132701
rect 397453 132696 400108 132698
rect 397453 132640 397458 132696
rect 397514 132640 400108 132696
rect 397453 132638 400108 132640
rect 397453 132635 397519 132638
rect 169753 131066 169819 131069
rect 398373 131066 398439 131069
rect 169753 131064 170108 131066
rect 169753 131008 169758 131064
rect 169814 131008 170108 131064
rect 169753 131006 170108 131008
rect 398373 131064 400108 131066
rect 398373 131008 398378 131064
rect 398434 131008 400108 131064
rect 398373 131006 400108 131008
rect 169753 131003 169819 131006
rect 398373 131003 398439 131006
rect 169150 129372 169156 129436
rect 169220 129434 169226 129436
rect 397453 129434 397519 129437
rect 169220 129374 170108 129434
rect 397453 129432 400108 129434
rect 397453 129376 397458 129432
rect 397514 129376 400108 129432
rect 397453 129374 400108 129376
rect 169220 129372 169226 129374
rect 397453 129371 397519 129374
rect 167862 127740 167868 127804
rect 167932 127802 167938 127804
rect 399569 127802 399635 127805
rect 167932 127742 170108 127802
rect 399569 127800 400108 127802
rect 399569 127744 399574 127800
rect 399630 127744 400108 127800
rect 399569 127742 400108 127744
rect 167932 127740 167938 127742
rect 399569 127739 399635 127742
rect 400581 126714 400647 126717
rect 400581 126712 400690 126714
rect 400581 126656 400586 126712
rect 400642 126656 400690 126712
rect 400581 126651 400690 126656
rect 168833 126170 168899 126173
rect 168833 126168 170108 126170
rect 168833 126112 168838 126168
rect 168894 126112 170108 126168
rect 400630 126140 400690 126651
rect 168833 126110 170108 126112
rect 168833 126107 168899 126110
rect 579705 126034 579771 126037
rect 583520 126034 584960 126124
rect 579705 126032 584960 126034
rect 579705 125976 579710 126032
rect 579766 125976 584960 126032
rect 579705 125974 584960 125976
rect 579705 125971 579771 125974
rect 583520 125884 584960 125974
rect 168925 124538 168991 124541
rect 397453 124538 397519 124541
rect 168925 124536 170108 124538
rect 168925 124480 168930 124536
rect 168986 124480 170108 124536
rect 168925 124478 170108 124480
rect 397453 124536 400108 124538
rect 397453 124480 397458 124536
rect 397514 124480 400108 124536
rect 397453 124478 400108 124480
rect 168925 124475 168991 124478
rect 397453 124475 397519 124478
rect -960 123572 480 123812
rect 167310 122844 167316 122908
rect 167380 122906 167386 122908
rect 397453 122906 397519 122909
rect 167380 122846 170108 122906
rect 397453 122904 400108 122906
rect 397453 122848 397458 122904
rect 397514 122848 400108 122904
rect 397453 122846 400108 122848
rect 167380 122844 167386 122846
rect 397453 122843 397519 122846
rect 400581 121410 400647 121413
rect 400581 121408 400690 121410
rect 400581 121352 400586 121408
rect 400642 121352 400690 121408
rect 400581 121347 400690 121352
rect 168230 121212 168236 121276
rect 168300 121274 168306 121276
rect 168300 121214 170108 121274
rect 400630 121244 400690 121347
rect 168300 121212 168306 121214
rect 282453 119914 282519 119917
rect 512085 119914 512151 119917
rect 279926 119912 282519 119914
rect 279926 119856 282458 119912
rect 282514 119856 282519 119912
rect 279926 119854 282519 119856
rect 169201 119642 169267 119645
rect 169201 119640 170108 119642
rect 169201 119584 169206 119640
rect 169262 119584 170108 119640
rect 169201 119582 170108 119584
rect 169201 119579 169267 119582
rect 279926 119340 279986 119854
rect 282453 119851 282519 119854
rect 509926 119912 512151 119914
rect 509926 119856 512090 119912
rect 512146 119856 512151 119912
rect 509926 119854 512151 119856
rect 397453 119642 397519 119645
rect 397453 119640 400108 119642
rect 397453 119584 397458 119640
rect 397514 119584 400108 119640
rect 397453 119582 400108 119584
rect 397453 119579 397519 119582
rect 509926 119340 509986 119854
rect 512085 119851 512151 119854
rect 166901 117874 166967 117877
rect 398097 117874 398163 117877
rect 166901 117872 170108 117874
rect 166901 117816 166906 117872
rect 166962 117816 170108 117872
rect 166901 117814 170108 117816
rect 398097 117872 400108 117874
rect 398097 117816 398102 117872
rect 398158 117816 400108 117872
rect 398097 117814 400108 117816
rect 166901 117811 166967 117814
rect 398097 117811 398163 117814
rect 169109 116242 169175 116245
rect 397821 116242 397887 116245
rect 169109 116240 170108 116242
rect 169109 116184 169114 116240
rect 169170 116184 170108 116240
rect 169109 116182 170108 116184
rect 397821 116240 400108 116242
rect 397821 116184 397826 116240
rect 397882 116184 400108 116240
rect 397821 116182 400108 116184
rect 169109 116179 169175 116182
rect 397821 116179 397887 116182
rect 168281 114610 168347 114613
rect 398005 114610 398071 114613
rect 168281 114608 170108 114610
rect 168281 114552 168286 114608
rect 168342 114552 170108 114608
rect 168281 114550 170108 114552
rect 398005 114608 400108 114610
rect 398005 114552 398010 114608
rect 398066 114552 400108 114608
rect 398005 114550 400108 114552
rect 168281 114547 168347 114550
rect 398005 114547 398071 114550
rect 169293 112978 169359 112981
rect 397545 112978 397611 112981
rect 169293 112976 170108 112978
rect 169293 112920 169298 112976
rect 169354 112920 170108 112976
rect 169293 112918 170108 112920
rect 397545 112976 400108 112978
rect 397545 112920 397550 112976
rect 397606 112920 400108 112976
rect 397545 112918 400108 112920
rect 169293 112915 169359 112918
rect 397545 112915 397611 112918
rect 579705 112842 579771 112845
rect 583520 112842 584960 112932
rect 579705 112840 584960 112842
rect 579705 112784 579710 112840
rect 579766 112784 584960 112840
rect 579705 112782 584960 112784
rect 579705 112779 579771 112782
rect 583520 112692 584960 112782
rect 167637 111346 167703 111349
rect 398833 111346 398899 111349
rect 167637 111344 170108 111346
rect 167637 111288 167642 111344
rect 167698 111288 170108 111344
rect 167637 111286 170108 111288
rect 398833 111344 400108 111346
rect 398833 111288 398838 111344
rect 398894 111288 400108 111344
rect 398833 111286 400108 111288
rect 167637 111283 167703 111286
rect 398833 111283 398899 111286
rect -960 110516 480 110756
rect 169385 109714 169451 109717
rect 398189 109714 398255 109717
rect 169385 109712 170108 109714
rect 169385 109656 169390 109712
rect 169446 109656 170108 109712
rect 169385 109654 170108 109656
rect 398189 109712 400108 109714
rect 398189 109656 398194 109712
rect 398250 109656 400108 109712
rect 398189 109654 400108 109656
rect 169385 109651 169451 109654
rect 398189 109651 398255 109654
rect 169477 108082 169543 108085
rect 169477 108080 170108 108082
rect 169477 108024 169482 108080
rect 169538 108024 170108 108080
rect 169477 108022 170108 108024
rect 169477 108019 169543 108022
rect 398782 108020 398788 108084
rect 398852 108082 398858 108084
rect 398852 108022 400108 108082
rect 398852 108020 398858 108022
rect 167729 106450 167795 106453
rect 167729 106448 170108 106450
rect 167729 106392 167734 106448
rect 167790 106392 170108 106448
rect 167729 106390 170108 106392
rect 167729 106387 167795 106390
rect 398046 106388 398052 106452
rect 398116 106450 398122 106452
rect 398116 106390 400108 106450
rect 398116 106388 398122 106390
rect 282361 106178 282427 106181
rect 510797 106178 510863 106181
rect 279926 106176 282427 106178
rect 279926 106120 282366 106176
rect 282422 106120 282427 106176
rect 279926 106118 282427 106120
rect 279926 105604 279986 106118
rect 282361 106115 282427 106118
rect 509926 106176 510863 106178
rect 509926 106120 510802 106176
rect 510858 106120 510863 106176
rect 509926 106118 510863 106120
rect 509926 105604 509986 106118
rect 510797 106115 510863 106118
rect 170121 104954 170187 104957
rect 170078 104952 170187 104954
rect 170078 104896 170126 104952
rect 170182 104896 170187 104952
rect 170078 104891 170187 104896
rect 170078 104788 170138 104891
rect 397453 104818 397519 104821
rect 397453 104816 400108 104818
rect 397453 104760 397458 104816
rect 397514 104760 400108 104816
rect 397453 104758 400108 104760
rect 397453 104755 397519 104758
rect 170029 103322 170095 103325
rect 400213 103322 400279 103325
rect 170029 103320 170138 103322
rect 170029 103264 170034 103320
rect 170090 103264 170138 103320
rect 170029 103259 170138 103264
rect 400213 103320 400322 103322
rect 400213 103264 400218 103320
rect 400274 103264 400322 103320
rect 400213 103259 400322 103264
rect 170078 103156 170138 103259
rect 400262 103156 400322 103259
rect 169569 101554 169635 101557
rect 397453 101554 397519 101557
rect 169569 101552 170108 101554
rect 169569 101496 169574 101552
rect 169630 101496 170108 101552
rect 169569 101494 170108 101496
rect 397453 101552 400108 101554
rect 397453 101496 397458 101552
rect 397514 101496 400108 101552
rect 397453 101494 400108 101496
rect 169569 101491 169635 101494
rect 397453 101491 397519 101494
rect 169661 99922 169727 99925
rect 398373 99922 398439 99925
rect 169661 99920 170108 99922
rect 169661 99864 169666 99920
rect 169722 99864 170108 99920
rect 169661 99862 170108 99864
rect 398373 99920 400108 99922
rect 398373 99864 398378 99920
rect 398434 99864 400108 99920
rect 398373 99862 400108 99864
rect 169661 99859 169727 99862
rect 398373 99859 398439 99862
rect 580533 99514 580599 99517
rect 583520 99514 584960 99604
rect 580533 99512 584960 99514
rect 580533 99456 580538 99512
rect 580594 99456 584960 99512
rect 580533 99454 584960 99456
rect 580533 99451 580599 99454
rect 583520 99364 584960 99454
rect 167821 98290 167887 98293
rect 397453 98290 397519 98293
rect 167821 98288 170108 98290
rect 167821 98232 167826 98288
rect 167882 98232 170108 98288
rect 167821 98230 170108 98232
rect 397453 98288 400108 98290
rect 397453 98232 397458 98288
rect 397514 98232 400108 98288
rect 397453 98230 400108 98232
rect 167821 98227 167887 98230
rect 397453 98227 397519 98230
rect -960 97460 480 97700
rect 166993 96522 167059 96525
rect 396809 96522 396875 96525
rect 166993 96520 170108 96522
rect 166993 96464 166998 96520
rect 167054 96464 170108 96520
rect 166993 96462 170108 96464
rect 396809 96520 400108 96522
rect 396809 96464 396814 96520
rect 396870 96464 400108 96520
rect 396809 96462 400108 96464
rect 166993 96459 167059 96462
rect 396809 96459 396875 96462
rect 169937 95162 170003 95165
rect 169937 95160 170138 95162
rect 169937 95104 169942 95160
rect 169998 95104 170138 95160
rect 169937 95102 170138 95104
rect 169937 95099 170003 95102
rect 170078 94860 170138 95102
rect 397453 94890 397519 94893
rect 397453 94888 400108 94890
rect 397453 94832 397458 94888
rect 397514 94832 400108 94888
rect 397453 94830 400108 94832
rect 397453 94827 397519 94830
rect 169518 93196 169524 93260
rect 169588 93258 169594 93260
rect 398097 93258 398163 93261
rect 169588 93198 170108 93258
rect 398097 93256 400108 93258
rect 398097 93200 398102 93256
rect 398158 93200 400108 93256
rect 398097 93198 400108 93200
rect 169588 93196 169594 93198
rect 398097 93195 398163 93198
rect 280245 92442 280311 92445
rect 511993 92442 512059 92445
rect 279926 92440 280311 92442
rect 279926 92384 280250 92440
rect 280306 92384 280311 92440
rect 279926 92382 280311 92384
rect 279926 91868 279986 92382
rect 280245 92379 280311 92382
rect 509926 92440 512059 92442
rect 509926 92384 511998 92440
rect 512054 92384 512059 92440
rect 509926 92382 512059 92384
rect 509926 91868 509986 92382
rect 511993 92379 512059 92382
rect 169334 91564 169340 91628
rect 169404 91626 169410 91628
rect 397453 91626 397519 91629
rect 169404 91566 170108 91626
rect 397453 91624 400108 91626
rect 397453 91568 397458 91624
rect 397514 91568 400108 91624
rect 397453 91566 400108 91568
rect 169404 91564 169410 91566
rect 397453 91563 397519 91566
rect 167913 89994 167979 89997
rect 397913 89994 397979 89997
rect 167913 89992 170108 89994
rect 167913 89936 167918 89992
rect 167974 89936 170108 89992
rect 167913 89934 170108 89936
rect 397913 89992 400108 89994
rect 397913 89936 397918 89992
rect 397974 89936 400108 89992
rect 397913 89934 400108 89936
rect 167913 89931 167979 89934
rect 397913 89931 397979 89934
rect 168005 88362 168071 88365
rect 397453 88362 397519 88365
rect 168005 88360 170108 88362
rect 168005 88304 168010 88360
rect 168066 88304 170108 88360
rect 168005 88302 170108 88304
rect 397453 88360 400108 88362
rect 397453 88304 397458 88360
rect 397514 88304 400108 88360
rect 397453 88302 400108 88304
rect 168005 88299 168071 88302
rect 397453 88299 397519 88302
rect 168189 86730 168255 86733
rect 397729 86730 397795 86733
rect 168189 86728 170108 86730
rect 168189 86672 168194 86728
rect 168250 86672 170108 86728
rect 168189 86670 170108 86672
rect 397729 86728 400108 86730
rect 397729 86672 397734 86728
rect 397790 86672 400108 86728
rect 397729 86670 400108 86672
rect 168189 86667 168255 86670
rect 397729 86667 397795 86670
rect 579981 86186 580047 86189
rect 583520 86186 584960 86276
rect 579981 86184 584960 86186
rect 579981 86128 579986 86184
rect 580042 86128 584960 86184
rect 579981 86126 584960 86128
rect 579981 86123 580047 86126
rect 583520 86036 584960 86126
rect 167678 85036 167684 85100
rect 167748 85098 167754 85100
rect 397545 85098 397611 85101
rect 167748 85038 170108 85098
rect 397545 85096 400108 85098
rect 397545 85040 397550 85096
rect 397606 85040 400108 85096
rect 397545 85038 400108 85040
rect 167748 85036 167754 85038
rect 397545 85035 397611 85038
rect -960 84540 480 84780
rect 168097 83466 168163 83469
rect 399569 83466 399635 83469
rect 168097 83464 170108 83466
rect 168097 83408 168102 83464
rect 168158 83408 170108 83464
rect 168097 83406 170108 83408
rect 399569 83464 400108 83466
rect 399569 83408 399574 83464
rect 399630 83408 400108 83464
rect 399569 83406 400108 83408
rect 168097 83403 168163 83406
rect 399569 83403 399635 83406
rect 168097 81834 168163 81837
rect 397453 81834 397519 81837
rect 168097 81832 170108 81834
rect 168097 81776 168102 81832
rect 168158 81776 170108 81832
rect 168097 81774 170108 81776
rect 397453 81832 400108 81834
rect 397453 81776 397458 81832
rect 397514 81776 400108 81832
rect 397453 81774 400108 81776
rect 168097 81771 168163 81774
rect 397453 81771 397519 81774
rect 167453 80202 167519 80205
rect 398189 80202 398255 80205
rect 167453 80200 170108 80202
rect 167453 80144 167458 80200
rect 167514 80144 170108 80200
rect 167453 80142 170108 80144
rect 398189 80200 400108 80202
rect 398189 80144 398194 80200
rect 398250 80144 400108 80200
rect 398189 80142 400108 80144
rect 167453 80139 167519 80142
rect 398189 80139 398255 80142
rect 168230 78508 168236 78572
rect 168300 78570 168306 78572
rect 282177 78570 282243 78573
rect 168300 78510 170108 78570
rect 279926 78568 282243 78570
rect 279926 78512 282182 78568
rect 282238 78512 282243 78568
rect 279926 78510 282243 78512
rect 168300 78508 168306 78510
rect 279926 78132 279986 78510
rect 282177 78507 282243 78510
rect 397453 78570 397519 78573
rect 510613 78570 510679 78573
rect 397453 78568 400108 78570
rect 397453 78512 397458 78568
rect 397514 78512 400108 78568
rect 397453 78510 400108 78512
rect 509926 78568 510679 78570
rect 509926 78512 510618 78568
rect 510674 78512 510679 78568
rect 509926 78510 510679 78512
rect 397453 78507 397519 78510
rect 509926 78132 509986 78510
rect 510613 78507 510679 78510
rect 168189 76938 168255 76941
rect 398005 76938 398071 76941
rect 398833 76938 398899 76941
rect 168189 76936 170108 76938
rect 168189 76880 168194 76936
rect 168250 76880 170108 76936
rect 168189 76878 170108 76880
rect 398005 76936 400108 76938
rect 398005 76880 398010 76936
rect 398066 76880 398838 76936
rect 398894 76880 400108 76936
rect 398005 76878 400108 76880
rect 168189 76875 168255 76878
rect 398005 76875 398071 76878
rect 398833 76875 398899 76878
rect 168005 75306 168071 75309
rect 398097 75306 398163 75309
rect 168005 75304 170108 75306
rect 168005 75248 168010 75304
rect 168066 75248 170108 75304
rect 168005 75246 170108 75248
rect 398097 75304 400108 75306
rect 398097 75248 398102 75304
rect 398158 75248 400108 75304
rect 398097 75246 400108 75248
rect 168005 75243 168071 75246
rect 398097 75243 398163 75246
rect 167269 73538 167335 73541
rect 398189 73538 398255 73541
rect 167269 73536 170108 73538
rect 167269 73480 167274 73536
rect 167330 73480 170108 73536
rect 167269 73478 170108 73480
rect 398189 73536 400108 73538
rect 398189 73480 398194 73536
rect 398250 73480 400108 73536
rect 398189 73478 400108 73480
rect 167269 73475 167335 73478
rect 398189 73475 398255 73478
rect 580441 72994 580507 72997
rect 583520 72994 584960 73084
rect 580441 72992 584960 72994
rect 580441 72936 580446 72992
rect 580502 72936 584960 72992
rect 580441 72934 584960 72936
rect 580441 72931 580507 72934
rect 583520 72844 584960 72934
rect 167637 71906 167703 71909
rect 397913 71906 397979 71909
rect 398281 71906 398347 71909
rect 167637 71904 170108 71906
rect 167637 71848 167642 71904
rect 167698 71848 170108 71904
rect 167637 71846 170108 71848
rect 397913 71904 400108 71906
rect 397913 71848 397918 71904
rect 397974 71848 398286 71904
rect 398342 71848 400108 71904
rect 397913 71846 400108 71848
rect 167637 71843 167703 71846
rect 397913 71843 397979 71846
rect 398281 71843 398347 71846
rect -960 71484 480 71724
rect 400581 70410 400647 70413
rect 400078 70408 400647 70410
rect 400078 70352 400586 70408
rect 400642 70352 400647 70408
rect 400078 70350 400647 70352
rect 167913 70274 167979 70277
rect 398281 70274 398347 70277
rect 400078 70274 400138 70350
rect 400581 70347 400647 70350
rect 167913 70272 170108 70274
rect 167913 70216 167918 70272
rect 167974 70216 170108 70272
rect 167913 70214 170108 70216
rect 398281 70272 400138 70274
rect 398281 70216 398286 70272
rect 398342 70244 400138 70272
rect 398342 70216 400108 70244
rect 398281 70214 400108 70216
rect 167913 70211 167979 70214
rect 398281 70211 398347 70214
rect 167729 68642 167795 68645
rect 398373 68642 398439 68645
rect 399201 68642 399267 68645
rect 167729 68640 170108 68642
rect 167729 68584 167734 68640
rect 167790 68584 170108 68640
rect 167729 68582 170108 68584
rect 398373 68640 400108 68642
rect 398373 68584 398378 68640
rect 398434 68584 399206 68640
rect 399262 68584 400108 68640
rect 398373 68582 400108 68584
rect 167729 68579 167795 68582
rect 398373 68579 398439 68582
rect 399201 68579 399267 68582
rect 169753 67010 169819 67013
rect 397453 67010 397519 67013
rect 169753 67008 170108 67010
rect 169753 66952 169758 67008
rect 169814 66952 170108 67008
rect 169753 66950 170108 66952
rect 397453 67008 400108 67010
rect 397453 66952 397458 67008
rect 397514 66952 400108 67008
rect 397453 66950 400108 66952
rect 169753 66947 169819 66950
rect 397453 66947 397519 66950
rect 168281 65378 168347 65381
rect 398465 65378 398531 65381
rect 168281 65376 170108 65378
rect 168281 65320 168286 65376
rect 168342 65320 170108 65376
rect 168281 65318 170108 65320
rect 398465 65376 400108 65378
rect 398465 65320 398470 65376
rect 398526 65320 400108 65376
rect 398465 65318 400108 65320
rect 168281 65315 168347 65318
rect 398465 65315 398531 65318
rect 282269 64698 282335 64701
rect 510889 64698 510955 64701
rect 279926 64696 282335 64698
rect 279926 64640 282274 64696
rect 282330 64640 282335 64696
rect 279926 64638 282335 64640
rect 279926 64396 279986 64638
rect 282269 64635 282335 64638
rect 509926 64696 510955 64698
rect 509926 64640 510894 64696
rect 510950 64640 510955 64696
rect 509926 64638 510955 64640
rect 509926 64396 509986 64638
rect 510889 64635 510955 64638
rect 168046 63684 168052 63748
rect 168116 63746 168122 63748
rect 168116 63686 170108 63746
rect 168116 63684 168122 63686
rect 400078 63610 400138 63716
rect 398790 63550 400138 63610
rect 394417 63474 394483 63477
rect 397862 63474 397868 63476
rect 394417 63472 397868 63474
rect 394417 63416 394422 63472
rect 394478 63416 397868 63472
rect 394417 63414 397868 63416
rect 394417 63411 394483 63414
rect 397862 63412 397868 63414
rect 397932 63474 397938 63476
rect 398790 63474 398850 63550
rect 397932 63414 398850 63474
rect 397932 63412 397938 63414
rect 169661 62114 169727 62117
rect 399201 62114 399267 62117
rect 399477 62114 399543 62117
rect 169661 62112 170108 62114
rect 169661 62056 169666 62112
rect 169722 62056 170108 62112
rect 169661 62054 170108 62056
rect 399201 62112 400108 62114
rect 399201 62056 399206 62112
rect 399262 62056 399482 62112
rect 399538 62056 400108 62112
rect 399201 62054 400108 62056
rect 169661 62051 169727 62054
rect 399201 62051 399267 62054
rect 399477 62051 399543 62054
rect 167678 60420 167684 60484
rect 167748 60482 167754 60484
rect 397453 60482 397519 60485
rect 167748 60422 170108 60482
rect 397453 60480 400108 60482
rect 397453 60424 397458 60480
rect 397514 60424 400108 60480
rect 397453 60422 400108 60424
rect 167748 60420 167754 60422
rect 397453 60419 397519 60422
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect 393129 59258 393195 59261
rect 397453 59258 397519 59261
rect 397678 59258 397684 59260
rect 393129 59256 397684 59258
rect 393129 59200 393134 59256
rect 393190 59200 397458 59256
rect 397514 59200 397684 59256
rect 393129 59198 397684 59200
rect 393129 59195 393195 59198
rect 397453 59195 397519 59198
rect 397678 59196 397684 59198
rect 397748 59196 397754 59260
rect 169477 58850 169543 58853
rect 398557 58850 398623 58853
rect 169477 58848 170108 58850
rect 169477 58792 169482 58848
rect 169538 58792 170108 58848
rect 169477 58790 170108 58792
rect 398557 58848 400108 58850
rect 398557 58792 398562 58848
rect 398618 58792 400108 58848
rect 398557 58790 400108 58792
rect 169477 58787 169543 58790
rect 398557 58787 398623 58790
rect -960 58428 480 58668
rect 167862 57156 167868 57220
rect 167932 57218 167938 57220
rect 397453 57218 397519 57221
rect 167932 57158 170108 57218
rect 397453 57216 400108 57218
rect 397453 57160 397458 57216
rect 397514 57160 400108 57216
rect 397453 57158 400108 57160
rect 167932 57156 167938 57158
rect 397453 57155 397519 57158
rect 169569 55586 169635 55589
rect 399109 55586 399175 55589
rect 169569 55584 170108 55586
rect 169569 55528 169574 55584
rect 169630 55528 170108 55584
rect 169569 55526 170108 55528
rect 399109 55584 400108 55586
rect 399109 55528 399114 55584
rect 399170 55528 400108 55584
rect 399109 55526 400108 55528
rect 169569 55523 169635 55526
rect 399109 55523 399175 55526
rect 167361 53954 167427 53957
rect 396993 53954 397059 53957
rect 167361 53952 170108 53954
rect 167361 53896 167366 53952
rect 167422 53896 170108 53952
rect 167361 53894 170108 53896
rect 396993 53952 400108 53954
rect 396993 53896 396998 53952
rect 397054 53896 400108 53952
rect 396993 53894 400108 53896
rect 167361 53891 167427 53894
rect 396993 53891 397059 53894
rect 169385 52186 169451 52189
rect 398649 52186 398715 52189
rect 169385 52184 170108 52186
rect 169385 52128 169390 52184
rect 169446 52128 170108 52184
rect 169385 52126 170108 52128
rect 398649 52184 400108 52186
rect 398649 52128 398654 52184
rect 398710 52128 400108 52184
rect 398649 52126 400108 52128
rect 169385 52123 169451 52126
rect 398649 52123 398715 52126
rect 512269 50962 512335 50965
rect 509926 50960 512335 50962
rect 509926 50904 512274 50960
rect 512330 50904 512335 50960
rect 509926 50902 512335 50904
rect 282821 50826 282887 50829
rect 279926 50824 282887 50826
rect 279926 50768 282826 50824
rect 282882 50768 282887 50824
rect 279926 50766 282887 50768
rect 279926 50660 279986 50766
rect 282821 50763 282887 50766
rect 509926 50660 509986 50902
rect 512269 50899 512335 50902
rect 169845 50554 169911 50557
rect 397913 50554 397979 50557
rect 399385 50554 399451 50557
rect 169845 50552 170108 50554
rect 169845 50496 169850 50552
rect 169906 50496 170108 50552
rect 169845 50494 170108 50496
rect 397913 50552 400108 50554
rect 397913 50496 397918 50552
rect 397974 50496 399390 50552
rect 399446 50496 400108 50552
rect 397913 50494 400108 50496
rect 169845 50491 169911 50494
rect 397913 50491 397979 50494
rect 399385 50491 399451 50494
rect 167545 48922 167611 48925
rect 397453 48922 397519 48925
rect 167545 48920 170108 48922
rect 167545 48864 167550 48920
rect 167606 48864 170108 48920
rect 167545 48862 170108 48864
rect 397453 48920 400108 48922
rect 397453 48864 397458 48920
rect 397514 48864 400108 48920
rect 397453 48862 400108 48864
rect 167545 48859 167611 48862
rect 397453 48859 397519 48862
rect 167453 47290 167519 47293
rect 397453 47290 397519 47293
rect 398741 47290 398807 47293
rect 167453 47288 170108 47290
rect 167453 47232 167458 47288
rect 167514 47232 170108 47288
rect 167453 47230 170108 47232
rect 397453 47288 400108 47290
rect 397453 47232 397458 47288
rect 397514 47232 398746 47288
rect 398802 47232 400108 47288
rect 397453 47230 400108 47232
rect 167453 47227 167519 47230
rect 397453 47227 397519 47230
rect 398741 47227 398807 47230
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect 169937 45794 170003 45797
rect 169937 45792 170138 45794
rect 169937 45736 169942 45792
rect 169998 45736 170138 45792
rect 169937 45734 170138 45736
rect 169937 45731 170003 45734
rect 170078 45628 170138 45734
rect 398741 45658 398807 45661
rect 398741 45656 400108 45658
rect -960 45372 480 45612
rect 398741 45600 398746 45656
rect 398802 45600 400108 45656
rect 398741 45598 400108 45600
rect 398741 45595 398807 45598
rect 167177 44026 167243 44029
rect 397177 44026 397243 44029
rect 167177 44024 170108 44026
rect 167177 43968 167182 44024
rect 167238 43968 170108 44024
rect 167177 43966 170108 43968
rect 397177 44024 400108 44026
rect 397177 43968 397182 44024
rect 397238 43968 400108 44024
rect 397177 43966 400108 43968
rect 167177 43963 167243 43966
rect 397177 43963 397243 43966
rect 397453 42394 397519 42397
rect 398833 42394 398899 42397
rect 397453 42392 400108 42394
rect 167821 41850 167887 41853
rect 170078 41850 170138 42364
rect 397453 42336 397458 42392
rect 397514 42336 398838 42392
rect 398894 42336 400108 42392
rect 397453 42334 400108 42336
rect 397453 42331 397519 42334
rect 398833 42331 398899 42334
rect 167821 41848 170138 41850
rect 167821 41792 167826 41848
rect 167882 41792 170138 41848
rect 167821 41790 170138 41792
rect 167821 41787 167887 41790
rect 168281 41444 168347 41445
rect 168230 41442 168236 41444
rect 168190 41382 168236 41442
rect 168300 41440 168347 41444
rect 168342 41384 168347 41440
rect 168230 41380 168236 41382
rect 168300 41380 168347 41384
rect 168281 41379 168347 41380
rect 168230 40700 168236 40764
rect 168300 40762 168306 40764
rect 397453 40762 397519 40765
rect 168300 40702 170108 40762
rect 397453 40760 400108 40762
rect 397453 40704 397458 40760
rect 397514 40704 400108 40760
rect 397453 40702 400108 40704
rect 168300 40700 168306 40702
rect 397453 40699 397519 40702
rect 168281 39946 168347 39949
rect 168966 39946 168972 39948
rect 168281 39944 168972 39946
rect 168281 39888 168286 39944
rect 168342 39888 168972 39944
rect 168281 39886 168972 39888
rect 168281 39883 168347 39886
rect 168966 39884 168972 39886
rect 169036 39884 169042 39948
rect 168005 39130 168071 39133
rect 397453 39130 397519 39133
rect 168005 39128 170108 39130
rect 168005 39072 168010 39128
rect 168066 39072 170108 39128
rect 168005 39070 170108 39072
rect 397453 39128 400108 39130
rect 397453 39072 397458 39128
rect 397514 39072 400108 39128
rect 397453 39070 400108 39072
rect 168005 39067 168071 39070
rect 397453 39067 397519 39070
rect 168281 37498 168347 37501
rect 397545 37498 397611 37501
rect 399293 37498 399359 37501
rect 168281 37496 170108 37498
rect 168281 37440 168286 37496
rect 168342 37440 170108 37496
rect 168281 37438 170108 37440
rect 397545 37496 400108 37498
rect 397545 37440 397550 37496
rect 397606 37440 399298 37496
rect 399354 37440 400108 37496
rect 397545 37438 400108 37440
rect 168281 37435 168347 37438
rect 397545 37435 397611 37438
rect 399293 37435 399359 37438
rect 280153 37226 280219 37229
rect 279926 37224 280219 37226
rect 279926 37168 280158 37224
rect 280214 37168 280219 37224
rect 279926 37166 280219 37168
rect 279926 36924 279986 37166
rect 280153 37163 280219 37166
rect 509509 37226 509575 37229
rect 509509 37224 509618 37226
rect 509509 37168 509514 37224
rect 509570 37168 509618 37224
rect 509509 37163 509618 37168
rect 509558 36924 509618 37163
rect 399753 35866 399819 35869
rect 399753 35864 400108 35866
rect 168281 35322 168347 35325
rect 170078 35322 170138 35836
rect 399753 35808 399758 35864
rect 399814 35808 400108 35864
rect 399753 35806 400108 35808
rect 399753 35803 399819 35806
rect 168281 35320 170138 35322
rect 168281 35264 168286 35320
rect 168342 35264 170138 35320
rect 168281 35262 170138 35264
rect 168281 35259 168347 35262
rect 397453 34234 397519 34237
rect 397453 34232 400108 34234
rect 170630 33693 170690 34204
rect 397453 34176 397458 34232
rect 397514 34176 400108 34232
rect 397453 34174 400108 34176
rect 397453 34171 397519 34174
rect 170581 33688 170690 33693
rect 170581 33632 170586 33688
rect 170642 33632 170690 33688
rect 170581 33630 170690 33632
rect 170581 33627 170647 33630
rect 397361 33146 397427 33149
rect 397494 33146 397500 33148
rect 397361 33144 397500 33146
rect 397361 33088 397366 33144
rect 397422 33088 397500 33144
rect 397361 33086 397500 33088
rect 397361 33083 397427 33086
rect 397494 33084 397500 33086
rect 397564 33084 397570 33148
rect 583520 32996 584960 33236
rect 397453 32602 397519 32605
rect 397453 32600 400108 32602
rect -960 32316 480 32556
rect 170446 32061 170506 32572
rect 397453 32544 397458 32600
rect 397514 32544 400108 32600
rect 397453 32542 400108 32544
rect 397453 32539 397519 32542
rect 170446 32056 170555 32061
rect 170446 32000 170494 32056
rect 170550 32000 170555 32056
rect 170446 31998 170555 32000
rect 170489 31995 170555 31998
rect 170397 31106 170463 31109
rect 170397 31104 170506 31106
rect 170397 31048 170402 31104
rect 170458 31048 170506 31104
rect 170397 31043 170506 31048
rect 170446 30940 170506 31043
rect 397453 30970 397519 30973
rect 397453 30968 400108 30970
rect 397453 30912 397458 30968
rect 397514 30912 400108 30968
rect 397453 30910 400108 30912
rect 397453 30907 397519 30910
rect 168046 30636 168052 30700
rect 168116 30698 168122 30700
rect 397862 30698 397868 30700
rect 168116 30638 397868 30698
rect 168116 30636 168122 30638
rect 397862 30636 397868 30638
rect 397932 30636 397938 30700
rect 170581 30290 170647 30293
rect 397494 30290 397500 30292
rect 170581 30288 397500 30290
rect 170581 30232 170586 30288
rect 170642 30232 397500 30288
rect 170581 30230 397500 30232
rect 170581 30227 170647 30230
rect 397494 30228 397500 30230
rect 397564 30228 397570 30292
rect 168966 30092 168972 30156
rect 169036 30154 169042 30156
rect 393957 30154 394023 30157
rect 169036 30152 394023 30154
rect 169036 30096 393962 30152
rect 394018 30096 394023 30152
rect 169036 30094 394023 30096
rect 169036 30092 169042 30094
rect 393957 30091 394023 30094
rect 167862 29956 167868 30020
rect 167932 30018 167938 30020
rect 280797 30018 280863 30021
rect 167932 30016 280863 30018
rect 167932 29960 280802 30016
rect 280858 29960 280863 30016
rect 167932 29958 280863 29960
rect 167932 29956 167938 29958
rect 280797 29955 280863 29958
rect 168230 29820 168236 29884
rect 168300 29882 168306 29884
rect 280981 29882 281047 29885
rect 168300 29880 281047 29882
rect 168300 29824 280986 29880
rect 281042 29824 281047 29880
rect 168300 29822 281047 29824
rect 168300 29820 168306 29822
rect 280981 29819 281047 29822
rect 170489 29746 170555 29749
rect 279325 29746 279391 29749
rect 170489 29744 279391 29746
rect 170489 29688 170494 29744
rect 170550 29688 279330 29744
rect 279386 29688 279391 29744
rect 170489 29686 279391 29688
rect 170489 29683 170555 29686
rect 279325 29683 279391 29686
rect 78673 28930 78739 28933
rect 454677 28930 454743 28933
rect 78673 28928 454743 28930
rect 78673 28872 78678 28928
rect 78734 28872 454682 28928
rect 454738 28872 454743 28928
rect 78673 28870 454743 28872
rect 78673 28867 78739 28870
rect 454677 28867 454743 28870
rect 191465 28794 191531 28797
rect 556797 28794 556863 28797
rect 191465 28792 556863 28794
rect 191465 28736 191470 28792
rect 191526 28736 556802 28792
rect 556858 28736 556863 28792
rect 191465 28734 556863 28736
rect 191465 28731 191531 28734
rect 556797 28731 556863 28734
rect 199837 28658 199903 28661
rect 551369 28658 551435 28661
rect 199837 28656 551435 28658
rect 199837 28600 199842 28656
rect 199898 28600 551374 28656
rect 551430 28600 551435 28656
rect 199837 28598 551435 28600
rect 199837 28595 199903 28598
rect 551369 28595 551435 28598
rect 233785 28522 233851 28525
rect 399518 28522 399524 28524
rect 233785 28520 399524 28522
rect 233785 28464 233790 28520
rect 233846 28464 399524 28520
rect 233785 28462 399524 28464
rect 233785 28459 233851 28462
rect 399518 28460 399524 28462
rect 399588 28460 399594 28524
rect 242249 28386 242315 28389
rect 399334 28386 399340 28388
rect 242249 28384 399340 28386
rect 242249 28328 242254 28384
rect 242310 28328 399340 28384
rect 242249 28326 399340 28328
rect 242249 28323 242315 28326
rect 399334 28324 399340 28326
rect 399404 28324 399410 28388
rect 168230 27508 168236 27572
rect 168300 27570 168306 27572
rect 397494 27570 397500 27572
rect 168300 27510 397500 27570
rect 168300 27508 168306 27510
rect 397494 27508 397500 27510
rect 397564 27508 397570 27572
rect 580257 19818 580323 19821
rect 583520 19818 584960 19908
rect 580257 19816 584960 19818
rect 580257 19760 580262 19816
rect 580318 19760 584960 19816
rect 580257 19758 584960 19760
rect 580257 19755 580323 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6340 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 435772 499700 435836 499764
rect 436046 499700 436110 499764
rect 67220 498204 67284 498268
rect 74212 498204 74276 498268
rect 77708 498204 77772 498268
rect 91876 498204 91940 498268
rect 95924 498204 95988 498268
rect 103284 498204 103348 498268
rect 120948 498204 121012 498268
rect 145972 498204 146036 498268
rect 153332 498204 153396 498268
rect 419580 498204 419644 498268
rect 455644 498204 455708 498268
rect 463556 498204 463620 498268
rect 73108 498068 73172 498132
rect 78812 498068 78876 498132
rect 80100 498068 80164 498132
rect 85804 498068 85868 498132
rect 86172 498068 86236 498132
rect 89484 498128 89548 498132
rect 89484 498072 89534 498128
rect 89534 498072 89548 498128
rect 89484 498068 89548 498072
rect 103652 498068 103716 498132
rect 113404 498068 113468 498132
rect 115980 498068 116044 498132
rect 118372 498068 118436 498132
rect 125916 498068 125980 498132
rect 128492 498068 128556 498132
rect 150940 498128 151004 498132
rect 150940 498072 150990 498128
rect 150990 498072 151004 498128
rect 150940 498068 151004 498072
rect 434484 498068 434548 498132
rect 441108 498068 441172 498132
rect 456196 498068 456260 498132
rect 96292 497856 96356 497860
rect 96292 497800 96342 497856
rect 96342 497800 96356 497856
rect 96292 497796 96356 497800
rect 71820 497388 71884 497452
rect 458036 497252 458100 497316
rect 432276 497116 432340 497180
rect 80836 496980 80900 497044
rect 83412 496980 83476 497044
rect 87092 496980 87156 497044
rect 92796 496980 92860 497044
rect 95188 496980 95252 497044
rect 98316 496980 98380 497044
rect 100892 496980 100956 497044
rect 106044 497040 106108 497044
rect 106044 496984 106094 497040
rect 106094 496984 106108 497040
rect 106044 496980 106108 496984
rect 108068 496980 108132 497044
rect 426572 496980 426636 497044
rect 428228 496980 428292 497044
rect 431172 496980 431236 497044
rect 433564 496980 433628 497044
rect 435956 496980 436020 497044
rect 438532 496980 438596 497044
rect 442764 496980 442828 497044
rect 443868 496980 443932 497044
rect 446260 496980 446324 497044
rect 448284 496980 448348 497044
rect 449756 496980 449820 497044
rect 451044 496980 451108 497044
rect 453620 496980 453684 497044
rect 458956 496980 459020 497044
rect 498516 496980 498580 497044
rect 66116 496904 66180 496908
rect 66116 496848 66166 496904
rect 66166 496848 66180 496904
rect 66116 496844 66180 496848
rect 68324 496844 68388 496908
rect 69612 496844 69676 496908
rect 70532 496844 70596 496908
rect 75500 496844 75564 496908
rect 76604 496844 76668 496908
rect 78260 496904 78324 496908
rect 78260 496848 78310 496904
rect 78310 496848 78324 496904
rect 78260 496844 78324 496848
rect 81020 496844 81084 496908
rect 82492 496844 82556 496908
rect 83596 496844 83660 496908
rect 84516 496844 84580 496908
rect 88196 496904 88260 496908
rect 88196 496848 88246 496904
rect 88246 496848 88260 496904
rect 88196 496844 88260 496848
rect 88564 496844 88628 496908
rect 90772 496844 90836 496908
rect 91140 496904 91204 496908
rect 91140 496848 91190 496904
rect 91190 496848 91204 496904
rect 91140 496844 91204 496848
rect 93532 496844 93596 496908
rect 93900 496844 93964 496908
rect 97580 496844 97644 496908
rect 98684 496844 98748 496908
rect 99972 496844 100036 496908
rect 101260 496844 101324 496908
rect 102180 496844 102244 496908
rect 104388 496844 104452 496908
rect 105860 496844 105924 496908
rect 106964 496844 107028 496908
rect 108436 496844 108500 496908
rect 109172 496844 109236 496908
rect 111012 496844 111076 496908
rect 123524 496844 123588 496908
rect 130884 496844 130948 496908
rect 133460 496844 133524 496908
rect 136036 496844 136100 496908
rect 138612 496844 138676 496908
rect 141004 496844 141068 496908
rect 143396 496904 143460 496908
rect 143396 496848 143446 496904
rect 143446 496848 143460 496904
rect 143396 496844 143460 496848
rect 148548 496844 148612 496908
rect 155908 496844 155972 496908
rect 415532 496844 415596 496908
rect 417188 496844 417252 496908
rect 418292 496844 418356 496908
rect 420500 496844 420564 496908
rect 421788 496844 421852 496908
rect 423076 496844 423140 496908
rect 424180 496844 424244 496908
rect 425468 496844 425532 496908
rect 427676 496844 427740 496908
rect 428596 496844 428660 496908
rect 430068 496844 430132 496908
rect 430804 496844 430868 496908
rect 433380 496904 433444 496908
rect 433380 496848 433394 496904
rect 433394 496848 433444 496904
rect 433380 496844 433444 496848
rect 435772 496844 435836 496908
rect 436876 496844 436940 496908
rect 438348 496844 438412 496908
rect 439452 496844 439516 496908
rect 440556 496844 440620 496908
rect 442028 496844 442092 496908
rect 443500 496844 443564 496908
rect 444788 496844 444852 496908
rect 445892 496904 445956 496908
rect 445892 496848 445942 496904
rect 445942 496848 445956 496904
rect 445892 496844 445956 496848
rect 447548 496844 447612 496908
rect 448652 496844 448716 496908
rect 450860 496844 450924 496908
rect 452516 496844 452580 496908
rect 453252 496844 453316 496908
rect 454356 496844 454420 496908
rect 456932 496904 456996 496908
rect 456932 496848 456946 496904
rect 456946 496848 456996 496904
rect 456932 496844 456996 496848
rect 458404 496844 458468 496908
rect 460980 496904 461044 496908
rect 460980 496848 460994 496904
rect 460994 496848 461044 496904
rect 460980 496844 461044 496848
rect 465948 496844 466012 496908
rect 468156 496844 468220 496908
rect 470916 496844 470980 496908
rect 473308 496904 473372 496908
rect 473308 496848 473358 496904
rect 473358 496848 473372 496904
rect 473308 496844 473372 496848
rect 475884 496844 475948 496908
rect 478460 496844 478524 496908
rect 480668 496844 480732 496908
rect 483428 496844 483492 496908
rect 486004 496844 486068 496908
rect 488580 496904 488644 496908
rect 488580 496848 488594 496904
rect 488594 496848 488644 496904
rect 488580 496844 488644 496848
rect 490972 496844 491036 496908
rect 493364 496844 493428 496908
rect 495940 496844 496004 496908
rect 500908 496904 500972 496908
rect 500908 496848 500958 496904
rect 500958 496848 500972 496904
rect 500908 496844 500972 496848
rect 503300 496844 503364 496908
rect 505508 496844 505572 496908
rect 412772 422316 412836 422380
rect 169156 420956 169220 421020
rect 414612 420956 414676 421020
rect 408540 420140 408604 420204
rect 409828 408852 409892 408916
rect 412956 406676 413020 406740
rect 412404 401916 412468 401980
rect 410012 377300 410076 377364
rect 411300 301684 411364 301748
rect 411484 297604 411548 297668
rect 411668 240076 411732 240140
rect 409460 224980 409524 225044
rect 411852 215324 411916 215388
rect 399524 199548 399588 199612
rect 409092 199548 409156 199612
rect 411852 199412 411916 199476
rect 399340 199276 399404 199340
rect 412772 199276 412836 199340
rect 398604 196556 398668 196620
rect 408540 196012 408604 196076
rect 409828 195332 409892 195396
rect 410012 195196 410076 195260
rect 399708 194108 399772 194172
rect 411484 194108 411548 194172
rect 168236 193972 168300 194036
rect 167316 193836 167380 193900
rect 412956 192476 413020 192540
rect 412404 145556 412468 145620
rect 411668 144060 411732 144124
rect 411300 142700 411364 142764
rect 414612 142700 414676 142764
rect 169340 139980 169404 140044
rect 168052 139844 168116 139908
rect 169524 139844 169588 139908
rect 167684 139436 167748 139500
rect 398052 139436 398116 139500
rect 398788 139436 398852 139500
rect 399708 139436 399772 139500
rect 168052 137532 168116 137596
rect 398604 137532 398668 137596
rect 167868 136580 167932 136644
rect 167684 135900 167748 135964
rect 167684 135628 167748 135692
rect 169156 129372 169220 129436
rect 167868 127740 167932 127804
rect 167316 122844 167380 122908
rect 168236 121212 168300 121276
rect 398788 108020 398852 108084
rect 398052 106388 398116 106452
rect 169524 93196 169588 93260
rect 169340 91564 169404 91628
rect 167684 85036 167748 85100
rect 168236 78508 168300 78572
rect 168052 63684 168116 63748
rect 397868 63412 397932 63476
rect 167684 60420 167748 60484
rect 397684 59196 397748 59260
rect 167868 57156 167932 57220
rect 168236 41440 168300 41444
rect 168236 41384 168286 41440
rect 168286 41384 168300 41440
rect 168236 41380 168300 41384
rect 168236 40700 168300 40764
rect 168972 39884 169036 39948
rect 397500 33084 397564 33148
rect 168052 30636 168116 30700
rect 397868 30636 397932 30700
rect 397500 30228 397564 30292
rect 168972 30092 169036 30156
rect 167868 29956 167932 30020
rect 168236 29820 168300 29884
rect 399524 28460 399588 28524
rect 399340 28324 399404 28388
rect 168236 27508 168300 27572
rect 397500 27508 397564 27572
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 402000 31574 428058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 402000 38414 434898
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 402000 42134 402618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 585308 49574 590058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 585308 56414 596898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 585308 60134 600618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 585308 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 585308 67574 608058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 585308 74414 614898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 585308 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 585308 81854 586338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 585308 85574 590058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 585308 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 585308 96134 600618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 585308 99854 604338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 585308 103574 608058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 585308 110414 614898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 585308 114134 618618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 585308 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 585308 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 585308 128414 596898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 585308 132134 600618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 585308 135854 604338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 585308 139574 608058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 585308 146414 614898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 585308 150134 618618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 585308 153854 586338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 585308 157574 590058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 585308 164414 596898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 585308 168134 600618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 585308 171854 604338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 585308 175574 608058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 585308 182414 614898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 585308 186134 618618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 50952 579454 51300 579486
rect 50952 579218 51008 579454
rect 51244 579218 51300 579454
rect 50952 579134 51300 579218
rect 50952 578898 51008 579134
rect 51244 578898 51300 579134
rect 50952 578866 51300 578898
rect 185320 579454 185668 579486
rect 185320 579218 185376 579454
rect 185612 579218 185668 579454
rect 185320 579134 185668 579218
rect 185320 578898 185376 579134
rect 185612 578898 185668 579134
rect 185320 578866 185668 578898
rect 50272 561454 50620 561486
rect 50272 561218 50328 561454
rect 50564 561218 50620 561454
rect 50272 561134 50620 561218
rect 50272 560898 50328 561134
rect 50564 560898 50620 561134
rect 50272 560866 50620 560898
rect 186000 561454 186348 561486
rect 186000 561218 186056 561454
rect 186292 561218 186348 561454
rect 186000 561134 186348 561218
rect 186000 560898 186056 561134
rect 186292 560898 186348 561134
rect 186000 560866 186348 560898
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 50952 543454 51300 543486
rect 50952 543218 51008 543454
rect 51244 543218 51300 543454
rect 50952 543134 51300 543218
rect 50952 542898 51008 543134
rect 51244 542898 51300 543134
rect 50952 542866 51300 542898
rect 185320 543454 185668 543486
rect 185320 543218 185376 543454
rect 185612 543218 185668 543454
rect 185320 543134 185668 543218
rect 185320 542898 185376 543134
rect 185612 542898 185668 543134
rect 185320 542866 185668 542898
rect 50272 525454 50620 525486
rect 50272 525218 50328 525454
rect 50564 525218 50620 525454
rect 50272 525134 50620 525218
rect 50272 524898 50328 525134
rect 50564 524898 50620 525134
rect 50272 524866 50620 524898
rect 186000 525454 186348 525486
rect 186000 525218 186056 525454
rect 186292 525218 186348 525454
rect 186000 525134 186348 525218
rect 186000 524898 186056 525134
rect 186292 524898 186348 525134
rect 186000 524866 186348 524898
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 50952 507454 51300 507486
rect 50952 507218 51008 507454
rect 51244 507218 51300 507454
rect 50952 507134 51300 507218
rect 50952 506898 51008 507134
rect 51244 506898 51300 507134
rect 50952 506866 51300 506898
rect 185320 507454 185668 507486
rect 185320 507218 185376 507454
rect 185612 507218 185668 507454
rect 185320 507134 185668 507218
rect 185320 506898 185376 507134
rect 185612 506898 185668 507134
rect 185320 506866 185668 506898
rect 66056 499590 66116 500106
rect 67144 499590 67204 500106
rect 68232 499590 68292 500106
rect 69592 499590 69652 500106
rect 70544 499590 70604 500106
rect 66056 499530 66178 499590
rect 67144 499530 67282 499590
rect 68232 499530 68386 499590
rect 69592 499530 69674 499590
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 402000 45854 406338
rect 48954 482614 49574 498000
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 402000 49574 410058
rect 55794 489454 56414 498000
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 402000 56414 416898
rect 59514 493174 60134 498000
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 402000 60134 420618
rect 63234 496894 63854 498000
rect 66118 496909 66178 499530
rect 67222 498269 67282 499530
rect 67219 498268 67285 498269
rect 67219 498204 67220 498268
rect 67284 498204 67285 498268
rect 67219 498203 67285 498204
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 66115 496908 66181 496909
rect 66115 496844 66116 496908
rect 66180 496844 66181 496908
rect 66115 496843 66181 496844
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 402000 63854 424338
rect 66954 464614 67574 498000
rect 68326 496909 68386 499530
rect 69614 496909 69674 499530
rect 70534 499530 70604 499590
rect 71768 499590 71828 500106
rect 73128 499590 73188 500106
rect 74216 499590 74276 500106
rect 71768 499530 71882 499590
rect 70534 496909 70594 499530
rect 71822 497453 71882 499530
rect 73110 499530 73188 499590
rect 74214 499530 74276 499590
rect 75440 499590 75500 500106
rect 76528 499590 76588 500106
rect 77616 499590 77676 500106
rect 78296 499590 78356 500106
rect 75440 499530 75562 499590
rect 76528 499530 76666 499590
rect 77616 499530 77770 499590
rect 73110 498133 73170 499530
rect 74214 498269 74274 499530
rect 74211 498268 74277 498269
rect 74211 498204 74212 498268
rect 74276 498204 74277 498268
rect 74211 498203 74277 498204
rect 73107 498132 73173 498133
rect 73107 498068 73108 498132
rect 73172 498068 73173 498132
rect 73107 498067 73173 498068
rect 71819 497452 71885 497453
rect 71819 497388 71820 497452
rect 71884 497388 71885 497452
rect 71819 497387 71885 497388
rect 68323 496908 68389 496909
rect 68323 496844 68324 496908
rect 68388 496844 68389 496908
rect 68323 496843 68389 496844
rect 69611 496908 69677 496909
rect 69611 496844 69612 496908
rect 69676 496844 69677 496908
rect 69611 496843 69677 496844
rect 70531 496908 70597 496909
rect 70531 496844 70532 496908
rect 70596 496844 70597 496908
rect 70531 496843 70597 496844
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 428614 67574 464058
rect 66954 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 67574 428614
rect 66954 428294 67574 428378
rect 66954 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 67574 428294
rect 66954 402000 67574 428058
rect 73794 471454 74414 498000
rect 75502 496909 75562 499530
rect 76606 496909 76666 499530
rect 77710 498269 77770 499530
rect 78262 499530 78356 499590
rect 78704 499590 78764 500106
rect 80064 499590 80124 500106
rect 80744 499590 80804 500106
rect 81288 499590 81348 500106
rect 78704 499530 78874 499590
rect 80064 499530 80162 499590
rect 80744 499530 80898 499590
rect 77707 498268 77773 498269
rect 77707 498204 77708 498268
rect 77772 498204 77773 498268
rect 77707 498203 77773 498204
rect 75499 496908 75565 496909
rect 75499 496844 75500 496908
rect 75564 496844 75565 496908
rect 75499 496843 75565 496844
rect 76603 496908 76669 496909
rect 76603 496844 76604 496908
rect 76668 496844 76669 496908
rect 76603 496843 76669 496844
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 73794 402000 74414 434898
rect 77514 475174 78134 498000
rect 78262 496909 78322 499530
rect 78814 498133 78874 499530
rect 80102 498133 80162 499530
rect 78811 498132 78877 498133
rect 78811 498068 78812 498132
rect 78876 498068 78877 498132
rect 78811 498067 78877 498068
rect 80099 498132 80165 498133
rect 80099 498068 80100 498132
rect 80164 498068 80165 498132
rect 80099 498067 80165 498068
rect 80838 497045 80898 499530
rect 81022 499530 81348 499590
rect 82376 499590 82436 500106
rect 83464 499590 83524 500106
rect 83600 499590 83660 500106
rect 84552 499590 84612 500106
rect 85912 499590 85972 500106
rect 82376 499530 82554 499590
rect 80835 497044 80901 497045
rect 80835 496980 80836 497044
rect 80900 496980 80901 497044
rect 80835 496979 80901 496980
rect 81022 496909 81082 499530
rect 78259 496908 78325 496909
rect 78259 496844 78260 496908
rect 78324 496844 78325 496908
rect 78259 496843 78325 496844
rect 81019 496908 81085 496909
rect 81019 496844 81020 496908
rect 81084 496844 81085 496908
rect 81019 496843 81085 496844
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 402000 78134 402618
rect 81234 478894 81854 498000
rect 82494 496909 82554 499530
rect 83414 499530 83524 499590
rect 83598 499530 83660 499590
rect 84518 499530 84612 499590
rect 85806 499530 85972 499590
rect 86048 499590 86108 500106
rect 87000 499590 87060 500106
rect 88088 499590 88148 500106
rect 88496 499590 88556 500106
rect 89448 499590 89508 500106
rect 90672 499590 90732 500106
rect 91080 499590 91140 500106
rect 91760 499590 91820 500106
rect 92848 499590 92908 500106
rect 86048 499530 86234 499590
rect 87000 499530 87154 499590
rect 88088 499530 88258 499590
rect 88496 499530 88626 499590
rect 89448 499530 89546 499590
rect 90672 499530 90834 499590
rect 91080 499530 91202 499590
rect 91760 499530 91938 499590
rect 83414 497045 83474 499530
rect 83411 497044 83477 497045
rect 83411 496980 83412 497044
rect 83476 496980 83477 497044
rect 83411 496979 83477 496980
rect 83598 496909 83658 499530
rect 84518 496909 84578 499530
rect 85806 498133 85866 499530
rect 86174 498133 86234 499530
rect 85803 498132 85869 498133
rect 85803 498068 85804 498132
rect 85868 498068 85869 498132
rect 85803 498067 85869 498068
rect 86171 498132 86237 498133
rect 86171 498068 86172 498132
rect 86236 498068 86237 498132
rect 86171 498067 86237 498068
rect 82491 496908 82557 496909
rect 82491 496844 82492 496908
rect 82556 496844 82557 496908
rect 82491 496843 82557 496844
rect 83595 496908 83661 496909
rect 83595 496844 83596 496908
rect 83660 496844 83661 496908
rect 83595 496843 83661 496844
rect 84515 496908 84581 496909
rect 84515 496844 84516 496908
rect 84580 496844 84581 496908
rect 84515 496843 84581 496844
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 81234 402000 81854 406338
rect 84954 482614 85574 498000
rect 87094 497045 87154 499530
rect 87091 497044 87157 497045
rect 87091 496980 87092 497044
rect 87156 496980 87157 497044
rect 87091 496979 87157 496980
rect 88198 496909 88258 499530
rect 88566 496909 88626 499530
rect 89486 498133 89546 499530
rect 89483 498132 89549 498133
rect 89483 498068 89484 498132
rect 89548 498068 89549 498132
rect 89483 498067 89549 498068
rect 90774 496909 90834 499530
rect 91142 496909 91202 499530
rect 91878 498269 91938 499530
rect 92798 499530 92908 499590
rect 93528 499590 93588 500106
rect 93936 499590 93996 500106
rect 95296 499590 95356 500106
rect 95976 499590 96036 500106
rect 96384 499590 96444 500106
rect 97608 499590 97668 500106
rect 93528 499530 93594 499590
rect 91875 498268 91941 498269
rect 91875 498204 91876 498268
rect 91940 498204 91941 498268
rect 91875 498203 91941 498204
rect 88195 496908 88261 496909
rect 88195 496844 88196 496908
rect 88260 496844 88261 496908
rect 88195 496843 88261 496844
rect 88563 496908 88629 496909
rect 88563 496844 88564 496908
rect 88628 496844 88629 496908
rect 88563 496843 88629 496844
rect 90771 496908 90837 496909
rect 90771 496844 90772 496908
rect 90836 496844 90837 496908
rect 90771 496843 90837 496844
rect 91139 496908 91205 496909
rect 91139 496844 91140 496908
rect 91204 496844 91205 496908
rect 91139 496843 91205 496844
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 402000 85574 410058
rect 91794 489454 92414 498000
rect 92798 497045 92858 499530
rect 92795 497044 92861 497045
rect 92795 496980 92796 497044
rect 92860 496980 92861 497044
rect 92795 496979 92861 496980
rect 93534 496909 93594 499530
rect 93902 499530 93996 499590
rect 95190 499530 95356 499590
rect 95926 499530 96036 499590
rect 96294 499530 96444 499590
rect 97582 499530 97668 499590
rect 98288 499590 98348 500106
rect 98696 499590 98756 500106
rect 98288 499530 98378 499590
rect 93902 496909 93962 499530
rect 95190 497045 95250 499530
rect 95926 498269 95986 499530
rect 95923 498268 95989 498269
rect 95923 498204 95924 498268
rect 95988 498204 95989 498268
rect 95923 498203 95989 498204
rect 95187 497044 95253 497045
rect 95187 496980 95188 497044
rect 95252 496980 95253 497044
rect 95187 496979 95253 496980
rect 93531 496908 93597 496909
rect 93531 496844 93532 496908
rect 93596 496844 93597 496908
rect 93531 496843 93597 496844
rect 93899 496908 93965 496909
rect 93899 496844 93900 496908
rect 93964 496844 93965 496908
rect 93899 496843 93965 496844
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 453454 92414 488898
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 417454 92414 452898
rect 91794 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 92414 417454
rect 91794 417134 92414 417218
rect 91794 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 92414 417134
rect 91794 402000 92414 416898
rect 95514 493174 96134 498000
rect 96294 497861 96354 499530
rect 96291 497860 96357 497861
rect 96291 497796 96292 497860
rect 96356 497796 96357 497860
rect 96291 497795 96357 497796
rect 97582 496909 97642 499530
rect 98318 497045 98378 499530
rect 98686 499530 98756 499590
rect 99784 499590 99844 500106
rect 101008 499590 101068 500106
rect 99784 499530 100034 499590
rect 98315 497044 98381 497045
rect 98315 496980 98316 497044
rect 98380 496980 98381 497044
rect 98315 496979 98381 496980
rect 98686 496909 98746 499530
rect 97579 496908 97645 496909
rect 97579 496844 97580 496908
rect 97644 496844 97645 496908
rect 97579 496843 97645 496844
rect 98683 496908 98749 496909
rect 98683 496844 98684 496908
rect 98748 496844 98749 496908
rect 98683 496843 98749 496844
rect 99234 496894 99854 498000
rect 99974 496909 100034 499530
rect 100894 499530 101068 499590
rect 101144 499590 101204 500106
rect 102232 499590 102292 500106
rect 103320 499590 103380 500106
rect 101144 499530 101322 499590
rect 100894 497045 100954 499530
rect 100891 497044 100957 497045
rect 100891 496980 100892 497044
rect 100956 496980 100957 497044
rect 100891 496979 100957 496980
rect 101262 496909 101322 499530
rect 102182 499530 102292 499590
rect 103286 499530 103380 499590
rect 103592 499590 103652 500106
rect 104408 499590 104468 500106
rect 103592 499530 103714 499590
rect 102182 496909 102242 499530
rect 103286 498269 103346 499530
rect 103283 498268 103349 498269
rect 103283 498204 103284 498268
rect 103348 498204 103349 498268
rect 103283 498203 103349 498204
rect 103654 498133 103714 499530
rect 104390 499530 104468 499590
rect 105768 499590 105828 500106
rect 106040 499590 106100 500106
rect 106992 499590 107052 500106
rect 108080 499590 108140 500106
rect 108488 499590 108548 500106
rect 105768 499530 105922 499590
rect 106040 499530 106106 499590
rect 103651 498132 103717 498133
rect 103651 498068 103652 498132
rect 103716 498068 103717 498132
rect 103651 498067 103717 498068
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95514 421174 96134 456618
rect 95514 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 96134 421174
rect 95514 420854 96134 420938
rect 95514 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 96134 420854
rect 95514 402000 96134 420618
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99971 496908 100037 496909
rect 99971 496844 99972 496908
rect 100036 496844 100037 496908
rect 99971 496843 100037 496844
rect 101259 496908 101325 496909
rect 101259 496844 101260 496908
rect 101324 496844 101325 496908
rect 101259 496843 101325 496844
rect 102179 496908 102245 496909
rect 102179 496844 102180 496908
rect 102244 496844 102245 496908
rect 102179 496843 102245 496844
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 424894 99854 460338
rect 99234 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 99854 424894
rect 99234 424574 99854 424658
rect 99234 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 99854 424574
rect 99234 402000 99854 424338
rect 102954 464614 103574 498000
rect 104390 496909 104450 499530
rect 105862 496909 105922 499530
rect 106046 497045 106106 499530
rect 106966 499530 107052 499590
rect 108070 499530 108140 499590
rect 108438 499530 108548 499590
rect 109168 499590 109228 500106
rect 110936 499590 110996 500106
rect 113520 499590 113580 500106
rect 109168 499530 109234 499590
rect 110936 499530 111074 499590
rect 106043 497044 106109 497045
rect 106043 496980 106044 497044
rect 106108 496980 106109 497044
rect 106043 496979 106109 496980
rect 106966 496909 107026 499530
rect 108070 497045 108130 499530
rect 108067 497044 108133 497045
rect 108067 496980 108068 497044
rect 108132 496980 108133 497044
rect 108067 496979 108133 496980
rect 108438 496909 108498 499530
rect 109174 496909 109234 499530
rect 104387 496908 104453 496909
rect 104387 496844 104388 496908
rect 104452 496844 104453 496908
rect 104387 496843 104453 496844
rect 105859 496908 105925 496909
rect 105859 496844 105860 496908
rect 105924 496844 105925 496908
rect 105859 496843 105925 496844
rect 106963 496908 107029 496909
rect 106963 496844 106964 496908
rect 107028 496844 107029 496908
rect 106963 496843 107029 496844
rect 108435 496908 108501 496909
rect 108435 496844 108436 496908
rect 108500 496844 108501 496908
rect 108435 496843 108501 496844
rect 109171 496908 109237 496909
rect 109171 496844 109172 496908
rect 109236 496844 109237 496908
rect 109171 496843 109237 496844
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 428614 103574 464058
rect 102954 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 103574 428614
rect 102954 428294 103574 428378
rect 102954 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 103574 428294
rect 102954 402000 103574 428058
rect 109794 471454 110414 498000
rect 111014 496909 111074 499530
rect 113406 499530 113580 499590
rect 115968 499590 116028 500106
rect 118280 499590 118340 500106
rect 121000 499590 121060 500106
rect 115968 499530 116042 499590
rect 118280 499530 118434 499590
rect 113406 498133 113466 499530
rect 115982 498133 116042 499530
rect 118374 498133 118434 499530
rect 120950 499530 121060 499590
rect 123448 499590 123508 500106
rect 125896 499590 125956 500106
rect 128480 499590 128540 500106
rect 130928 499590 130988 500106
rect 133512 499590 133572 500106
rect 123448 499530 123586 499590
rect 125896 499530 125978 499590
rect 128480 499530 128554 499590
rect 120950 498269 121010 499530
rect 120947 498268 121013 498269
rect 120947 498204 120948 498268
rect 121012 498204 121013 498268
rect 120947 498203 121013 498204
rect 113403 498132 113469 498133
rect 113403 498068 113404 498132
rect 113468 498068 113469 498132
rect 113403 498067 113469 498068
rect 115979 498132 116045 498133
rect 115979 498068 115980 498132
rect 116044 498068 116045 498132
rect 115979 498067 116045 498068
rect 118371 498132 118437 498133
rect 118371 498068 118372 498132
rect 118436 498068 118437 498132
rect 118371 498067 118437 498068
rect 111011 496908 111077 496909
rect 111011 496844 111012 496908
rect 111076 496844 111077 496908
rect 111011 496843 111077 496844
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 435454 110414 470898
rect 109794 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 110414 435454
rect 109794 435134 110414 435218
rect 109794 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 110414 435134
rect 109794 402000 110414 434898
rect 113514 475174 114134 498000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 113514 402000 114134 402618
rect 117234 478894 117854 498000
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 402000 117854 406338
rect 120954 482614 121574 498000
rect 123526 496909 123586 499530
rect 125918 498133 125978 499530
rect 128494 498133 128554 499530
rect 130886 499530 130988 499590
rect 133462 499530 133572 499590
rect 135960 499590 136020 500106
rect 138544 499590 138604 500106
rect 140992 499590 141052 500106
rect 143440 499590 143500 500106
rect 135960 499530 136098 499590
rect 138544 499530 138674 499590
rect 140992 499530 141066 499590
rect 125915 498132 125981 498133
rect 125915 498068 125916 498132
rect 125980 498068 125981 498132
rect 125915 498067 125981 498068
rect 128491 498132 128557 498133
rect 128491 498068 128492 498132
rect 128556 498068 128557 498132
rect 128491 498067 128557 498068
rect 123523 496908 123589 496909
rect 123523 496844 123524 496908
rect 123588 496844 123589 496908
rect 123523 496843 123589 496844
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 402000 121574 410058
rect 127794 489454 128414 498000
rect 130886 496909 130946 499530
rect 130883 496908 130949 496909
rect 130883 496844 130884 496908
rect 130948 496844 130949 496908
rect 130883 496843 130949 496844
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 402000 128414 416898
rect 131514 493174 132134 498000
rect 133462 496909 133522 499530
rect 133459 496908 133525 496909
rect 133459 496844 133460 496908
rect 133524 496844 133525 496908
rect 133459 496843 133525 496844
rect 135234 496894 135854 498000
rect 136038 496909 136098 499530
rect 138614 496909 138674 499530
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 402000 132134 420618
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 136035 496908 136101 496909
rect 136035 496844 136036 496908
rect 136100 496844 136101 496908
rect 136035 496843 136101 496844
rect 138611 496908 138677 496909
rect 138611 496844 138612 496908
rect 138676 496844 138677 496908
rect 138611 496843 138677 496844
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 49568 381454 49888 381486
rect 49568 381218 49610 381454
rect 49846 381218 49888 381454
rect 49568 381134 49888 381218
rect 49568 380898 49610 381134
rect 49846 380898 49888 381134
rect 49568 380866 49888 380898
rect 80288 381454 80608 381486
rect 80288 381218 80330 381454
rect 80566 381218 80608 381454
rect 80288 381134 80608 381218
rect 80288 380898 80330 381134
rect 80566 380898 80608 381134
rect 80288 380866 80608 380898
rect 111008 381454 111328 381486
rect 111008 381218 111050 381454
rect 111286 381218 111328 381454
rect 111008 381134 111328 381218
rect 111008 380898 111050 381134
rect 111286 380898 111328 381134
rect 111008 380866 111328 380898
rect 34208 363454 34528 363486
rect 34208 363218 34250 363454
rect 34486 363218 34528 363454
rect 34208 363134 34528 363218
rect 34208 362898 34250 363134
rect 34486 362898 34528 363134
rect 34208 362866 34528 362898
rect 64928 363454 65248 363486
rect 64928 363218 64970 363454
rect 65206 363218 65248 363454
rect 64928 363134 65248 363218
rect 64928 362898 64970 363134
rect 65206 362898 65248 363134
rect 64928 362866 65248 362898
rect 95648 363454 95968 363486
rect 95648 363218 95690 363454
rect 95926 363218 95968 363454
rect 95648 363134 95968 363218
rect 95648 362898 95690 363134
rect 95926 362898 95968 363134
rect 95648 362866 95968 362898
rect 126368 363454 126688 363486
rect 126368 363218 126410 363454
rect 126646 363218 126688 363454
rect 126368 363134 126688 363218
rect 126368 362898 126410 363134
rect 126646 362898 126688 363134
rect 126368 362866 126688 362898
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 49568 345454 49888 345486
rect 49568 345218 49610 345454
rect 49846 345218 49888 345454
rect 49568 345134 49888 345218
rect 49568 344898 49610 345134
rect 49846 344898 49888 345134
rect 49568 344866 49888 344898
rect 80288 345454 80608 345486
rect 80288 345218 80330 345454
rect 80566 345218 80608 345454
rect 80288 345134 80608 345218
rect 80288 344898 80330 345134
rect 80566 344898 80608 345134
rect 80288 344866 80608 344898
rect 111008 345454 111328 345486
rect 111008 345218 111050 345454
rect 111286 345218 111328 345454
rect 111008 345134 111328 345218
rect 111008 344898 111050 345134
rect 111286 344898 111328 345134
rect 111008 344866 111328 344898
rect 34208 327454 34528 327486
rect 34208 327218 34250 327454
rect 34486 327218 34528 327454
rect 34208 327134 34528 327218
rect 34208 326898 34250 327134
rect 34486 326898 34528 327134
rect 34208 326866 34528 326898
rect 64928 327454 65248 327486
rect 64928 327218 64970 327454
rect 65206 327218 65248 327454
rect 64928 327134 65248 327218
rect 64928 326898 64970 327134
rect 65206 326898 65248 327134
rect 64928 326866 65248 326898
rect 95648 327454 95968 327486
rect 95648 327218 95690 327454
rect 95926 327218 95968 327454
rect 95648 327134 95968 327218
rect 95648 326898 95690 327134
rect 95926 326898 95968 327134
rect 95648 326866 95968 326898
rect 126368 327454 126688 327486
rect 126368 327218 126410 327454
rect 126646 327218 126688 327454
rect 126368 327134 126688 327218
rect 126368 326898 126410 327134
rect 126646 326898 126688 327134
rect 126368 326866 126688 326898
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 49568 309454 49888 309486
rect 49568 309218 49610 309454
rect 49846 309218 49888 309454
rect 49568 309134 49888 309218
rect 49568 308898 49610 309134
rect 49846 308898 49888 309134
rect 49568 308866 49888 308898
rect 80288 309454 80608 309486
rect 80288 309218 80330 309454
rect 80566 309218 80608 309454
rect 80288 309134 80608 309218
rect 80288 308898 80330 309134
rect 80566 308898 80608 309134
rect 80288 308866 80608 308898
rect 111008 309454 111328 309486
rect 111008 309218 111050 309454
rect 111286 309218 111328 309454
rect 111008 309134 111328 309218
rect 111008 308898 111050 309134
rect 111286 308898 111328 309134
rect 111008 308866 111328 308898
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 284614 31574 298000
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 291454 38414 298000
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 295174 42134 298000
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 262894 45854 298000
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 266614 49574 298000
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 273454 56414 298000
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 277174 60134 298000
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 280894 63854 298000
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 284614 67574 298000
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 212614 67574 248058
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66954 176614 67574 212058
rect 66954 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 67574 176614
rect 66954 176294 67574 176378
rect 66954 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 67574 176294
rect 66954 140614 67574 176058
rect 66954 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 67574 140614
rect 66954 140294 67574 140378
rect 66954 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 67574 140294
rect 66954 104614 67574 140058
rect 66954 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 67574 104614
rect 66954 104294 67574 104378
rect 66954 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 67574 104294
rect 66954 68614 67574 104058
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 291454 74414 298000
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 219454 74414 254898
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 147454 74414 182898
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 111454 74414 146898
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 73794 75454 74414 110898
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 295174 78134 298000
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 223174 78134 258618
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 151174 78134 186618
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 115174 78134 150618
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 262894 81854 298000
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 226894 81854 262338
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 154894 81854 190338
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 118894 81854 154338
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 266614 85574 298000
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 158614 85574 194058
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 122614 85574 158058
rect 84954 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 85574 122614
rect 84954 122294 85574 122378
rect 84954 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 85574 122294
rect 84954 86614 85574 122058
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 273454 92414 298000
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 165454 92414 200898
rect 91794 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 92414 165454
rect 91794 165134 92414 165218
rect 91794 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 92414 165134
rect 91794 129454 92414 164898
rect 91794 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 92414 129454
rect 91794 129134 92414 129218
rect 91794 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 92414 129134
rect 91794 93454 92414 128898
rect 91794 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 92414 93454
rect 91794 93134 92414 93218
rect 91794 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 92414 93134
rect 91794 57454 92414 92898
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 277174 96134 298000
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 205174 96134 240618
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 169174 96134 204618
rect 95514 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 96134 169174
rect 95514 168854 96134 168938
rect 95514 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 96134 168854
rect 95514 133174 96134 168618
rect 95514 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 96134 133174
rect 95514 132854 96134 132938
rect 95514 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 96134 132854
rect 95514 97174 96134 132618
rect 95514 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 96134 97174
rect 95514 96854 96134 96938
rect 95514 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 96134 96854
rect 95514 61174 96134 96618
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 280894 99854 298000
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 208894 99854 244338
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 99234 172894 99854 208338
rect 99234 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 99854 172894
rect 99234 172574 99854 172658
rect 99234 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 99854 172574
rect 99234 136894 99854 172338
rect 99234 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 99854 136894
rect 99234 136574 99854 136658
rect 99234 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 99854 136574
rect 99234 100894 99854 136338
rect 99234 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 99854 100894
rect 99234 100574 99854 100658
rect 99234 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 99854 100574
rect 99234 64894 99854 100338
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 284614 103574 298000
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 212614 103574 248058
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 102954 176614 103574 212058
rect 102954 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 103574 176614
rect 102954 176294 103574 176378
rect 102954 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 103574 176294
rect 102954 140614 103574 176058
rect 102954 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 103574 140614
rect 102954 140294 103574 140378
rect 102954 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 103574 140294
rect 102954 104614 103574 140058
rect 102954 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 103574 104614
rect 102954 104294 103574 104378
rect 102954 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 103574 104294
rect 102954 68614 103574 104058
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 291454 110414 298000
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 219454 110414 254898
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109794 147454 110414 182898
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 111454 110414 146898
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 295174 114134 298000
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 151174 114134 186618
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 115174 114134 150618
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 262894 117854 298000
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 266614 121574 298000
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 273454 128414 298000
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 127794 165454 128414 200898
rect 127794 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 128414 165454
rect 127794 165134 128414 165218
rect 127794 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 128414 165134
rect 127794 129454 128414 164898
rect 127794 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 128414 129454
rect 127794 129134 128414 129218
rect 127794 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 128414 129134
rect 127794 93454 128414 128898
rect 127794 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 128414 93454
rect 127794 93134 128414 93218
rect 127794 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 128414 93134
rect 127794 57454 128414 92898
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 277174 132134 298000
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 205174 132134 240618
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 131514 169174 132134 204618
rect 131514 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 132134 169174
rect 131514 168854 132134 168938
rect 131514 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 132134 168854
rect 131514 133174 132134 168618
rect 131514 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 132134 133174
rect 131514 132854 132134 132938
rect 131514 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 132134 132854
rect 131514 97174 132134 132618
rect 131514 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 132134 97174
rect 131514 96854 132134 96938
rect 131514 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 132134 96854
rect 131514 61174 132134 96618
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 208894 135854 244338
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 135234 172894 135854 208338
rect 135234 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 135854 172894
rect 135234 172574 135854 172658
rect 135234 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 135854 172574
rect 135234 136894 135854 172338
rect 135234 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 135854 136894
rect 135234 136574 135854 136658
rect 135234 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 135854 136574
rect 135234 100894 135854 136338
rect 135234 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 135854 100894
rect 135234 100574 135854 100658
rect 135234 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 135854 100574
rect 135234 64894 135854 100338
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 464614 139574 498000
rect 141006 496909 141066 499530
rect 143398 499530 143500 499590
rect 145888 499590 145948 500106
rect 148472 499590 148532 500106
rect 150920 499590 150980 500106
rect 153368 499590 153428 500106
rect 155952 499590 156012 500106
rect 145888 499530 146034 499590
rect 148472 499530 148610 499590
rect 150920 499530 151002 499590
rect 143398 496909 143458 499530
rect 145974 498269 146034 499530
rect 145971 498268 146037 498269
rect 145971 498204 145972 498268
rect 146036 498204 146037 498268
rect 145971 498203 146037 498204
rect 141003 496908 141069 496909
rect 141003 496844 141004 496908
rect 141068 496844 141069 496908
rect 141003 496843 141069 496844
rect 143395 496908 143461 496909
rect 143395 496844 143396 496908
rect 143460 496844 143461 496908
rect 143395 496843 143461 496844
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 212614 139574 248058
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 138954 176614 139574 212058
rect 138954 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 139574 176614
rect 138954 176294 139574 176378
rect 138954 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 139574 176294
rect 138954 140614 139574 176058
rect 138954 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 139574 140614
rect 138954 140294 139574 140378
rect 138954 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 139574 140294
rect 138954 104614 139574 140058
rect 138954 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 139574 104614
rect 138954 104294 139574 104378
rect 138954 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 139574 104294
rect 138954 68614 139574 104058
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 471454 146414 498000
rect 148550 496909 148610 499530
rect 150942 498133 151002 499530
rect 153334 499530 153428 499590
rect 155910 499530 156012 499590
rect 153334 498269 153394 499530
rect 153331 498268 153397 498269
rect 153331 498204 153332 498268
rect 153396 498204 153397 498268
rect 153331 498203 153397 498204
rect 150939 498132 151005 498133
rect 150939 498068 150940 498132
rect 151004 498068 151005 498132
rect 150939 498067 151005 498068
rect 148547 496908 148613 496909
rect 148547 496844 148548 496908
rect 148612 496844 148613 496908
rect 148547 496843 148613 496844
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 475174 150134 498000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 478894 153854 498000
rect 155910 496909 155970 499530
rect 155907 496908 155973 496909
rect 155907 496844 155908 496908
rect 155972 496844 155973 496908
rect 155907 496843 155973 496844
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 482614 157574 498000
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 489454 164414 498000
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 163794 165454 164414 200898
rect 167514 493174 168134 498000
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 171234 496894 171854 498000
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 169155 421020 169221 421021
rect 169155 420956 169156 421020
rect 169220 420956 169221 421020
rect 169155 420955 169221 420956
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167315 193900 167381 193901
rect 167315 193836 167316 193900
rect 167380 193836 167381 193900
rect 167315 193835 167381 193836
rect 163794 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 164414 165454
rect 163794 165134 164414 165218
rect 163794 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 164414 165134
rect 163794 129454 164414 164898
rect 163794 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 164414 129454
rect 163794 129134 164414 129218
rect 163794 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 164414 129134
rect 163794 93454 164414 128898
rect 167318 122909 167378 193835
rect 167514 169174 168134 204618
rect 168235 194036 168301 194037
rect 168235 193972 168236 194036
rect 168300 193972 168301 194036
rect 168235 193971 168301 193972
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 142000 168134 168618
rect 168051 139908 168117 139909
rect 168051 139844 168052 139908
rect 168116 139844 168117 139908
rect 168051 139843 168117 139844
rect 167683 139500 167749 139501
rect 167683 139436 167684 139500
rect 167748 139436 167749 139500
rect 167683 139435 167749 139436
rect 167686 135965 167746 139435
rect 168054 137597 168114 139843
rect 168051 137596 168117 137597
rect 168051 137532 168052 137596
rect 168116 137532 168117 137596
rect 168051 137531 168117 137532
rect 167867 136644 167933 136645
rect 167867 136580 167868 136644
rect 167932 136580 167933 136644
rect 167867 136579 167933 136580
rect 167683 135964 167749 135965
rect 167683 135900 167684 135964
rect 167748 135900 167749 135964
rect 167683 135899 167749 135900
rect 167683 135692 167749 135693
rect 167683 135628 167684 135692
rect 167748 135628 167749 135692
rect 167683 135627 167749 135628
rect 167315 122908 167381 122909
rect 167315 122844 167316 122908
rect 167380 122844 167381 122908
rect 167315 122843 167381 122844
rect 163794 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 164414 93454
rect 163794 93134 164414 93218
rect 163794 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 164414 93134
rect 163794 57454 164414 92898
rect 167686 85101 167746 135627
rect 167870 127805 167930 136579
rect 167867 127804 167933 127805
rect 167867 127740 167868 127804
rect 167932 127740 167933 127804
rect 167867 127739 167933 127740
rect 168238 121277 168298 193971
rect 169158 129437 169218 420955
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 142000 171854 172338
rect 174954 464614 175574 498000
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 142000 175574 176058
rect 181794 471454 182414 498000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 142000 182414 146898
rect 185514 475174 186134 498000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 422000 189854 442338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 422000 193574 446058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 422000 200414 452898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 422000 204134 456618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 422000 207854 424338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 422000 211574 428058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 422000 218414 434898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 422000 222134 438618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 422000 225854 442338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 422000 229574 446058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 422000 236414 452898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 422000 240134 456618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 422000 243854 424338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 422000 247574 428058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 422000 254414 434898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 422000 258134 438618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 422000 261854 442338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 422000 265574 446058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 422000 272414 452898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 422000 276134 456618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 422000 279854 424338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 422000 283574 428058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 422000 290414 434898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 422000 294134 438618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 422000 297854 442338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 422000 301574 446058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 422000 308414 452898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 422000 312134 456618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 422000 315854 424338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 422000 319574 428058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 422000 326414 434898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 422000 330134 438618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 422000 333854 442338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 422000 337574 446058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 422000 344414 452898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 422000 348134 456618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 422000 351854 424338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 422000 355574 428058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 422000 362414 434898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 422000 366134 438618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 422000 369854 442338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 422000 373574 446058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 422000 380414 452898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 422000 384134 456618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 422000 387854 424338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 585308 398414 614898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 585308 402134 618618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 585308 405854 586338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 585308 409574 590058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 585308 416414 596898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 585308 420134 600618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 585308 423854 604338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 585308 427574 608058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 585308 434414 614898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 585308 438134 618618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 585308 441854 586338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 585308 445574 590058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 585308 452414 596898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 585308 456134 600618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 585308 459854 604338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 585308 463574 608058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 585308 470414 614898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 585308 474134 618618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 585308 477854 586338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 585308 481574 590058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 585308 488414 596898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 585308 492134 600618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 585308 495854 604338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 585308 499574 608058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 585308 506414 614898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 585308 510134 618618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 585308 513854 586338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 585308 517574 590058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 585308 524414 596898
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 585308 528134 600618
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 585308 531854 604338
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 585308 535574 608058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 400952 579454 401300 579486
rect 400952 579218 401008 579454
rect 401244 579218 401300 579454
rect 400952 579134 401300 579218
rect 400952 578898 401008 579134
rect 401244 578898 401300 579134
rect 400952 578866 401300 578898
rect 535320 579454 535668 579486
rect 535320 579218 535376 579454
rect 535612 579218 535668 579454
rect 535320 579134 535668 579218
rect 535320 578898 535376 579134
rect 535612 578898 535668 579134
rect 535320 578866 535668 578898
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 400272 561454 400620 561486
rect 400272 561218 400328 561454
rect 400564 561218 400620 561454
rect 400272 561134 400620 561218
rect 400272 560898 400328 561134
rect 400564 560898 400620 561134
rect 400272 560866 400620 560898
rect 536000 561454 536348 561486
rect 536000 561218 536056 561454
rect 536292 561218 536348 561454
rect 536000 561134 536348 561218
rect 536000 560898 536056 561134
rect 536292 560898 536348 561134
rect 536000 560866 536348 560898
rect 400952 543454 401300 543486
rect 400952 543218 401008 543454
rect 401244 543218 401300 543454
rect 400952 543134 401300 543218
rect 400952 542898 401008 543134
rect 401244 542898 401300 543134
rect 400952 542866 401300 542898
rect 535320 543454 535668 543486
rect 535320 543218 535376 543454
rect 535612 543218 535668 543454
rect 535320 543134 535668 543218
rect 535320 542898 535376 543134
rect 535612 542898 535668 543134
rect 535320 542866 535668 542898
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 400272 525454 400620 525486
rect 400272 525218 400328 525454
rect 400564 525218 400620 525454
rect 400272 525134 400620 525218
rect 400272 524898 400328 525134
rect 400564 524898 400620 525134
rect 400272 524866 400620 524898
rect 536000 525454 536348 525486
rect 536000 525218 536056 525454
rect 536292 525218 536348 525454
rect 536000 525134 536348 525218
rect 536000 524898 536056 525134
rect 536292 524898 536348 525134
rect 536000 524866 536348 524898
rect 400952 507454 401300 507486
rect 400952 507218 401008 507454
rect 401244 507218 401300 507454
rect 400952 507134 401300 507218
rect 400952 506898 401008 507134
rect 401244 506898 401300 507134
rect 400952 506866 401300 506898
rect 535320 507454 535668 507486
rect 535320 507218 535376 507454
rect 535612 507218 535668 507454
rect 535320 507134 535668 507218
rect 535320 506898 535376 507134
rect 535612 506898 535668 507134
rect 535320 506866 535668 506898
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 416056 499590 416116 500106
rect 415534 499530 416116 499590
rect 417144 499590 417204 500106
rect 418232 499590 418292 500106
rect 419592 499590 419652 500106
rect 420544 499590 420604 500106
rect 417144 499530 417250 499590
rect 418232 499530 418354 499590
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 422000 391574 428058
rect 397794 471454 398414 498000
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 422000 398414 434898
rect 401514 475174 402134 498000
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 422000 402134 438618
rect 405234 478894 405854 498000
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 422000 405854 442338
rect 408954 482614 409574 498000
rect 415534 496909 415594 499530
rect 415531 496908 415597 496909
rect 415531 496844 415532 496908
rect 415596 496844 415597 496908
rect 415531 496843 415597 496844
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 422000 409574 446058
rect 415794 489454 416414 498000
rect 417190 496909 417250 499530
rect 418294 496909 418354 499530
rect 419582 499530 419652 499590
rect 420502 499530 420604 499590
rect 421768 499590 421828 500106
rect 423128 499590 423188 500106
rect 424216 499590 424276 500106
rect 421768 499530 421850 499590
rect 419582 498269 419642 499530
rect 419579 498268 419645 498269
rect 419579 498204 419580 498268
rect 419644 498204 419645 498268
rect 419579 498203 419645 498204
rect 417187 496908 417253 496909
rect 417187 496844 417188 496908
rect 417252 496844 417253 496908
rect 417187 496843 417253 496844
rect 418291 496908 418357 496909
rect 418291 496844 418292 496908
rect 418356 496844 418357 496908
rect 418291 496843 418357 496844
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 412771 422380 412837 422381
rect 412771 422316 412772 422380
rect 412836 422316 412837 422380
rect 412771 422315 412837 422316
rect 408539 420204 408605 420205
rect 408539 420140 408540 420204
rect 408604 420140 408605 420204
rect 408539 420139 408605 420140
rect 209568 417454 209888 417486
rect 209568 417218 209610 417454
rect 209846 417218 209888 417454
rect 209568 417134 209888 417218
rect 209568 416898 209610 417134
rect 209846 416898 209888 417134
rect 209568 416866 209888 416898
rect 240288 417454 240608 417486
rect 240288 417218 240330 417454
rect 240566 417218 240608 417454
rect 240288 417134 240608 417218
rect 240288 416898 240330 417134
rect 240566 416898 240608 417134
rect 240288 416866 240608 416898
rect 271008 417454 271328 417486
rect 271008 417218 271050 417454
rect 271286 417218 271328 417454
rect 271008 417134 271328 417218
rect 271008 416898 271050 417134
rect 271286 416898 271328 417134
rect 271008 416866 271328 416898
rect 301728 417454 302048 417486
rect 301728 417218 301770 417454
rect 302006 417218 302048 417454
rect 301728 417134 302048 417218
rect 301728 416898 301770 417134
rect 302006 416898 302048 417134
rect 301728 416866 302048 416898
rect 332448 417454 332768 417486
rect 332448 417218 332490 417454
rect 332726 417218 332768 417454
rect 332448 417134 332768 417218
rect 332448 416898 332490 417134
rect 332726 416898 332768 417134
rect 332448 416866 332768 416898
rect 363168 417454 363488 417486
rect 363168 417218 363210 417454
rect 363446 417218 363488 417454
rect 363168 417134 363488 417218
rect 363168 416898 363210 417134
rect 363446 416898 363488 417134
rect 363168 416866 363488 416898
rect 393888 417454 394208 417486
rect 393888 417218 393930 417454
rect 394166 417218 394208 417454
rect 393888 417134 394208 417218
rect 393888 416898 393930 417134
rect 394166 416898 394208 417134
rect 393888 416866 394208 416898
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 194208 399454 194528 399486
rect 194208 399218 194250 399454
rect 194486 399218 194528 399454
rect 194208 399134 194528 399218
rect 194208 398898 194250 399134
rect 194486 398898 194528 399134
rect 194208 398866 194528 398898
rect 224928 399454 225248 399486
rect 224928 399218 224970 399454
rect 225206 399218 225248 399454
rect 224928 399134 225248 399218
rect 224928 398898 224970 399134
rect 225206 398898 225248 399134
rect 224928 398866 225248 398898
rect 255648 399454 255968 399486
rect 255648 399218 255690 399454
rect 255926 399218 255968 399454
rect 255648 399134 255968 399218
rect 255648 398898 255690 399134
rect 255926 398898 255968 399134
rect 255648 398866 255968 398898
rect 286368 399454 286688 399486
rect 286368 399218 286410 399454
rect 286646 399218 286688 399454
rect 286368 399134 286688 399218
rect 286368 398898 286410 399134
rect 286646 398898 286688 399134
rect 286368 398866 286688 398898
rect 317088 399454 317408 399486
rect 317088 399218 317130 399454
rect 317366 399218 317408 399454
rect 317088 399134 317408 399218
rect 317088 398898 317130 399134
rect 317366 398898 317408 399134
rect 317088 398866 317408 398898
rect 347808 399454 348128 399486
rect 347808 399218 347850 399454
rect 348086 399218 348128 399454
rect 347808 399134 348128 399218
rect 347808 398898 347850 399134
rect 348086 398898 348128 399134
rect 347808 398866 348128 398898
rect 378528 399454 378848 399486
rect 378528 399218 378570 399454
rect 378806 399218 378848 399454
rect 378528 399134 378848 399218
rect 378528 398898 378570 399134
rect 378806 398898 378848 399134
rect 378528 398866 378848 398898
rect 209568 381454 209888 381486
rect 209568 381218 209610 381454
rect 209846 381218 209888 381454
rect 209568 381134 209888 381218
rect 209568 380898 209610 381134
rect 209846 380898 209888 381134
rect 209568 380866 209888 380898
rect 240288 381454 240608 381486
rect 240288 381218 240330 381454
rect 240566 381218 240608 381454
rect 240288 381134 240608 381218
rect 240288 380898 240330 381134
rect 240566 380898 240608 381134
rect 240288 380866 240608 380898
rect 271008 381454 271328 381486
rect 271008 381218 271050 381454
rect 271286 381218 271328 381454
rect 271008 381134 271328 381218
rect 271008 380898 271050 381134
rect 271286 380898 271328 381134
rect 271008 380866 271328 380898
rect 301728 381454 302048 381486
rect 301728 381218 301770 381454
rect 302006 381218 302048 381454
rect 301728 381134 302048 381218
rect 301728 380898 301770 381134
rect 302006 380898 302048 381134
rect 301728 380866 302048 380898
rect 332448 381454 332768 381486
rect 332448 381218 332490 381454
rect 332726 381218 332768 381454
rect 332448 381134 332768 381218
rect 332448 380898 332490 381134
rect 332726 380898 332768 381134
rect 332448 380866 332768 380898
rect 363168 381454 363488 381486
rect 363168 381218 363210 381454
rect 363446 381218 363488 381454
rect 363168 381134 363488 381218
rect 363168 380898 363210 381134
rect 363446 380898 363488 381134
rect 363168 380866 363488 380898
rect 393888 381454 394208 381486
rect 393888 381218 393930 381454
rect 394166 381218 394208 381454
rect 393888 381134 394208 381218
rect 393888 380898 393930 381134
rect 394166 380898 394208 381134
rect 393888 380866 394208 380898
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 194208 363454 194528 363486
rect 194208 363218 194250 363454
rect 194486 363218 194528 363454
rect 194208 363134 194528 363218
rect 194208 362898 194250 363134
rect 194486 362898 194528 363134
rect 194208 362866 194528 362898
rect 224928 363454 225248 363486
rect 224928 363218 224970 363454
rect 225206 363218 225248 363454
rect 224928 363134 225248 363218
rect 224928 362898 224970 363134
rect 225206 362898 225248 363134
rect 224928 362866 225248 362898
rect 255648 363454 255968 363486
rect 255648 363218 255690 363454
rect 255926 363218 255968 363454
rect 255648 363134 255968 363218
rect 255648 362898 255690 363134
rect 255926 362898 255968 363134
rect 255648 362866 255968 362898
rect 286368 363454 286688 363486
rect 286368 363218 286410 363454
rect 286646 363218 286688 363454
rect 286368 363134 286688 363218
rect 286368 362898 286410 363134
rect 286646 362898 286688 363134
rect 286368 362866 286688 362898
rect 317088 363454 317408 363486
rect 317088 363218 317130 363454
rect 317366 363218 317408 363454
rect 317088 363134 317408 363218
rect 317088 362898 317130 363134
rect 317366 362898 317408 363134
rect 317088 362866 317408 362898
rect 347808 363454 348128 363486
rect 347808 363218 347850 363454
rect 348086 363218 348128 363454
rect 347808 363134 348128 363218
rect 347808 362898 347850 363134
rect 348086 362898 348128 363134
rect 347808 362866 348128 362898
rect 378528 363454 378848 363486
rect 378528 363218 378570 363454
rect 378806 363218 378848 363454
rect 378528 363134 378848 363218
rect 378528 362898 378570 363134
rect 378806 362898 378848 363134
rect 378528 362866 378848 362898
rect 209568 345454 209888 345486
rect 209568 345218 209610 345454
rect 209846 345218 209888 345454
rect 209568 345134 209888 345218
rect 209568 344898 209610 345134
rect 209846 344898 209888 345134
rect 209568 344866 209888 344898
rect 240288 345454 240608 345486
rect 240288 345218 240330 345454
rect 240566 345218 240608 345454
rect 240288 345134 240608 345218
rect 240288 344898 240330 345134
rect 240566 344898 240608 345134
rect 240288 344866 240608 344898
rect 271008 345454 271328 345486
rect 271008 345218 271050 345454
rect 271286 345218 271328 345454
rect 271008 345134 271328 345218
rect 271008 344898 271050 345134
rect 271286 344898 271328 345134
rect 271008 344866 271328 344898
rect 301728 345454 302048 345486
rect 301728 345218 301770 345454
rect 302006 345218 302048 345454
rect 301728 345134 302048 345218
rect 301728 344898 301770 345134
rect 302006 344898 302048 345134
rect 301728 344866 302048 344898
rect 332448 345454 332768 345486
rect 332448 345218 332490 345454
rect 332726 345218 332768 345454
rect 332448 345134 332768 345218
rect 332448 344898 332490 345134
rect 332726 344898 332768 345134
rect 332448 344866 332768 344898
rect 363168 345454 363488 345486
rect 363168 345218 363210 345454
rect 363446 345218 363488 345454
rect 363168 345134 363488 345218
rect 363168 344898 363210 345134
rect 363446 344898 363488 345134
rect 363168 344866 363488 344898
rect 393888 345454 394208 345486
rect 393888 345218 393930 345454
rect 394166 345218 394208 345454
rect 393888 345134 394208 345218
rect 393888 344898 393930 345134
rect 394166 344898 394208 345134
rect 393888 344866 394208 344898
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 194208 327454 194528 327486
rect 194208 327218 194250 327454
rect 194486 327218 194528 327454
rect 194208 327134 194528 327218
rect 194208 326898 194250 327134
rect 194486 326898 194528 327134
rect 194208 326866 194528 326898
rect 224928 327454 225248 327486
rect 224928 327218 224970 327454
rect 225206 327218 225248 327454
rect 224928 327134 225248 327218
rect 224928 326898 224970 327134
rect 225206 326898 225248 327134
rect 224928 326866 225248 326898
rect 255648 327454 255968 327486
rect 255648 327218 255690 327454
rect 255926 327218 255968 327454
rect 255648 327134 255968 327218
rect 255648 326898 255690 327134
rect 255926 326898 255968 327134
rect 255648 326866 255968 326898
rect 286368 327454 286688 327486
rect 286368 327218 286410 327454
rect 286646 327218 286688 327454
rect 286368 327134 286688 327218
rect 286368 326898 286410 327134
rect 286646 326898 286688 327134
rect 286368 326866 286688 326898
rect 317088 327454 317408 327486
rect 317088 327218 317130 327454
rect 317366 327218 317408 327454
rect 317088 327134 317408 327218
rect 317088 326898 317130 327134
rect 317366 326898 317408 327134
rect 317088 326866 317408 326898
rect 347808 327454 348128 327486
rect 347808 327218 347850 327454
rect 348086 327218 348128 327454
rect 347808 327134 348128 327218
rect 347808 326898 347850 327134
rect 348086 326898 348128 327134
rect 347808 326866 348128 326898
rect 378528 327454 378848 327486
rect 378528 327218 378570 327454
rect 378806 327218 378848 327454
rect 378528 327134 378848 327218
rect 378528 326898 378570 327134
rect 378806 326898 378848 327134
rect 378528 326866 378848 326898
rect 209568 309454 209888 309486
rect 209568 309218 209610 309454
rect 209846 309218 209888 309454
rect 209568 309134 209888 309218
rect 209568 308898 209610 309134
rect 209846 308898 209888 309134
rect 209568 308866 209888 308898
rect 240288 309454 240608 309486
rect 240288 309218 240330 309454
rect 240566 309218 240608 309454
rect 240288 309134 240608 309218
rect 240288 308898 240330 309134
rect 240566 308898 240608 309134
rect 240288 308866 240608 308898
rect 271008 309454 271328 309486
rect 271008 309218 271050 309454
rect 271286 309218 271328 309454
rect 271008 309134 271328 309218
rect 271008 308898 271050 309134
rect 271286 308898 271328 309134
rect 271008 308866 271328 308898
rect 301728 309454 302048 309486
rect 301728 309218 301770 309454
rect 302006 309218 302048 309454
rect 301728 309134 302048 309218
rect 301728 308898 301770 309134
rect 302006 308898 302048 309134
rect 301728 308866 302048 308898
rect 332448 309454 332768 309486
rect 332448 309218 332490 309454
rect 332726 309218 332768 309454
rect 332448 309134 332768 309218
rect 332448 308898 332490 309134
rect 332726 308898 332768 309134
rect 332448 308866 332768 308898
rect 363168 309454 363488 309486
rect 363168 309218 363210 309454
rect 363446 309218 363488 309454
rect 363168 309134 363488 309218
rect 363168 308898 363210 309134
rect 363446 308898 363488 309134
rect 363168 308866 363488 308898
rect 393888 309454 394208 309486
rect 393888 309218 393930 309454
rect 394166 309218 394208 309454
rect 393888 309134 394208 309218
rect 393888 308898 393930 309134
rect 394166 308898 394208 309134
rect 393888 308866 394208 308898
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 194208 291454 194528 291486
rect 194208 291218 194250 291454
rect 194486 291218 194528 291454
rect 194208 291134 194528 291218
rect 194208 290898 194250 291134
rect 194486 290898 194528 291134
rect 194208 290866 194528 290898
rect 224928 291454 225248 291486
rect 224928 291218 224970 291454
rect 225206 291218 225248 291454
rect 224928 291134 225248 291218
rect 224928 290898 224970 291134
rect 225206 290898 225248 291134
rect 224928 290866 225248 290898
rect 255648 291454 255968 291486
rect 255648 291218 255690 291454
rect 255926 291218 255968 291454
rect 255648 291134 255968 291218
rect 255648 290898 255690 291134
rect 255926 290898 255968 291134
rect 255648 290866 255968 290898
rect 286368 291454 286688 291486
rect 286368 291218 286410 291454
rect 286646 291218 286688 291454
rect 286368 291134 286688 291218
rect 286368 290898 286410 291134
rect 286646 290898 286688 291134
rect 286368 290866 286688 290898
rect 317088 291454 317408 291486
rect 317088 291218 317130 291454
rect 317366 291218 317408 291454
rect 317088 291134 317408 291218
rect 317088 290898 317130 291134
rect 317366 290898 317408 291134
rect 317088 290866 317408 290898
rect 347808 291454 348128 291486
rect 347808 291218 347850 291454
rect 348086 291218 348128 291454
rect 347808 291134 348128 291218
rect 347808 290898 347850 291134
rect 348086 290898 348128 291134
rect 347808 290866 348128 290898
rect 378528 291454 378848 291486
rect 378528 291218 378570 291454
rect 378806 291218 378848 291454
rect 378528 291134 378848 291218
rect 378528 290898 378570 291134
rect 378806 290898 378848 291134
rect 378528 290866 378848 290898
rect 209568 273454 209888 273486
rect 209568 273218 209610 273454
rect 209846 273218 209888 273454
rect 209568 273134 209888 273218
rect 209568 272898 209610 273134
rect 209846 272898 209888 273134
rect 209568 272866 209888 272898
rect 240288 273454 240608 273486
rect 240288 273218 240330 273454
rect 240566 273218 240608 273454
rect 240288 273134 240608 273218
rect 240288 272898 240330 273134
rect 240566 272898 240608 273134
rect 240288 272866 240608 272898
rect 271008 273454 271328 273486
rect 271008 273218 271050 273454
rect 271286 273218 271328 273454
rect 271008 273134 271328 273218
rect 271008 272898 271050 273134
rect 271286 272898 271328 273134
rect 271008 272866 271328 272898
rect 301728 273454 302048 273486
rect 301728 273218 301770 273454
rect 302006 273218 302048 273454
rect 301728 273134 302048 273218
rect 301728 272898 301770 273134
rect 302006 272898 302048 273134
rect 301728 272866 302048 272898
rect 332448 273454 332768 273486
rect 332448 273218 332490 273454
rect 332726 273218 332768 273454
rect 332448 273134 332768 273218
rect 332448 272898 332490 273134
rect 332726 272898 332768 273134
rect 332448 272866 332768 272898
rect 363168 273454 363488 273486
rect 363168 273218 363210 273454
rect 363446 273218 363488 273454
rect 363168 273134 363488 273218
rect 363168 272898 363210 273134
rect 363446 272898 363488 273134
rect 363168 272866 363488 272898
rect 393888 273454 394208 273486
rect 393888 273218 393930 273454
rect 394166 273218 394208 273454
rect 393888 273134 394208 273218
rect 393888 272898 393930 273134
rect 394166 272898 394208 273134
rect 393888 272866 394208 272898
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 194208 255454 194528 255486
rect 194208 255218 194250 255454
rect 194486 255218 194528 255454
rect 194208 255134 194528 255218
rect 194208 254898 194250 255134
rect 194486 254898 194528 255134
rect 194208 254866 194528 254898
rect 224928 255454 225248 255486
rect 224928 255218 224970 255454
rect 225206 255218 225248 255454
rect 224928 255134 225248 255218
rect 224928 254898 224970 255134
rect 225206 254898 225248 255134
rect 224928 254866 225248 254898
rect 255648 255454 255968 255486
rect 255648 255218 255690 255454
rect 255926 255218 255968 255454
rect 255648 255134 255968 255218
rect 255648 254898 255690 255134
rect 255926 254898 255968 255134
rect 255648 254866 255968 254898
rect 286368 255454 286688 255486
rect 286368 255218 286410 255454
rect 286646 255218 286688 255454
rect 286368 255134 286688 255218
rect 286368 254898 286410 255134
rect 286646 254898 286688 255134
rect 286368 254866 286688 254898
rect 317088 255454 317408 255486
rect 317088 255218 317130 255454
rect 317366 255218 317408 255454
rect 317088 255134 317408 255218
rect 317088 254898 317130 255134
rect 317366 254898 317408 255134
rect 317088 254866 317408 254898
rect 347808 255454 348128 255486
rect 347808 255218 347850 255454
rect 348086 255218 348128 255454
rect 347808 255134 348128 255218
rect 347808 254898 347850 255134
rect 348086 254898 348128 255134
rect 347808 254866 348128 254898
rect 378528 255454 378848 255486
rect 378528 255218 378570 255454
rect 378806 255218 378848 255454
rect 378528 255134 378848 255218
rect 378528 254898 378570 255134
rect 378806 254898 378848 255134
rect 378528 254866 378848 254898
rect 209568 237454 209888 237486
rect 209568 237218 209610 237454
rect 209846 237218 209888 237454
rect 209568 237134 209888 237218
rect 209568 236898 209610 237134
rect 209846 236898 209888 237134
rect 209568 236866 209888 236898
rect 240288 237454 240608 237486
rect 240288 237218 240330 237454
rect 240566 237218 240608 237454
rect 240288 237134 240608 237218
rect 240288 236898 240330 237134
rect 240566 236898 240608 237134
rect 240288 236866 240608 236898
rect 271008 237454 271328 237486
rect 271008 237218 271050 237454
rect 271286 237218 271328 237454
rect 271008 237134 271328 237218
rect 271008 236898 271050 237134
rect 271286 236898 271328 237134
rect 271008 236866 271328 236898
rect 301728 237454 302048 237486
rect 301728 237218 301770 237454
rect 302006 237218 302048 237454
rect 301728 237134 302048 237218
rect 301728 236898 301770 237134
rect 302006 236898 302048 237134
rect 301728 236866 302048 236898
rect 332448 237454 332768 237486
rect 332448 237218 332490 237454
rect 332726 237218 332768 237454
rect 332448 237134 332768 237218
rect 332448 236898 332490 237134
rect 332726 236898 332768 237134
rect 332448 236866 332768 236898
rect 363168 237454 363488 237486
rect 363168 237218 363210 237454
rect 363446 237218 363488 237454
rect 363168 237134 363488 237218
rect 363168 236898 363210 237134
rect 363446 236898 363488 237134
rect 363168 236866 363488 236898
rect 393888 237454 394208 237486
rect 393888 237218 393930 237454
rect 394166 237218 394208 237454
rect 393888 237134 394208 237218
rect 393888 236898 393930 237134
rect 394166 236898 394208 237134
rect 393888 236866 394208 236898
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 194208 219454 194528 219486
rect 194208 219218 194250 219454
rect 194486 219218 194528 219454
rect 194208 219134 194528 219218
rect 194208 218898 194250 219134
rect 194486 218898 194528 219134
rect 194208 218866 194528 218898
rect 224928 219454 225248 219486
rect 224928 219218 224970 219454
rect 225206 219218 225248 219454
rect 224928 219134 225248 219218
rect 224928 218898 224970 219134
rect 225206 218898 225248 219134
rect 224928 218866 225248 218898
rect 255648 219454 255968 219486
rect 255648 219218 255690 219454
rect 255926 219218 255968 219454
rect 255648 219134 255968 219218
rect 255648 218898 255690 219134
rect 255926 218898 255968 219134
rect 255648 218866 255968 218898
rect 286368 219454 286688 219486
rect 286368 219218 286410 219454
rect 286646 219218 286688 219454
rect 286368 219134 286688 219218
rect 286368 218898 286410 219134
rect 286646 218898 286688 219134
rect 286368 218866 286688 218898
rect 317088 219454 317408 219486
rect 317088 219218 317130 219454
rect 317366 219218 317408 219454
rect 317088 219134 317408 219218
rect 317088 218898 317130 219134
rect 317366 218898 317408 219134
rect 317088 218866 317408 218898
rect 347808 219454 348128 219486
rect 347808 219218 347850 219454
rect 348086 219218 348128 219454
rect 347808 219134 348128 219218
rect 347808 218898 347850 219134
rect 348086 218898 348128 219134
rect 347808 218866 348128 218898
rect 378528 219454 378848 219486
rect 378528 219218 378570 219454
rect 378806 219218 378848 219454
rect 378528 219134 378848 219218
rect 378528 218898 378570 219134
rect 378806 218898 378848 219134
rect 378528 218866 378848 218898
rect 399523 199612 399589 199613
rect 399523 199548 399524 199612
rect 399588 199548 399589 199612
rect 399523 199547 399589 199548
rect 399339 199340 399405 199341
rect 399339 199276 399340 199340
rect 399404 199276 399405 199340
rect 399339 199275 399405 199276
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 142000 186134 150618
rect 189234 190894 189854 198000
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 142000 189854 154338
rect 192954 194614 193574 198000
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 142000 193574 158058
rect 199794 165454 200414 198000
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 142000 200414 164898
rect 203514 169174 204134 198000
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 142000 204134 168618
rect 207234 172894 207854 198000
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 142000 207854 172338
rect 210954 176614 211574 198000
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 142000 211574 176058
rect 217794 183454 218414 198000
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 147454 218414 182898
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 142000 218414 146898
rect 221514 187174 222134 198000
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 151174 222134 186618
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 142000 222134 150618
rect 225234 190894 225854 198000
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 154894 225854 190338
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 142000 225854 154338
rect 228954 194614 229574 198000
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 142000 229574 158058
rect 235794 165454 236414 198000
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 142000 236414 164898
rect 239514 169174 240134 198000
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 142000 240134 168618
rect 243234 172894 243854 198000
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 142000 243854 172338
rect 246954 176614 247574 198000
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 142000 247574 176058
rect 253794 183454 254414 198000
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 142000 254414 146898
rect 257514 187174 258134 198000
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 142000 258134 150618
rect 261234 190894 261854 198000
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 142000 261854 154338
rect 264954 194614 265574 198000
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 142000 265574 158058
rect 271794 165454 272414 198000
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 142000 272414 164898
rect 275514 169174 276134 198000
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 142000 276134 168618
rect 279234 172894 279854 198000
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 142000 279854 172338
rect 282954 176614 283574 198000
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 169339 140044 169405 140045
rect 169339 139980 169340 140044
rect 169404 139980 169405 140044
rect 169339 139979 169405 139980
rect 169155 129436 169221 129437
rect 169155 129372 169156 129436
rect 169220 129372 169221 129436
rect 169155 129371 169221 129372
rect 168235 121276 168301 121277
rect 168235 121212 168236 121276
rect 168300 121212 168301 121276
rect 168235 121211 168301 121212
rect 169342 91629 169402 139979
rect 169523 139908 169589 139909
rect 169523 139844 169524 139908
rect 169588 139844 169589 139908
rect 169523 139843 169589 139844
rect 169526 93261 169586 139843
rect 189568 129454 189888 129486
rect 189568 129218 189610 129454
rect 189846 129218 189888 129454
rect 189568 129134 189888 129218
rect 189568 128898 189610 129134
rect 189846 128898 189888 129134
rect 189568 128866 189888 128898
rect 220288 129454 220608 129486
rect 220288 129218 220330 129454
rect 220566 129218 220608 129454
rect 220288 129134 220608 129218
rect 220288 128898 220330 129134
rect 220566 128898 220608 129134
rect 220288 128866 220608 128898
rect 251008 129454 251328 129486
rect 251008 129218 251050 129454
rect 251286 129218 251328 129454
rect 251008 129134 251328 129218
rect 251008 128898 251050 129134
rect 251286 128898 251328 129134
rect 251008 128866 251328 128898
rect 174208 111454 174528 111486
rect 174208 111218 174250 111454
rect 174486 111218 174528 111454
rect 174208 111134 174528 111218
rect 174208 110898 174250 111134
rect 174486 110898 174528 111134
rect 174208 110866 174528 110898
rect 204928 111454 205248 111486
rect 204928 111218 204970 111454
rect 205206 111218 205248 111454
rect 204928 111134 205248 111218
rect 204928 110898 204970 111134
rect 205206 110898 205248 111134
rect 204928 110866 205248 110898
rect 235648 111454 235968 111486
rect 235648 111218 235690 111454
rect 235926 111218 235968 111454
rect 235648 111134 235968 111218
rect 235648 110898 235690 111134
rect 235926 110898 235968 111134
rect 235648 110866 235968 110898
rect 266368 111454 266688 111486
rect 266368 111218 266410 111454
rect 266646 111218 266688 111454
rect 266368 111134 266688 111218
rect 266368 110898 266410 111134
rect 266646 110898 266688 111134
rect 266368 110866 266688 110898
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 189568 93454 189888 93486
rect 169523 93260 169589 93261
rect 169523 93196 169524 93260
rect 169588 93196 169589 93260
rect 169523 93195 169589 93196
rect 189568 93218 189610 93454
rect 189846 93218 189888 93454
rect 189568 93134 189888 93218
rect 189568 92898 189610 93134
rect 189846 92898 189888 93134
rect 189568 92866 189888 92898
rect 220288 93454 220608 93486
rect 220288 93218 220330 93454
rect 220566 93218 220608 93454
rect 220288 93134 220608 93218
rect 220288 92898 220330 93134
rect 220566 92898 220608 93134
rect 220288 92866 220608 92898
rect 251008 93454 251328 93486
rect 251008 93218 251050 93454
rect 251286 93218 251328 93454
rect 251008 93134 251328 93218
rect 251008 92898 251050 93134
rect 251286 92898 251328 93134
rect 251008 92866 251328 92898
rect 169339 91628 169405 91629
rect 169339 91564 169340 91628
rect 169404 91564 169405 91628
rect 169339 91563 169405 91564
rect 167683 85100 167749 85101
rect 167683 85036 167684 85100
rect 167748 85036 167749 85100
rect 167683 85035 167749 85036
rect 168235 78572 168301 78573
rect 168235 78508 168236 78572
rect 168300 78508 168301 78572
rect 168235 78507 168301 78508
rect 168051 63748 168117 63749
rect 168051 63684 168052 63748
rect 168116 63684 168117 63748
rect 168051 63683 168117 63684
rect 167683 60484 167749 60485
rect 167683 60420 167684 60484
rect 167748 60420 167749 60484
rect 167683 60419 167749 60420
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 167686 29610 167746 60419
rect 167867 57220 167933 57221
rect 167867 57156 167868 57220
rect 167932 57156 167933 57220
rect 167867 57155 167933 57156
rect 167870 30021 167930 57155
rect 168054 30701 168114 63683
rect 168238 41445 168298 78507
rect 174208 75454 174528 75486
rect 174208 75218 174250 75454
rect 174486 75218 174528 75454
rect 174208 75134 174528 75218
rect 174208 74898 174250 75134
rect 174486 74898 174528 75134
rect 174208 74866 174528 74898
rect 204928 75454 205248 75486
rect 204928 75218 204970 75454
rect 205206 75218 205248 75454
rect 204928 75134 205248 75218
rect 204928 74898 204970 75134
rect 205206 74898 205248 75134
rect 204928 74866 205248 74898
rect 235648 75454 235968 75486
rect 235648 75218 235690 75454
rect 235926 75218 235968 75454
rect 235648 75134 235968 75218
rect 235648 74898 235690 75134
rect 235926 74898 235968 75134
rect 235648 74866 235968 74898
rect 266368 75454 266688 75486
rect 266368 75218 266410 75454
rect 266646 75218 266688 75454
rect 266368 75134 266688 75218
rect 266368 74898 266410 75134
rect 266646 74898 266688 75134
rect 266368 74866 266688 74898
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 189568 57454 189888 57486
rect 189568 57218 189610 57454
rect 189846 57218 189888 57454
rect 189568 57134 189888 57218
rect 189568 56898 189610 57134
rect 189846 56898 189888 57134
rect 189568 56866 189888 56898
rect 220288 57454 220608 57486
rect 220288 57218 220330 57454
rect 220566 57218 220608 57454
rect 220288 57134 220608 57218
rect 220288 56898 220330 57134
rect 220566 56898 220608 57134
rect 220288 56866 220608 56898
rect 251008 57454 251328 57486
rect 251008 57218 251050 57454
rect 251286 57218 251328 57454
rect 251008 57134 251328 57218
rect 251008 56898 251050 57134
rect 251286 56898 251328 57134
rect 251008 56866 251328 56898
rect 168235 41444 168301 41445
rect 168235 41380 168236 41444
rect 168300 41380 168301 41444
rect 168235 41379 168301 41380
rect 168235 40764 168301 40765
rect 168235 40700 168236 40764
rect 168300 40700 168301 40764
rect 168235 40699 168301 40700
rect 168051 30700 168117 30701
rect 168051 30636 168052 30700
rect 168116 30636 168117 30700
rect 168051 30635 168117 30636
rect 167867 30020 167933 30021
rect 167867 29956 167868 30020
rect 167932 29956 167933 30020
rect 167867 29955 167933 29956
rect 168238 29885 168298 40699
rect 168971 39948 169037 39949
rect 168971 39884 168972 39948
rect 169036 39884 169037 39948
rect 168971 39883 169037 39884
rect 168974 30157 169034 39883
rect 174208 39454 174528 39486
rect 174208 39218 174250 39454
rect 174486 39218 174528 39454
rect 174208 39134 174528 39218
rect 174208 38898 174250 39134
rect 174486 38898 174528 39134
rect 174208 38866 174528 38898
rect 204928 39454 205248 39486
rect 204928 39218 204970 39454
rect 205206 39218 205248 39454
rect 204928 39134 205248 39218
rect 204928 38898 204970 39134
rect 205206 38898 205248 39134
rect 204928 38866 205248 38898
rect 235648 39454 235968 39486
rect 235648 39218 235690 39454
rect 235926 39218 235968 39454
rect 235648 39134 235968 39218
rect 235648 38898 235690 39134
rect 235926 38898 235968 39134
rect 235648 38866 235968 38898
rect 266368 39454 266688 39486
rect 266368 39218 266410 39454
rect 266646 39218 266688 39454
rect 266368 39134 266688 39218
rect 266368 38898 266410 39134
rect 266646 38898 266688 39134
rect 266368 38866 266688 38898
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 168971 30156 169037 30157
rect 168971 30092 168972 30156
rect 169036 30092 169037 30156
rect 168971 30091 169037 30092
rect 168235 29884 168301 29885
rect 168235 29820 168236 29884
rect 168300 29820 168301 29884
rect 168235 29819 168301 29820
rect 167686 29550 168298 29610
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 28000
rect 168238 27573 168298 29550
rect 168235 27572 168301 27573
rect 168235 27508 168236 27572
rect 168300 27508 168301 27572
rect 168235 27507 168301 27508
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 28000
rect 181794 3454 182414 28000
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 7174 186134 28000
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 28000
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 14614 193574 28000
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 28000
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 28000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 28000
rect 217794 3454 218414 28000
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 7174 222134 28000
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 10894 225854 28000
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 28000
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 28000
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 28000
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 28000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 28000
rect 253794 3454 254414 28000
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 28000
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 28000
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 28000
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 28000
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 28000
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 28000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 183454 290414 198000
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 187174 294134 198000
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 190894 297854 198000
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 194614 301574 198000
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 165454 308414 198000
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 169174 312134 198000
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 172894 315854 198000
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 176614 319574 198000
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 183454 326414 198000
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 187174 330134 198000
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 190894 333854 198000
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 194614 337574 198000
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 165454 344414 198000
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 169174 348134 198000
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 172894 351854 198000
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 176614 355574 198000
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 183454 362414 198000
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 187174 366134 198000
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 190894 369854 198000
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 194614 373574 198000
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 165454 380414 198000
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 169174 384134 198000
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 172894 387854 198000
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 176614 391574 198000
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 397794 183454 398414 198000
rect 398603 196620 398669 196621
rect 398603 196556 398604 196620
rect 398668 196556 398669 196620
rect 398603 196555 398669 196556
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 142000 398414 146898
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 398051 139500 398117 139501
rect 398051 139436 398052 139500
rect 398116 139436 398117 139500
rect 398051 139435 398117 139436
rect 398054 106453 398114 139435
rect 398606 137597 398666 196555
rect 398787 139500 398853 139501
rect 398787 139436 398788 139500
rect 398852 139436 398853 139500
rect 398787 139435 398853 139436
rect 398603 137596 398669 137597
rect 398603 137532 398604 137596
rect 398668 137532 398669 137596
rect 398603 137531 398669 137532
rect 398790 108085 398850 139435
rect 398787 108084 398853 108085
rect 398787 108020 398788 108084
rect 398852 108020 398853 108084
rect 398787 108019 398853 108020
rect 398051 106452 398117 106453
rect 398051 106388 398052 106452
rect 398116 106388 398117 106452
rect 398051 106387 398117 106388
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 397867 63476 397933 63477
rect 397867 63412 397868 63476
rect 397932 63412 397933 63476
rect 397867 63411 397933 63412
rect 397683 59260 397749 59261
rect 397683 59196 397684 59260
rect 397748 59196 397749 59260
rect 397683 59195 397749 59196
rect 397499 33148 397565 33149
rect 397499 33084 397500 33148
rect 397564 33084 397565 33148
rect 397499 33083 397565 33084
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397502 30293 397562 33083
rect 397499 30292 397565 30293
rect 397499 30228 397500 30292
rect 397564 30228 397565 30292
rect 397499 30227 397565 30228
rect 397686 28250 397746 59195
rect 397870 30701 397930 63411
rect 397867 30700 397933 30701
rect 397867 30636 397868 30700
rect 397932 30636 397933 30700
rect 397867 30635 397933 30636
rect 399342 28389 399402 199275
rect 399526 28525 399586 199547
rect 399707 194172 399773 194173
rect 399707 194108 399708 194172
rect 399772 194108 399773 194172
rect 399707 194107 399773 194108
rect 399710 139501 399770 194107
rect 401514 187174 402134 198000
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 142000 402134 150618
rect 405234 190894 405854 198000
rect 408542 196077 408602 420139
rect 409827 408916 409893 408917
rect 409827 408852 409828 408916
rect 409892 408852 409893 408916
rect 409827 408851 409893 408852
rect 409459 225044 409525 225045
rect 409459 224980 409460 225044
rect 409524 224980 409525 225044
rect 409459 224979 409525 224980
rect 409462 219450 409522 224979
rect 409094 219390 409522 219450
rect 409094 199613 409154 219390
rect 409091 199612 409157 199613
rect 409091 199548 409092 199612
rect 409156 199548 409157 199612
rect 409091 199547 409157 199548
rect 408539 196076 408605 196077
rect 408539 196012 408540 196076
rect 408604 196012 408605 196076
rect 408539 196011 408605 196012
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 142000 405854 154338
rect 408954 194614 409574 198000
rect 409830 195397 409890 408851
rect 412403 401980 412469 401981
rect 412403 401916 412404 401980
rect 412468 401916 412469 401980
rect 412403 401915 412469 401916
rect 410011 377364 410077 377365
rect 410011 377300 410012 377364
rect 410076 377300 410077 377364
rect 410011 377299 410077 377300
rect 409827 195396 409893 195397
rect 409827 195332 409828 195396
rect 409892 195332 409893 195396
rect 409827 195331 409893 195332
rect 410014 195261 410074 377299
rect 411299 301748 411365 301749
rect 411299 301684 411300 301748
rect 411364 301684 411365 301748
rect 411299 301683 411365 301684
rect 410011 195260 410077 195261
rect 410011 195196 410012 195260
rect 410076 195196 410077 195260
rect 410011 195195 410077 195196
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 142000 409574 158058
rect 411302 142765 411362 301683
rect 411483 297668 411549 297669
rect 411483 297604 411484 297668
rect 411548 297604 411549 297668
rect 411483 297603 411549 297604
rect 411486 194173 411546 297603
rect 411667 240140 411733 240141
rect 411667 240076 411668 240140
rect 411732 240076 411733 240140
rect 411667 240075 411733 240076
rect 411483 194172 411549 194173
rect 411483 194108 411484 194172
rect 411548 194108 411549 194172
rect 411483 194107 411549 194108
rect 411670 144125 411730 240075
rect 411851 215388 411917 215389
rect 411851 215324 411852 215388
rect 411916 215324 411917 215388
rect 411851 215323 411917 215324
rect 411854 199477 411914 215323
rect 411851 199476 411917 199477
rect 411851 199412 411852 199476
rect 411916 199412 411917 199476
rect 411851 199411 411917 199412
rect 412406 145621 412466 401915
rect 412774 199341 412834 422315
rect 414611 421020 414677 421021
rect 414611 420956 414612 421020
rect 414676 420956 414677 421020
rect 414611 420955 414677 420956
rect 412955 406740 413021 406741
rect 412955 406676 412956 406740
rect 413020 406676 413021 406740
rect 412955 406675 413021 406676
rect 412771 199340 412837 199341
rect 412771 199276 412772 199340
rect 412836 199276 412837 199340
rect 412771 199275 412837 199276
rect 412958 192541 413018 406675
rect 412955 192540 413021 192541
rect 412955 192476 412956 192540
rect 413020 192476 413021 192540
rect 412955 192475 413021 192476
rect 412403 145620 412469 145621
rect 412403 145556 412404 145620
rect 412468 145556 412469 145620
rect 412403 145555 412469 145556
rect 411667 144124 411733 144125
rect 411667 144060 411668 144124
rect 411732 144060 411733 144124
rect 411667 144059 411733 144060
rect 414614 142765 414674 420955
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 411299 142764 411365 142765
rect 411299 142700 411300 142764
rect 411364 142700 411365 142764
rect 411299 142699 411365 142700
rect 414611 142764 414677 142765
rect 414611 142700 414612 142764
rect 414676 142700 414677 142764
rect 414611 142699 414677 142700
rect 415794 142000 416414 164898
rect 419514 493174 420134 498000
rect 420502 496909 420562 499530
rect 421790 496909 421850 499530
rect 423078 499530 423188 499590
rect 424182 499530 424276 499590
rect 425440 499590 425500 500106
rect 426528 499590 426588 500106
rect 427616 499590 427676 500106
rect 428296 499590 428356 500106
rect 428704 499590 428764 500106
rect 425440 499530 425530 499590
rect 426528 499530 426634 499590
rect 427616 499530 427738 499590
rect 423078 496909 423138 499530
rect 420499 496908 420565 496909
rect 420499 496844 420500 496908
rect 420564 496844 420565 496908
rect 420499 496843 420565 496844
rect 421787 496908 421853 496909
rect 421787 496844 421788 496908
rect 421852 496844 421853 496908
rect 421787 496843 421853 496844
rect 423075 496908 423141 496909
rect 423075 496844 423076 496908
rect 423140 496844 423141 496908
rect 423075 496843 423141 496844
rect 423234 496894 423854 498000
rect 424182 496909 424242 499530
rect 425470 496909 425530 499530
rect 426574 497045 426634 499530
rect 426571 497044 426637 497045
rect 426571 496980 426572 497044
rect 426636 496980 426637 497044
rect 426571 496979 426637 496980
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 142000 420134 168618
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 424179 496908 424245 496909
rect 424179 496844 424180 496908
rect 424244 496844 424245 496908
rect 424179 496843 424245 496844
rect 425467 496908 425533 496909
rect 425467 496844 425468 496908
rect 425532 496844 425533 496908
rect 425467 496843 425533 496844
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 142000 423854 172338
rect 426954 464614 427574 498000
rect 427678 496909 427738 499530
rect 428230 499530 428356 499590
rect 428598 499530 428764 499590
rect 430064 499590 430124 500106
rect 430744 499590 430804 500106
rect 431288 499590 431348 500106
rect 432376 499590 432436 500106
rect 430064 499530 430130 499590
rect 430744 499530 430866 499590
rect 428230 497045 428290 499530
rect 428227 497044 428293 497045
rect 428227 496980 428228 497044
rect 428292 496980 428293 497044
rect 428227 496979 428293 496980
rect 428598 496909 428658 499530
rect 430070 496909 430130 499530
rect 430806 496909 430866 499530
rect 431174 499530 431348 499590
rect 432278 499530 432436 499590
rect 431174 497045 431234 499530
rect 432278 497181 432338 499530
rect 433464 499490 433524 500106
rect 433600 499590 433660 500106
rect 434552 499590 434612 500106
rect 435771 499764 435837 499765
rect 435771 499700 435772 499764
rect 435836 499700 435837 499764
rect 435771 499699 435837 499700
rect 433600 499530 433810 499590
rect 433382 499430 433524 499490
rect 432275 497180 432341 497181
rect 432275 497116 432276 497180
rect 432340 497116 432341 497180
rect 432275 497115 432341 497116
rect 431171 497044 431237 497045
rect 431171 496980 431172 497044
rect 431236 496980 431237 497044
rect 431171 496979 431237 496980
rect 433382 496909 433442 499430
rect 433750 498810 433810 499530
rect 433566 498750 433810 498810
rect 434486 499530 434612 499590
rect 433566 497045 433626 498750
rect 434486 498133 434546 499530
rect 434483 498132 434549 498133
rect 434483 498068 434484 498132
rect 434548 498068 434549 498132
rect 434483 498067 434549 498068
rect 433563 497044 433629 497045
rect 433563 496980 433564 497044
rect 433628 496980 433629 497044
rect 433563 496979 433629 496980
rect 427675 496908 427741 496909
rect 427675 496844 427676 496908
rect 427740 496844 427741 496908
rect 427675 496843 427741 496844
rect 428595 496908 428661 496909
rect 428595 496844 428596 496908
rect 428660 496844 428661 496908
rect 428595 496843 428661 496844
rect 430067 496908 430133 496909
rect 430067 496844 430068 496908
rect 430132 496844 430133 496908
rect 430067 496843 430133 496844
rect 430803 496908 430869 496909
rect 430803 496844 430804 496908
rect 430868 496844 430869 496908
rect 430803 496843 430869 496844
rect 433379 496908 433445 496909
rect 433379 496844 433380 496908
rect 433444 496844 433445 496908
rect 433379 496843 433445 496844
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 142000 427574 176058
rect 433794 471454 434414 498000
rect 435774 496909 435834 499699
rect 435912 499590 435972 500106
rect 436048 499765 436108 500106
rect 436045 499764 436111 499765
rect 436045 499700 436046 499764
rect 436110 499700 436111 499764
rect 436045 499699 436111 499700
rect 437000 499590 437060 500106
rect 435912 499530 436018 499590
rect 435958 497045 436018 499530
rect 436878 499530 437060 499590
rect 438088 499590 438148 500106
rect 438496 499590 438556 500106
rect 439448 499590 439508 500106
rect 440672 499590 440732 500106
rect 438088 499530 438410 499590
rect 438496 499530 438594 499590
rect 439448 499530 439514 499590
rect 435955 497044 436021 497045
rect 435955 496980 435956 497044
rect 436020 496980 436021 497044
rect 435955 496979 436021 496980
rect 436878 496909 436938 499530
rect 435771 496908 435837 496909
rect 435771 496844 435772 496908
rect 435836 496844 435837 496908
rect 435771 496843 435837 496844
rect 436875 496908 436941 496909
rect 436875 496844 436876 496908
rect 436940 496844 436941 496908
rect 436875 496843 436941 496844
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 437514 475174 438134 498000
rect 438350 496909 438410 499530
rect 438534 497045 438594 499530
rect 438531 497044 438597 497045
rect 438531 496980 438532 497044
rect 438596 496980 438597 497044
rect 438531 496979 438597 496980
rect 439454 496909 439514 499530
rect 440558 499530 440732 499590
rect 441080 499590 441140 500106
rect 441760 499590 441820 500106
rect 442848 499590 442908 500106
rect 443528 499590 443588 500106
rect 443936 499590 443996 500106
rect 445296 499590 445356 500106
rect 445976 499590 446036 500106
rect 446384 499590 446444 500106
rect 447608 499590 447668 500106
rect 448288 499590 448348 500106
rect 448696 499590 448756 500106
rect 449784 499590 449844 500106
rect 451008 499590 451068 500106
rect 441080 499530 441170 499590
rect 441760 499530 442090 499590
rect 440558 496909 440618 499530
rect 441110 498133 441170 499530
rect 441107 498132 441173 498133
rect 441107 498068 441108 498132
rect 441172 498068 441173 498132
rect 441107 498067 441173 498068
rect 438347 496908 438413 496909
rect 438347 496844 438348 496908
rect 438412 496844 438413 496908
rect 438347 496843 438413 496844
rect 439451 496908 439517 496909
rect 439451 496844 439452 496908
rect 439516 496844 439517 496908
rect 439451 496843 439517 496844
rect 440555 496908 440621 496909
rect 440555 496844 440556 496908
rect 440620 496844 440621 496908
rect 440555 496843 440621 496844
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 412000 438134 438618
rect 441234 478894 441854 498000
rect 442030 496909 442090 499530
rect 442766 499530 442908 499590
rect 443502 499530 443588 499590
rect 443870 499530 443996 499590
rect 444790 499530 445356 499590
rect 445894 499530 446036 499590
rect 446262 499530 446444 499590
rect 447550 499530 447668 499590
rect 448286 499530 448348 499590
rect 448654 499530 448756 499590
rect 449758 499530 449844 499590
rect 450862 499530 451068 499590
rect 442766 497045 442826 499530
rect 442763 497044 442829 497045
rect 442763 496980 442764 497044
rect 442828 496980 442829 497044
rect 442763 496979 442829 496980
rect 443502 496909 443562 499530
rect 443870 497045 443930 499530
rect 443867 497044 443933 497045
rect 443867 496980 443868 497044
rect 443932 496980 443933 497044
rect 443867 496979 443933 496980
rect 444790 496909 444850 499530
rect 442027 496908 442093 496909
rect 442027 496844 442028 496908
rect 442092 496844 442093 496908
rect 442027 496843 442093 496844
rect 443499 496908 443565 496909
rect 443499 496844 443500 496908
rect 443564 496844 443565 496908
rect 443499 496843 443565 496844
rect 444787 496908 444853 496909
rect 444787 496844 444788 496908
rect 444852 496844 444853 496908
rect 444787 496843 444853 496844
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 412000 441854 442338
rect 444954 482614 445574 498000
rect 445894 496909 445954 499530
rect 446262 497045 446322 499530
rect 446259 497044 446325 497045
rect 446259 496980 446260 497044
rect 446324 496980 446325 497044
rect 446259 496979 446325 496980
rect 447550 496909 447610 499530
rect 448286 497045 448346 499530
rect 448283 497044 448349 497045
rect 448283 496980 448284 497044
rect 448348 496980 448349 497044
rect 448283 496979 448349 496980
rect 448654 496909 448714 499530
rect 449758 497045 449818 499530
rect 449755 497044 449821 497045
rect 449755 496980 449756 497044
rect 449820 496980 449821 497044
rect 449755 496979 449821 496980
rect 450862 496909 450922 499530
rect 451144 498810 451204 500106
rect 452232 499590 452292 500106
rect 453320 499590 453380 500106
rect 452232 499530 452578 499590
rect 451046 498750 451204 498810
rect 451046 497045 451106 498750
rect 451043 497044 451109 497045
rect 451043 496980 451044 497044
rect 451108 496980 451109 497044
rect 451043 496979 451109 496980
rect 445891 496908 445957 496909
rect 445891 496844 445892 496908
rect 445956 496844 445957 496908
rect 445891 496843 445957 496844
rect 447547 496908 447613 496909
rect 447547 496844 447548 496908
rect 447612 496844 447613 496908
rect 447547 496843 447613 496844
rect 448651 496908 448717 496909
rect 448651 496844 448652 496908
rect 448716 496844 448717 496908
rect 448651 496843 448717 496844
rect 450859 496908 450925 496909
rect 450859 496844 450860 496908
rect 450924 496844 450925 496908
rect 450859 496843 450925 496844
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 412000 445574 446058
rect 451794 489454 452414 498000
rect 452518 496909 452578 499530
rect 453254 499530 453380 499590
rect 453592 499590 453652 500106
rect 454408 499590 454468 500106
rect 455768 499590 455828 500106
rect 453592 499530 453682 499590
rect 453254 496909 453314 499530
rect 453622 497045 453682 499530
rect 454358 499530 454468 499590
rect 455646 499530 455828 499590
rect 456040 499590 456100 500106
rect 456992 499590 457052 500106
rect 458080 499590 458140 500106
rect 458488 499590 458548 500106
rect 459168 499590 459228 500106
rect 456040 499530 456258 499590
rect 453619 497044 453685 497045
rect 453619 496980 453620 497044
rect 453684 496980 453685 497044
rect 453619 496979 453685 496980
rect 454358 496909 454418 499530
rect 455646 498269 455706 499530
rect 455643 498268 455709 498269
rect 455643 498204 455644 498268
rect 455708 498204 455709 498268
rect 455643 498203 455709 498204
rect 456198 498133 456258 499530
rect 456934 499530 457052 499590
rect 458038 499530 458140 499590
rect 458406 499530 458548 499590
rect 458958 499530 459228 499590
rect 460936 499590 460996 500106
rect 463520 499590 463580 500106
rect 465968 499590 466028 500106
rect 468280 499590 468340 500106
rect 471000 499590 471060 500106
rect 473448 499590 473508 500106
rect 475896 499590 475956 500106
rect 478480 499590 478540 500106
rect 480928 499590 480988 500106
rect 483512 499590 483572 500106
rect 460936 499530 461042 499590
rect 463520 499530 463618 499590
rect 456195 498132 456261 498133
rect 456195 498068 456196 498132
rect 456260 498068 456261 498132
rect 456195 498067 456261 498068
rect 452515 496908 452581 496909
rect 452515 496844 452516 496908
rect 452580 496844 452581 496908
rect 452515 496843 452581 496844
rect 453251 496908 453317 496909
rect 453251 496844 453252 496908
rect 453316 496844 453317 496908
rect 453251 496843 453317 496844
rect 454355 496908 454421 496909
rect 454355 496844 454356 496908
rect 454420 496844 454421 496908
rect 454355 496843 454421 496844
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 412000 452414 416898
rect 455514 493174 456134 498000
rect 456934 496909 456994 499530
rect 458038 497317 458098 499530
rect 458035 497316 458101 497317
rect 458035 497252 458036 497316
rect 458100 497252 458101 497316
rect 458035 497251 458101 497252
rect 458406 496909 458466 499530
rect 458958 497045 459018 499530
rect 458955 497044 459021 497045
rect 458955 496980 458956 497044
rect 459020 496980 459021 497044
rect 458955 496979 459021 496980
rect 456931 496908 456997 496909
rect 456931 496844 456932 496908
rect 456996 496844 456997 496908
rect 456931 496843 456997 496844
rect 458403 496908 458469 496909
rect 458403 496844 458404 496908
rect 458468 496844 458469 496908
rect 458403 496843 458469 496844
rect 459234 496894 459854 498000
rect 460982 496909 461042 499530
rect 463558 498269 463618 499530
rect 465950 499530 466028 499590
rect 468158 499530 468340 499590
rect 470918 499530 471060 499590
rect 473310 499530 473508 499590
rect 475886 499530 475956 499590
rect 478462 499530 478540 499590
rect 480670 499530 480988 499590
rect 483430 499530 483572 499590
rect 485960 499590 486020 500106
rect 488544 499590 488604 500106
rect 490992 499590 491052 500106
rect 493440 499590 493500 500106
rect 485960 499530 486066 499590
rect 488544 499530 488642 499590
rect 463555 498268 463621 498269
rect 463555 498204 463556 498268
rect 463620 498204 463621 498268
rect 463555 498203 463621 498204
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 412000 456134 420618
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 460979 496908 461045 496909
rect 460979 496844 460980 496908
rect 461044 496844 461045 496908
rect 460979 496843 461045 496844
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 412000 459854 424338
rect 462954 464614 463574 498000
rect 465950 496909 466010 499530
rect 468158 496909 468218 499530
rect 465947 496908 466013 496909
rect 465947 496844 465948 496908
rect 466012 496844 466013 496908
rect 465947 496843 466013 496844
rect 468155 496908 468221 496909
rect 468155 496844 468156 496908
rect 468220 496844 468221 496908
rect 468155 496843 468221 496844
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 412000 463574 428058
rect 469794 471454 470414 498000
rect 470918 496909 470978 499530
rect 473310 496909 473370 499530
rect 470915 496908 470981 496909
rect 470915 496844 470916 496908
rect 470980 496844 470981 496908
rect 470915 496843 470981 496844
rect 473307 496908 473373 496909
rect 473307 496844 473308 496908
rect 473372 496844 473373 496908
rect 473307 496843 473373 496844
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 412000 470414 434898
rect 473514 475174 474134 498000
rect 475886 496909 475946 499530
rect 475883 496908 475949 496909
rect 475883 496844 475884 496908
rect 475948 496844 475949 496908
rect 475883 496843 475949 496844
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 412000 474134 438618
rect 477234 478894 477854 498000
rect 478462 496909 478522 499530
rect 480670 496909 480730 499530
rect 478459 496908 478525 496909
rect 478459 496844 478460 496908
rect 478524 496844 478525 496908
rect 478459 496843 478525 496844
rect 480667 496908 480733 496909
rect 480667 496844 480668 496908
rect 480732 496844 480733 496908
rect 480667 496843 480733 496844
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 412000 477854 442338
rect 480954 482614 481574 498000
rect 483430 496909 483490 499530
rect 486006 496909 486066 499530
rect 483427 496908 483493 496909
rect 483427 496844 483428 496908
rect 483492 496844 483493 496908
rect 483427 496843 483493 496844
rect 486003 496908 486069 496909
rect 486003 496844 486004 496908
rect 486068 496844 486069 496908
rect 486003 496843 486069 496844
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 412000 481574 446058
rect 487794 489454 488414 498000
rect 488582 496909 488642 499530
rect 490974 499530 491052 499590
rect 493366 499530 493500 499590
rect 495888 499590 495948 500106
rect 498472 499590 498532 500106
rect 500920 499590 500980 500106
rect 503368 499590 503428 500106
rect 505952 499590 506012 500106
rect 495888 499530 496002 499590
rect 498472 499530 498578 499590
rect 490974 496909 491034 499530
rect 488579 496908 488645 496909
rect 488579 496844 488580 496908
rect 488644 496844 488645 496908
rect 488579 496843 488645 496844
rect 490971 496908 491037 496909
rect 490971 496844 490972 496908
rect 491036 496844 491037 496908
rect 490971 496843 491037 496844
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 412000 488414 416898
rect 491514 493174 492134 498000
rect 493366 496909 493426 499530
rect 493363 496908 493429 496909
rect 493363 496844 493364 496908
rect 493428 496844 493429 496908
rect 493363 496843 493429 496844
rect 495234 496894 495854 498000
rect 495942 496909 496002 499530
rect 498518 497045 498578 499530
rect 500910 499530 500980 499590
rect 503302 499530 503428 499590
rect 505510 499530 506012 499590
rect 498515 497044 498581 497045
rect 498515 496980 498516 497044
rect 498580 496980 498581 497044
rect 498515 496979 498581 496980
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 412000 492134 420618
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495939 496908 496005 496909
rect 495939 496844 495940 496908
rect 496004 496844 496005 496908
rect 495939 496843 496005 496844
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 412000 495854 424338
rect 498954 464614 499574 498000
rect 500910 496909 500970 499530
rect 503302 496909 503362 499530
rect 505510 496909 505570 499530
rect 500907 496908 500973 496909
rect 500907 496844 500908 496908
rect 500972 496844 500973 496908
rect 500907 496843 500973 496844
rect 503299 496908 503365 496909
rect 503299 496844 503300 496908
rect 503364 496844 503365 496908
rect 503299 496843 503365 496844
rect 505507 496908 505573 496909
rect 505507 496844 505508 496908
rect 505572 496844 505573 496908
rect 505507 496843 505573 496844
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 412000 499574 428058
rect 505794 471454 506414 498000
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 412000 506414 434898
rect 509514 475174 510134 498000
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 412000 510134 438618
rect 513234 478894 513854 498000
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 412000 513854 442338
rect 516954 482614 517574 498000
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 412000 517574 446058
rect 523794 489454 524414 498000
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 412000 524414 416898
rect 527514 493174 528134 498000
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 412000 528134 420618
rect 531234 496894 531854 498000
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 412000 531854 424338
rect 534954 464614 535574 498000
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 412000 535574 428058
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 412000 542414 434898
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 412000 546134 438618
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 412000 549854 442338
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 444208 399454 444528 399486
rect 444208 399218 444250 399454
rect 444486 399218 444528 399454
rect 444208 399134 444528 399218
rect 444208 398898 444250 399134
rect 444486 398898 444528 399134
rect 444208 398866 444528 398898
rect 474928 399454 475248 399486
rect 474928 399218 474970 399454
rect 475206 399218 475248 399454
rect 474928 399134 475248 399218
rect 474928 398898 474970 399134
rect 475206 398898 475248 399134
rect 474928 398866 475248 398898
rect 505648 399454 505968 399486
rect 505648 399218 505690 399454
rect 505926 399218 505968 399454
rect 505648 399134 505968 399218
rect 505648 398898 505690 399134
rect 505926 398898 505968 399134
rect 505648 398866 505968 398898
rect 536368 399454 536688 399486
rect 536368 399218 536410 399454
rect 536646 399218 536688 399454
rect 536368 399134 536688 399218
rect 536368 398898 536410 399134
rect 536646 398898 536688 399134
rect 536368 398866 536688 398898
rect 459568 381454 459888 381486
rect 459568 381218 459610 381454
rect 459846 381218 459888 381454
rect 459568 381134 459888 381218
rect 459568 380898 459610 381134
rect 459846 380898 459888 381134
rect 459568 380866 459888 380898
rect 490288 381454 490608 381486
rect 490288 381218 490330 381454
rect 490566 381218 490608 381454
rect 490288 381134 490608 381218
rect 490288 380898 490330 381134
rect 490566 380898 490608 381134
rect 490288 380866 490608 380898
rect 521008 381454 521328 381486
rect 521008 381218 521050 381454
rect 521286 381218 521328 381454
rect 521008 381134 521328 381218
rect 521008 380898 521050 381134
rect 521286 380898 521328 381134
rect 521008 380866 521328 380898
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 444208 363454 444528 363486
rect 444208 363218 444250 363454
rect 444486 363218 444528 363454
rect 444208 363134 444528 363218
rect 444208 362898 444250 363134
rect 444486 362898 444528 363134
rect 444208 362866 444528 362898
rect 474928 363454 475248 363486
rect 474928 363218 474970 363454
rect 475206 363218 475248 363454
rect 474928 363134 475248 363218
rect 474928 362898 474970 363134
rect 475206 362898 475248 363134
rect 474928 362866 475248 362898
rect 505648 363454 505968 363486
rect 505648 363218 505690 363454
rect 505926 363218 505968 363454
rect 505648 363134 505968 363218
rect 505648 362898 505690 363134
rect 505926 362898 505968 363134
rect 505648 362866 505968 362898
rect 536368 363454 536688 363486
rect 536368 363218 536410 363454
rect 536646 363218 536688 363454
rect 536368 363134 536688 363218
rect 536368 362898 536410 363134
rect 536646 362898 536688 363134
rect 536368 362866 536688 362898
rect 459568 345454 459888 345486
rect 459568 345218 459610 345454
rect 459846 345218 459888 345454
rect 459568 345134 459888 345218
rect 459568 344898 459610 345134
rect 459846 344898 459888 345134
rect 459568 344866 459888 344898
rect 490288 345454 490608 345486
rect 490288 345218 490330 345454
rect 490566 345218 490608 345454
rect 490288 345134 490608 345218
rect 490288 344898 490330 345134
rect 490566 344898 490608 345134
rect 490288 344866 490608 344898
rect 521008 345454 521328 345486
rect 521008 345218 521050 345454
rect 521286 345218 521328 345454
rect 521008 345134 521328 345218
rect 521008 344898 521050 345134
rect 521286 344898 521328 345134
rect 521008 344866 521328 344898
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 444208 327454 444528 327486
rect 444208 327218 444250 327454
rect 444486 327218 444528 327454
rect 444208 327134 444528 327218
rect 444208 326898 444250 327134
rect 444486 326898 444528 327134
rect 444208 326866 444528 326898
rect 474928 327454 475248 327486
rect 474928 327218 474970 327454
rect 475206 327218 475248 327454
rect 474928 327134 475248 327218
rect 474928 326898 474970 327134
rect 475206 326898 475248 327134
rect 474928 326866 475248 326898
rect 505648 327454 505968 327486
rect 505648 327218 505690 327454
rect 505926 327218 505968 327454
rect 505648 327134 505968 327218
rect 505648 326898 505690 327134
rect 505926 326898 505968 327134
rect 505648 326866 505968 326898
rect 536368 327454 536688 327486
rect 536368 327218 536410 327454
rect 536646 327218 536688 327454
rect 536368 327134 536688 327218
rect 536368 326898 536410 327134
rect 536646 326898 536688 327134
rect 536368 326866 536688 326898
rect 459568 309454 459888 309486
rect 459568 309218 459610 309454
rect 459846 309218 459888 309454
rect 459568 309134 459888 309218
rect 459568 308898 459610 309134
rect 459846 308898 459888 309134
rect 459568 308866 459888 308898
rect 490288 309454 490608 309486
rect 490288 309218 490330 309454
rect 490566 309218 490608 309454
rect 490288 309134 490608 309218
rect 490288 308898 490330 309134
rect 490566 308898 490608 309134
rect 490288 308866 490608 308898
rect 521008 309454 521328 309486
rect 521008 309218 521050 309454
rect 521286 309218 521328 309454
rect 521008 309134 521328 309218
rect 521008 308898 521050 309134
rect 521286 308898 521328 309134
rect 521008 308866 521328 308898
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 142000 434414 146898
rect 437514 295174 438134 298000
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 142000 438134 150618
rect 441234 262894 441854 298000
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 142000 441854 154338
rect 444954 266614 445574 298000
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 142000 445574 158058
rect 451794 273454 452414 298000
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 142000 452414 164898
rect 455514 277174 456134 298000
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 142000 456134 168618
rect 459234 280894 459854 298000
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 142000 459854 172338
rect 462954 284614 463574 298000
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 142000 463574 176058
rect 469794 291454 470414 298000
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 142000 470414 146898
rect 473514 295174 474134 298000
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 142000 474134 150618
rect 477234 262894 477854 298000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 142000 477854 154338
rect 480954 266614 481574 298000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 142000 481574 158058
rect 487794 273454 488414 298000
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 142000 488414 164898
rect 491514 277174 492134 298000
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 142000 492134 168618
rect 495234 280894 495854 298000
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 142000 495854 172338
rect 498954 284614 499574 298000
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 142000 499574 176058
rect 505794 291454 506414 298000
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 142000 506414 146898
rect 509514 295174 510134 298000
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 142000 510134 150618
rect 513234 262894 513854 298000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 399707 139500 399773 139501
rect 399707 139436 399708 139500
rect 399772 139436 399773 139500
rect 399707 139435 399773 139436
rect 419568 129454 419888 129486
rect 419568 129218 419610 129454
rect 419846 129218 419888 129454
rect 419568 129134 419888 129218
rect 419568 128898 419610 129134
rect 419846 128898 419888 129134
rect 419568 128866 419888 128898
rect 450288 129454 450608 129486
rect 450288 129218 450330 129454
rect 450566 129218 450608 129454
rect 450288 129134 450608 129218
rect 450288 128898 450330 129134
rect 450566 128898 450608 129134
rect 450288 128866 450608 128898
rect 481008 129454 481328 129486
rect 481008 129218 481050 129454
rect 481286 129218 481328 129454
rect 481008 129134 481328 129218
rect 481008 128898 481050 129134
rect 481286 128898 481328 129134
rect 481008 128866 481328 128898
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 404208 111454 404528 111486
rect 404208 111218 404250 111454
rect 404486 111218 404528 111454
rect 404208 111134 404528 111218
rect 404208 110898 404250 111134
rect 404486 110898 404528 111134
rect 404208 110866 404528 110898
rect 434928 111454 435248 111486
rect 434928 111218 434970 111454
rect 435206 111218 435248 111454
rect 434928 111134 435248 111218
rect 434928 110898 434970 111134
rect 435206 110898 435248 111134
rect 434928 110866 435248 110898
rect 465648 111454 465968 111486
rect 465648 111218 465690 111454
rect 465926 111218 465968 111454
rect 465648 111134 465968 111218
rect 465648 110898 465690 111134
rect 465926 110898 465968 111134
rect 465648 110866 465968 110898
rect 496368 111454 496688 111486
rect 496368 111218 496410 111454
rect 496646 111218 496688 111454
rect 496368 111134 496688 111218
rect 496368 110898 496410 111134
rect 496646 110898 496688 111134
rect 496368 110866 496688 110898
rect 419568 93454 419888 93486
rect 419568 93218 419610 93454
rect 419846 93218 419888 93454
rect 419568 93134 419888 93218
rect 419568 92898 419610 93134
rect 419846 92898 419888 93134
rect 419568 92866 419888 92898
rect 450288 93454 450608 93486
rect 450288 93218 450330 93454
rect 450566 93218 450608 93454
rect 450288 93134 450608 93218
rect 450288 92898 450330 93134
rect 450566 92898 450608 93134
rect 450288 92866 450608 92898
rect 481008 93454 481328 93486
rect 481008 93218 481050 93454
rect 481286 93218 481328 93454
rect 481008 93134 481328 93218
rect 481008 92898 481050 93134
rect 481286 92898 481328 93134
rect 481008 92866 481328 92898
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 404208 75454 404528 75486
rect 404208 75218 404250 75454
rect 404486 75218 404528 75454
rect 404208 75134 404528 75218
rect 404208 74898 404250 75134
rect 404486 74898 404528 75134
rect 404208 74866 404528 74898
rect 434928 75454 435248 75486
rect 434928 75218 434970 75454
rect 435206 75218 435248 75454
rect 434928 75134 435248 75218
rect 434928 74898 434970 75134
rect 435206 74898 435248 75134
rect 434928 74866 435248 74898
rect 465648 75454 465968 75486
rect 465648 75218 465690 75454
rect 465926 75218 465968 75454
rect 465648 75134 465968 75218
rect 465648 74898 465690 75134
rect 465926 74898 465968 75134
rect 465648 74866 465968 74898
rect 496368 75454 496688 75486
rect 496368 75218 496410 75454
rect 496646 75218 496688 75454
rect 496368 75134 496688 75218
rect 496368 74898 496410 75134
rect 496646 74898 496688 75134
rect 496368 74866 496688 74898
rect 419568 57454 419888 57486
rect 419568 57218 419610 57454
rect 419846 57218 419888 57454
rect 419568 57134 419888 57218
rect 419568 56898 419610 57134
rect 419846 56898 419888 57134
rect 419568 56866 419888 56898
rect 450288 57454 450608 57486
rect 450288 57218 450330 57454
rect 450566 57218 450608 57454
rect 450288 57134 450608 57218
rect 450288 56898 450330 57134
rect 450566 56898 450608 57134
rect 450288 56866 450608 56898
rect 481008 57454 481328 57486
rect 481008 57218 481050 57454
rect 481286 57218 481328 57454
rect 481008 57134 481328 57218
rect 481008 56898 481050 57134
rect 481286 56898 481328 57134
rect 481008 56866 481328 56898
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 404208 39454 404528 39486
rect 404208 39218 404250 39454
rect 404486 39218 404528 39454
rect 404208 39134 404528 39218
rect 404208 38898 404250 39134
rect 404486 38898 404528 39134
rect 404208 38866 404528 38898
rect 434928 39454 435248 39486
rect 434928 39218 434970 39454
rect 435206 39218 435248 39454
rect 434928 39134 435248 39218
rect 434928 38898 434970 39134
rect 435206 38898 435248 39134
rect 434928 38866 435248 38898
rect 465648 39454 465968 39486
rect 465648 39218 465690 39454
rect 465926 39218 465968 39454
rect 465648 39134 465968 39218
rect 465648 38898 465690 39134
rect 465926 38898 465968 39134
rect 465648 38866 465968 38898
rect 496368 39454 496688 39486
rect 496368 39218 496410 39454
rect 496646 39218 496688 39454
rect 496368 39134 496688 39218
rect 496368 38898 496410 39134
rect 496646 38898 496688 39134
rect 496368 38866 496688 38898
rect 399523 28524 399589 28525
rect 399523 28460 399524 28524
rect 399588 28460 399589 28524
rect 399523 28459 399589 28460
rect 399339 28388 399405 28389
rect 399339 28324 399340 28388
rect 399404 28324 399405 28388
rect 399339 28323 399405 28324
rect 397502 28190 397746 28250
rect 397502 27573 397562 28190
rect 397499 27572 397565 27573
rect 397499 27508 397500 27572
rect 397564 27508 397565 27572
rect 397499 27507 397565 27508
rect 397794 3454 398414 28000
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 7174 402134 28000
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 10894 405854 28000
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 14614 409574 28000
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 28000
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 28000
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 28000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 28000
rect 433794 3454 434414 28000
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 7174 438134 28000
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 10894 441854 28000
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 14614 445574 28000
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 21454 452414 28000
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 28000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 28000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 28000
rect 469794 3454 470414 28000
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 7174 474134 28000
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 10894 477854 28000
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 14614 481574 28000
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 21454 488414 28000
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 28000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 28000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 28000
rect 505794 3454 506414 28000
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 7174 510134 28000
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 266614 517574 298000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 273454 524414 298000
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 277174 528134 298000
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 280894 531854 298000
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 284614 535574 298000
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 291454 542414 298000
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 295174 546134 298000
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 262894 549854 298000
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 51008 579218 51244 579454
rect 51008 578898 51244 579134
rect 185376 579218 185612 579454
rect 185376 578898 185612 579134
rect 50328 561218 50564 561454
rect 50328 560898 50564 561134
rect 186056 561218 186292 561454
rect 186056 560898 186292 561134
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 51008 543218 51244 543454
rect 51008 542898 51244 543134
rect 185376 543218 185612 543454
rect 185376 542898 185612 543134
rect 50328 525218 50564 525454
rect 50328 524898 50564 525134
rect 186056 525218 186292 525454
rect 186056 524898 186292 525134
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 51008 507218 51244 507454
rect 51008 506898 51244 507134
rect 185376 507218 185612 507454
rect 185376 506898 185612 507134
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 66986 428378 67222 428614
rect 67306 428378 67542 428614
rect 66986 428058 67222 428294
rect 67306 428058 67542 428294
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 91826 417218 92062 417454
rect 92146 417218 92382 417454
rect 91826 416898 92062 417134
rect 92146 416898 92382 417134
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 95546 420938 95782 421174
rect 95866 420938 96102 421174
rect 95546 420618 95782 420854
rect 95866 420618 96102 420854
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 99266 424658 99502 424894
rect 99586 424658 99822 424894
rect 99266 424338 99502 424574
rect 99586 424338 99822 424574
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 102986 428378 103222 428614
rect 103306 428378 103542 428614
rect 102986 428058 103222 428294
rect 103306 428058 103542 428294
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 109826 435218 110062 435454
rect 110146 435218 110382 435454
rect 109826 434898 110062 435134
rect 110146 434898 110382 435134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 49610 381218 49846 381454
rect 49610 380898 49846 381134
rect 80330 381218 80566 381454
rect 80330 380898 80566 381134
rect 111050 381218 111286 381454
rect 111050 380898 111286 381134
rect 34250 363218 34486 363454
rect 34250 362898 34486 363134
rect 64970 363218 65206 363454
rect 64970 362898 65206 363134
rect 95690 363218 95926 363454
rect 95690 362898 95926 363134
rect 126410 363218 126646 363454
rect 126410 362898 126646 363134
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 49610 345218 49846 345454
rect 49610 344898 49846 345134
rect 80330 345218 80566 345454
rect 80330 344898 80566 345134
rect 111050 345218 111286 345454
rect 111050 344898 111286 345134
rect 34250 327218 34486 327454
rect 34250 326898 34486 327134
rect 64970 327218 65206 327454
rect 64970 326898 65206 327134
rect 95690 327218 95926 327454
rect 95690 326898 95926 327134
rect 126410 327218 126646 327454
rect 126410 326898 126646 327134
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 49610 309218 49846 309454
rect 49610 308898 49846 309134
rect 80330 309218 80566 309454
rect 80330 308898 80566 309134
rect 111050 309218 111286 309454
rect 111050 308898 111286 309134
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 176378 67222 176614
rect 67306 176378 67542 176614
rect 66986 176058 67222 176294
rect 67306 176058 67542 176294
rect 66986 140378 67222 140614
rect 67306 140378 67542 140614
rect 66986 140058 67222 140294
rect 67306 140058 67542 140294
rect 66986 104378 67222 104614
rect 67306 104378 67542 104614
rect 66986 104058 67222 104294
rect 67306 104058 67542 104294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 84986 122378 85222 122614
rect 85306 122378 85542 122614
rect 84986 122058 85222 122294
rect 85306 122058 85542 122294
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 91826 165218 92062 165454
rect 92146 165218 92382 165454
rect 91826 164898 92062 165134
rect 92146 164898 92382 165134
rect 91826 129218 92062 129454
rect 92146 129218 92382 129454
rect 91826 128898 92062 129134
rect 92146 128898 92382 129134
rect 91826 93218 92062 93454
rect 92146 93218 92382 93454
rect 91826 92898 92062 93134
rect 92146 92898 92382 93134
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 95546 168938 95782 169174
rect 95866 168938 96102 169174
rect 95546 168618 95782 168854
rect 95866 168618 96102 168854
rect 95546 132938 95782 133174
rect 95866 132938 96102 133174
rect 95546 132618 95782 132854
rect 95866 132618 96102 132854
rect 95546 96938 95782 97174
rect 95866 96938 96102 97174
rect 95546 96618 95782 96854
rect 95866 96618 96102 96854
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 99266 172658 99502 172894
rect 99586 172658 99822 172894
rect 99266 172338 99502 172574
rect 99586 172338 99822 172574
rect 99266 136658 99502 136894
rect 99586 136658 99822 136894
rect 99266 136338 99502 136574
rect 99586 136338 99822 136574
rect 99266 100658 99502 100894
rect 99586 100658 99822 100894
rect 99266 100338 99502 100574
rect 99586 100338 99822 100574
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 102986 176378 103222 176614
rect 103306 176378 103542 176614
rect 102986 176058 103222 176294
rect 103306 176058 103542 176294
rect 102986 140378 103222 140614
rect 103306 140378 103542 140614
rect 102986 140058 103222 140294
rect 103306 140058 103542 140294
rect 102986 104378 103222 104614
rect 103306 104378 103542 104614
rect 102986 104058 103222 104294
rect 103306 104058 103542 104294
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 127826 165218 128062 165454
rect 128146 165218 128382 165454
rect 127826 164898 128062 165134
rect 128146 164898 128382 165134
rect 127826 129218 128062 129454
rect 128146 129218 128382 129454
rect 127826 128898 128062 129134
rect 128146 128898 128382 129134
rect 127826 93218 128062 93454
rect 128146 93218 128382 93454
rect 127826 92898 128062 93134
rect 128146 92898 128382 93134
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 131546 168938 131782 169174
rect 131866 168938 132102 169174
rect 131546 168618 131782 168854
rect 131866 168618 132102 168854
rect 131546 132938 131782 133174
rect 131866 132938 132102 133174
rect 131546 132618 131782 132854
rect 131866 132618 132102 132854
rect 131546 96938 131782 97174
rect 131866 96938 132102 97174
rect 131546 96618 131782 96854
rect 131866 96618 132102 96854
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 135266 172658 135502 172894
rect 135586 172658 135822 172894
rect 135266 172338 135502 172574
rect 135586 172338 135822 172574
rect 135266 136658 135502 136894
rect 135586 136658 135822 136894
rect 135266 136338 135502 136574
rect 135586 136338 135822 136574
rect 135266 100658 135502 100894
rect 135586 100658 135822 100894
rect 135266 100338 135502 100574
rect 135586 100338 135822 100574
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 138986 176378 139222 176614
rect 139306 176378 139542 176614
rect 138986 176058 139222 176294
rect 139306 176058 139542 176294
rect 138986 140378 139222 140614
rect 139306 140378 139542 140614
rect 138986 140058 139222 140294
rect 139306 140058 139542 140294
rect 138986 104378 139222 104614
rect 139306 104378 139542 104614
rect 138986 104058 139222 104294
rect 139306 104058 139542 104294
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 163826 165218 164062 165454
rect 164146 165218 164382 165454
rect 163826 164898 164062 165134
rect 164146 164898 164382 165134
rect 163826 129218 164062 129454
rect 164146 129218 164382 129454
rect 163826 128898 164062 129134
rect 164146 128898 164382 129134
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 163826 93218 164062 93454
rect 164146 93218 164382 93454
rect 163826 92898 164062 93134
rect 164146 92898 164382 93134
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 401008 579218 401244 579454
rect 401008 578898 401244 579134
rect 535376 579218 535612 579454
rect 535376 578898 535612 579134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 400328 561218 400564 561454
rect 400328 560898 400564 561134
rect 536056 561218 536292 561454
rect 536056 560898 536292 561134
rect 401008 543218 401244 543454
rect 401008 542898 401244 543134
rect 535376 543218 535612 543454
rect 535376 542898 535612 543134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 400328 525218 400564 525454
rect 400328 524898 400564 525134
rect 536056 525218 536292 525454
rect 536056 524898 536292 525134
rect 401008 507218 401244 507454
rect 401008 506898 401244 507134
rect 535376 507218 535612 507454
rect 535376 506898 535612 507134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 209610 417218 209846 417454
rect 209610 416898 209846 417134
rect 240330 417218 240566 417454
rect 240330 416898 240566 417134
rect 271050 417218 271286 417454
rect 271050 416898 271286 417134
rect 301770 417218 302006 417454
rect 301770 416898 302006 417134
rect 332490 417218 332726 417454
rect 332490 416898 332726 417134
rect 363210 417218 363446 417454
rect 363210 416898 363446 417134
rect 393930 417218 394166 417454
rect 393930 416898 394166 417134
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 194250 399218 194486 399454
rect 194250 398898 194486 399134
rect 224970 399218 225206 399454
rect 224970 398898 225206 399134
rect 255690 399218 255926 399454
rect 255690 398898 255926 399134
rect 286410 399218 286646 399454
rect 286410 398898 286646 399134
rect 317130 399218 317366 399454
rect 317130 398898 317366 399134
rect 347850 399218 348086 399454
rect 347850 398898 348086 399134
rect 378570 399218 378806 399454
rect 378570 398898 378806 399134
rect 209610 381218 209846 381454
rect 209610 380898 209846 381134
rect 240330 381218 240566 381454
rect 240330 380898 240566 381134
rect 271050 381218 271286 381454
rect 271050 380898 271286 381134
rect 301770 381218 302006 381454
rect 301770 380898 302006 381134
rect 332490 381218 332726 381454
rect 332490 380898 332726 381134
rect 363210 381218 363446 381454
rect 363210 380898 363446 381134
rect 393930 381218 394166 381454
rect 393930 380898 394166 381134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 194250 363218 194486 363454
rect 194250 362898 194486 363134
rect 224970 363218 225206 363454
rect 224970 362898 225206 363134
rect 255690 363218 255926 363454
rect 255690 362898 255926 363134
rect 286410 363218 286646 363454
rect 286410 362898 286646 363134
rect 317130 363218 317366 363454
rect 317130 362898 317366 363134
rect 347850 363218 348086 363454
rect 347850 362898 348086 363134
rect 378570 363218 378806 363454
rect 378570 362898 378806 363134
rect 209610 345218 209846 345454
rect 209610 344898 209846 345134
rect 240330 345218 240566 345454
rect 240330 344898 240566 345134
rect 271050 345218 271286 345454
rect 271050 344898 271286 345134
rect 301770 345218 302006 345454
rect 301770 344898 302006 345134
rect 332490 345218 332726 345454
rect 332490 344898 332726 345134
rect 363210 345218 363446 345454
rect 363210 344898 363446 345134
rect 393930 345218 394166 345454
rect 393930 344898 394166 345134
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 194250 327218 194486 327454
rect 194250 326898 194486 327134
rect 224970 327218 225206 327454
rect 224970 326898 225206 327134
rect 255690 327218 255926 327454
rect 255690 326898 255926 327134
rect 286410 327218 286646 327454
rect 286410 326898 286646 327134
rect 317130 327218 317366 327454
rect 317130 326898 317366 327134
rect 347850 327218 348086 327454
rect 347850 326898 348086 327134
rect 378570 327218 378806 327454
rect 378570 326898 378806 327134
rect 209610 309218 209846 309454
rect 209610 308898 209846 309134
rect 240330 309218 240566 309454
rect 240330 308898 240566 309134
rect 271050 309218 271286 309454
rect 271050 308898 271286 309134
rect 301770 309218 302006 309454
rect 301770 308898 302006 309134
rect 332490 309218 332726 309454
rect 332490 308898 332726 309134
rect 363210 309218 363446 309454
rect 363210 308898 363446 309134
rect 393930 309218 394166 309454
rect 393930 308898 394166 309134
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 194250 291218 194486 291454
rect 194250 290898 194486 291134
rect 224970 291218 225206 291454
rect 224970 290898 225206 291134
rect 255690 291218 255926 291454
rect 255690 290898 255926 291134
rect 286410 291218 286646 291454
rect 286410 290898 286646 291134
rect 317130 291218 317366 291454
rect 317130 290898 317366 291134
rect 347850 291218 348086 291454
rect 347850 290898 348086 291134
rect 378570 291218 378806 291454
rect 378570 290898 378806 291134
rect 209610 273218 209846 273454
rect 209610 272898 209846 273134
rect 240330 273218 240566 273454
rect 240330 272898 240566 273134
rect 271050 273218 271286 273454
rect 271050 272898 271286 273134
rect 301770 273218 302006 273454
rect 301770 272898 302006 273134
rect 332490 273218 332726 273454
rect 332490 272898 332726 273134
rect 363210 273218 363446 273454
rect 363210 272898 363446 273134
rect 393930 273218 394166 273454
rect 393930 272898 394166 273134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 194250 255218 194486 255454
rect 194250 254898 194486 255134
rect 224970 255218 225206 255454
rect 224970 254898 225206 255134
rect 255690 255218 255926 255454
rect 255690 254898 255926 255134
rect 286410 255218 286646 255454
rect 286410 254898 286646 255134
rect 317130 255218 317366 255454
rect 317130 254898 317366 255134
rect 347850 255218 348086 255454
rect 347850 254898 348086 255134
rect 378570 255218 378806 255454
rect 378570 254898 378806 255134
rect 209610 237218 209846 237454
rect 209610 236898 209846 237134
rect 240330 237218 240566 237454
rect 240330 236898 240566 237134
rect 271050 237218 271286 237454
rect 271050 236898 271286 237134
rect 301770 237218 302006 237454
rect 301770 236898 302006 237134
rect 332490 237218 332726 237454
rect 332490 236898 332726 237134
rect 363210 237218 363446 237454
rect 363210 236898 363446 237134
rect 393930 237218 394166 237454
rect 393930 236898 394166 237134
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 194250 219218 194486 219454
rect 194250 218898 194486 219134
rect 224970 219218 225206 219454
rect 224970 218898 225206 219134
rect 255690 219218 255926 219454
rect 255690 218898 255926 219134
rect 286410 219218 286646 219454
rect 286410 218898 286646 219134
rect 317130 219218 317366 219454
rect 317130 218898 317366 219134
rect 347850 219218 348086 219454
rect 347850 218898 348086 219134
rect 378570 219218 378806 219454
rect 378570 218898 378806 219134
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 189610 129218 189846 129454
rect 189610 128898 189846 129134
rect 220330 129218 220566 129454
rect 220330 128898 220566 129134
rect 251050 129218 251286 129454
rect 251050 128898 251286 129134
rect 174250 111218 174486 111454
rect 174250 110898 174486 111134
rect 204970 111218 205206 111454
rect 204970 110898 205206 111134
rect 235690 111218 235926 111454
rect 235690 110898 235926 111134
rect 266410 111218 266646 111454
rect 266410 110898 266646 111134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 189610 93218 189846 93454
rect 189610 92898 189846 93134
rect 220330 93218 220566 93454
rect 220330 92898 220566 93134
rect 251050 93218 251286 93454
rect 251050 92898 251286 93134
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 174250 75218 174486 75454
rect 174250 74898 174486 75134
rect 204970 75218 205206 75454
rect 204970 74898 205206 75134
rect 235690 75218 235926 75454
rect 235690 74898 235926 75134
rect 266410 75218 266646 75454
rect 266410 74898 266646 75134
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 189610 57218 189846 57454
rect 189610 56898 189846 57134
rect 220330 57218 220566 57454
rect 220330 56898 220566 57134
rect 251050 57218 251286 57454
rect 251050 56898 251286 57134
rect 174250 39218 174486 39454
rect 174250 38898 174486 39134
rect 204970 39218 205206 39454
rect 204970 38898 205206 39134
rect 235690 39218 235926 39454
rect 235690 38898 235926 39134
rect 266410 39218 266646 39454
rect 266410 38898 266646 39134
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 444250 399218 444486 399454
rect 444250 398898 444486 399134
rect 474970 399218 475206 399454
rect 474970 398898 475206 399134
rect 505690 399218 505926 399454
rect 505690 398898 505926 399134
rect 536410 399218 536646 399454
rect 536410 398898 536646 399134
rect 459610 381218 459846 381454
rect 459610 380898 459846 381134
rect 490330 381218 490566 381454
rect 490330 380898 490566 381134
rect 521050 381218 521286 381454
rect 521050 380898 521286 381134
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 444250 363218 444486 363454
rect 444250 362898 444486 363134
rect 474970 363218 475206 363454
rect 474970 362898 475206 363134
rect 505690 363218 505926 363454
rect 505690 362898 505926 363134
rect 536410 363218 536646 363454
rect 536410 362898 536646 363134
rect 459610 345218 459846 345454
rect 459610 344898 459846 345134
rect 490330 345218 490566 345454
rect 490330 344898 490566 345134
rect 521050 345218 521286 345454
rect 521050 344898 521286 345134
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 444250 327218 444486 327454
rect 444250 326898 444486 327134
rect 474970 327218 475206 327454
rect 474970 326898 475206 327134
rect 505690 327218 505926 327454
rect 505690 326898 505926 327134
rect 536410 327218 536646 327454
rect 536410 326898 536646 327134
rect 459610 309218 459846 309454
rect 459610 308898 459846 309134
rect 490330 309218 490566 309454
rect 490330 308898 490566 309134
rect 521050 309218 521286 309454
rect 521050 308898 521286 309134
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 419610 129218 419846 129454
rect 419610 128898 419846 129134
rect 450330 129218 450566 129454
rect 450330 128898 450566 129134
rect 481050 129218 481286 129454
rect 481050 128898 481286 129134
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 404250 111218 404486 111454
rect 404250 110898 404486 111134
rect 434970 111218 435206 111454
rect 434970 110898 435206 111134
rect 465690 111218 465926 111454
rect 465690 110898 465926 111134
rect 496410 111218 496646 111454
rect 496410 110898 496646 111134
rect 419610 93218 419846 93454
rect 419610 92898 419846 93134
rect 450330 93218 450566 93454
rect 450330 92898 450566 93134
rect 481050 93218 481286 93454
rect 481050 92898 481286 93134
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 404250 75218 404486 75454
rect 404250 74898 404486 75134
rect 434970 75218 435206 75454
rect 434970 74898 435206 75134
rect 465690 75218 465926 75454
rect 465690 74898 465926 75134
rect 496410 75218 496646 75454
rect 496410 74898 496646 75134
rect 419610 57218 419846 57454
rect 419610 56898 419846 57134
rect 450330 57218 450566 57454
rect 450330 56898 450566 57134
rect 481050 57218 481286 57454
rect 481050 56898 481286 57134
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 404250 39218 404486 39454
rect 404250 38898 404486 39134
rect 434970 39218 435206 39454
rect 434970 38898 435206 39134
rect 465690 39218 465926 39454
rect 465690 38898 465926 39134
rect 496410 39218 496646 39454
rect 496410 38898 496646 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 51008 579454
rect 51244 579218 185376 579454
rect 185612 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 401008 579454
rect 401244 579218 535376 579454
rect 535612 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 51008 579134
rect 51244 578898 185376 579134
rect 185612 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 401008 579134
rect 401244 578898 535376 579134
rect 535612 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 50328 561454
rect 50564 561218 186056 561454
rect 186292 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 400328 561454
rect 400564 561218 536056 561454
rect 536292 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 50328 561134
rect 50564 560898 186056 561134
rect 186292 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 400328 561134
rect 400564 560898 536056 561134
rect 536292 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 51008 543454
rect 51244 543218 185376 543454
rect 185612 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 401008 543454
rect 401244 543218 535376 543454
rect 535612 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 51008 543134
rect 51244 542898 185376 543134
rect 185612 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 401008 543134
rect 401244 542898 535376 543134
rect 535612 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 50328 525454
rect 50564 525218 186056 525454
rect 186292 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 400328 525454
rect 400564 525218 536056 525454
rect 536292 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 50328 525134
rect 50564 524898 186056 525134
rect 186292 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 400328 525134
rect 400564 524898 536056 525134
rect 536292 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 51008 507454
rect 51244 507218 185376 507454
rect 185612 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 401008 507454
rect 401244 507218 535376 507454
rect 535612 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 51008 507134
rect 51244 506898 185376 507134
rect 185612 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 401008 507134
rect 401244 506898 535376 507134
rect 535612 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 109826 435454
rect 110062 435218 110146 435454
rect 110382 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 109826 435134
rect 110062 434898 110146 435134
rect 110382 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 66986 428614
rect 67222 428378 67306 428614
rect 67542 428378 102986 428614
rect 103222 428378 103306 428614
rect 103542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 66986 428294
rect 67222 428058 67306 428294
rect 67542 428058 102986 428294
rect 103222 428058 103306 428294
rect 103542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 99266 424894
rect 99502 424658 99586 424894
rect 99822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 99266 424574
rect 99502 424338 99586 424574
rect 99822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 95546 421174
rect 95782 420938 95866 421174
rect 96102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 95546 420854
rect 95782 420618 95866 420854
rect 96102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 91826 417454
rect 92062 417218 92146 417454
rect 92382 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 209610 417454
rect 209846 417218 240330 417454
rect 240566 417218 271050 417454
rect 271286 417218 301770 417454
rect 302006 417218 332490 417454
rect 332726 417218 363210 417454
rect 363446 417218 393930 417454
rect 394166 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 91826 417134
rect 92062 416898 92146 417134
rect 92382 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 209610 417134
rect 209846 416898 240330 417134
rect 240566 416898 271050 417134
rect 271286 416898 301770 417134
rect 302006 416898 332490 417134
rect 332726 416898 363210 417134
rect 363446 416898 393930 417134
rect 394166 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 194250 399454
rect 194486 399218 224970 399454
rect 225206 399218 255690 399454
rect 255926 399218 286410 399454
rect 286646 399218 317130 399454
rect 317366 399218 347850 399454
rect 348086 399218 378570 399454
rect 378806 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 444250 399454
rect 444486 399218 474970 399454
rect 475206 399218 505690 399454
rect 505926 399218 536410 399454
rect 536646 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 194250 399134
rect 194486 398898 224970 399134
rect 225206 398898 255690 399134
rect 255926 398898 286410 399134
rect 286646 398898 317130 399134
rect 317366 398898 347850 399134
rect 348086 398898 378570 399134
rect 378806 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 444250 399134
rect 444486 398898 474970 399134
rect 475206 398898 505690 399134
rect 505926 398898 536410 399134
rect 536646 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 49610 381454
rect 49846 381218 80330 381454
rect 80566 381218 111050 381454
rect 111286 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 209610 381454
rect 209846 381218 240330 381454
rect 240566 381218 271050 381454
rect 271286 381218 301770 381454
rect 302006 381218 332490 381454
rect 332726 381218 363210 381454
rect 363446 381218 393930 381454
rect 394166 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 459610 381454
rect 459846 381218 490330 381454
rect 490566 381218 521050 381454
rect 521286 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 49610 381134
rect 49846 380898 80330 381134
rect 80566 380898 111050 381134
rect 111286 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 209610 381134
rect 209846 380898 240330 381134
rect 240566 380898 271050 381134
rect 271286 380898 301770 381134
rect 302006 380898 332490 381134
rect 332726 380898 363210 381134
rect 363446 380898 393930 381134
rect 394166 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 459610 381134
rect 459846 380898 490330 381134
rect 490566 380898 521050 381134
rect 521286 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 34250 363454
rect 34486 363218 64970 363454
rect 65206 363218 95690 363454
rect 95926 363218 126410 363454
rect 126646 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 194250 363454
rect 194486 363218 224970 363454
rect 225206 363218 255690 363454
rect 255926 363218 286410 363454
rect 286646 363218 317130 363454
rect 317366 363218 347850 363454
rect 348086 363218 378570 363454
rect 378806 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 444250 363454
rect 444486 363218 474970 363454
rect 475206 363218 505690 363454
rect 505926 363218 536410 363454
rect 536646 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 34250 363134
rect 34486 362898 64970 363134
rect 65206 362898 95690 363134
rect 95926 362898 126410 363134
rect 126646 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 194250 363134
rect 194486 362898 224970 363134
rect 225206 362898 255690 363134
rect 255926 362898 286410 363134
rect 286646 362898 317130 363134
rect 317366 362898 347850 363134
rect 348086 362898 378570 363134
rect 378806 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 444250 363134
rect 444486 362898 474970 363134
rect 475206 362898 505690 363134
rect 505926 362898 536410 363134
rect 536646 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 49610 345454
rect 49846 345218 80330 345454
rect 80566 345218 111050 345454
rect 111286 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 209610 345454
rect 209846 345218 240330 345454
rect 240566 345218 271050 345454
rect 271286 345218 301770 345454
rect 302006 345218 332490 345454
rect 332726 345218 363210 345454
rect 363446 345218 393930 345454
rect 394166 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 459610 345454
rect 459846 345218 490330 345454
rect 490566 345218 521050 345454
rect 521286 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 49610 345134
rect 49846 344898 80330 345134
rect 80566 344898 111050 345134
rect 111286 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 209610 345134
rect 209846 344898 240330 345134
rect 240566 344898 271050 345134
rect 271286 344898 301770 345134
rect 302006 344898 332490 345134
rect 332726 344898 363210 345134
rect 363446 344898 393930 345134
rect 394166 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 459610 345134
rect 459846 344898 490330 345134
rect 490566 344898 521050 345134
rect 521286 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 34250 327454
rect 34486 327218 64970 327454
rect 65206 327218 95690 327454
rect 95926 327218 126410 327454
rect 126646 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 194250 327454
rect 194486 327218 224970 327454
rect 225206 327218 255690 327454
rect 255926 327218 286410 327454
rect 286646 327218 317130 327454
rect 317366 327218 347850 327454
rect 348086 327218 378570 327454
rect 378806 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 444250 327454
rect 444486 327218 474970 327454
rect 475206 327218 505690 327454
rect 505926 327218 536410 327454
rect 536646 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 34250 327134
rect 34486 326898 64970 327134
rect 65206 326898 95690 327134
rect 95926 326898 126410 327134
rect 126646 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 194250 327134
rect 194486 326898 224970 327134
rect 225206 326898 255690 327134
rect 255926 326898 286410 327134
rect 286646 326898 317130 327134
rect 317366 326898 347850 327134
rect 348086 326898 378570 327134
rect 378806 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 444250 327134
rect 444486 326898 474970 327134
rect 475206 326898 505690 327134
rect 505926 326898 536410 327134
rect 536646 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 49610 309454
rect 49846 309218 80330 309454
rect 80566 309218 111050 309454
rect 111286 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 209610 309454
rect 209846 309218 240330 309454
rect 240566 309218 271050 309454
rect 271286 309218 301770 309454
rect 302006 309218 332490 309454
rect 332726 309218 363210 309454
rect 363446 309218 393930 309454
rect 394166 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 459610 309454
rect 459846 309218 490330 309454
rect 490566 309218 521050 309454
rect 521286 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 49610 309134
rect 49846 308898 80330 309134
rect 80566 308898 111050 309134
rect 111286 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 209610 309134
rect 209846 308898 240330 309134
rect 240566 308898 271050 309134
rect 271286 308898 301770 309134
rect 302006 308898 332490 309134
rect 332726 308898 363210 309134
rect 363446 308898 393930 309134
rect 394166 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 459610 309134
rect 459846 308898 490330 309134
rect 490566 308898 521050 309134
rect 521286 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 194250 291454
rect 194486 291218 224970 291454
rect 225206 291218 255690 291454
rect 255926 291218 286410 291454
rect 286646 291218 317130 291454
rect 317366 291218 347850 291454
rect 348086 291218 378570 291454
rect 378806 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 194250 291134
rect 194486 290898 224970 291134
rect 225206 290898 255690 291134
rect 255926 290898 286410 291134
rect 286646 290898 317130 291134
rect 317366 290898 347850 291134
rect 348086 290898 378570 291134
rect 378806 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 209610 273454
rect 209846 273218 240330 273454
rect 240566 273218 271050 273454
rect 271286 273218 301770 273454
rect 302006 273218 332490 273454
rect 332726 273218 363210 273454
rect 363446 273218 393930 273454
rect 394166 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 209610 273134
rect 209846 272898 240330 273134
rect 240566 272898 271050 273134
rect 271286 272898 301770 273134
rect 302006 272898 332490 273134
rect 332726 272898 363210 273134
rect 363446 272898 393930 273134
rect 394166 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 194250 255454
rect 194486 255218 224970 255454
rect 225206 255218 255690 255454
rect 255926 255218 286410 255454
rect 286646 255218 317130 255454
rect 317366 255218 347850 255454
rect 348086 255218 378570 255454
rect 378806 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 194250 255134
rect 194486 254898 224970 255134
rect 225206 254898 255690 255134
rect 255926 254898 286410 255134
rect 286646 254898 317130 255134
rect 317366 254898 347850 255134
rect 348086 254898 378570 255134
rect 378806 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 209610 237454
rect 209846 237218 240330 237454
rect 240566 237218 271050 237454
rect 271286 237218 301770 237454
rect 302006 237218 332490 237454
rect 332726 237218 363210 237454
rect 363446 237218 393930 237454
rect 394166 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 209610 237134
rect 209846 236898 240330 237134
rect 240566 236898 271050 237134
rect 271286 236898 301770 237134
rect 302006 236898 332490 237134
rect 332726 236898 363210 237134
rect 363446 236898 393930 237134
rect 394166 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 194250 219454
rect 194486 219218 224970 219454
rect 225206 219218 255690 219454
rect 255926 219218 286410 219454
rect 286646 219218 317130 219454
rect 317366 219218 347850 219454
rect 348086 219218 378570 219454
rect 378806 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 194250 219134
rect 194486 218898 224970 219134
rect 225206 218898 255690 219134
rect 255926 218898 286410 219134
rect 286646 218898 317130 219134
rect 317366 218898 347850 219134
rect 348086 218898 378570 219134
rect 378806 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 66986 176614
rect 67222 176378 67306 176614
rect 67542 176378 102986 176614
rect 103222 176378 103306 176614
rect 103542 176378 138986 176614
rect 139222 176378 139306 176614
rect 139542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 66986 176294
rect 67222 176058 67306 176294
rect 67542 176058 102986 176294
rect 103222 176058 103306 176294
rect 103542 176058 138986 176294
rect 139222 176058 139306 176294
rect 139542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 99266 172894
rect 99502 172658 99586 172894
rect 99822 172658 135266 172894
rect 135502 172658 135586 172894
rect 135822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 99266 172574
rect 99502 172338 99586 172574
rect 99822 172338 135266 172574
rect 135502 172338 135586 172574
rect 135822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 95546 169174
rect 95782 168938 95866 169174
rect 96102 168938 131546 169174
rect 131782 168938 131866 169174
rect 132102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 95546 168854
rect 95782 168618 95866 168854
rect 96102 168618 131546 168854
rect 131782 168618 131866 168854
rect 132102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 91826 165454
rect 92062 165218 92146 165454
rect 92382 165218 127826 165454
rect 128062 165218 128146 165454
rect 128382 165218 163826 165454
rect 164062 165218 164146 165454
rect 164382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 91826 165134
rect 92062 164898 92146 165134
rect 92382 164898 127826 165134
rect 128062 164898 128146 165134
rect 128382 164898 163826 165134
rect 164062 164898 164146 165134
rect 164382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 66986 140614
rect 67222 140378 67306 140614
rect 67542 140378 102986 140614
rect 103222 140378 103306 140614
rect 103542 140378 138986 140614
rect 139222 140378 139306 140614
rect 139542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 66986 140294
rect 67222 140058 67306 140294
rect 67542 140058 102986 140294
rect 103222 140058 103306 140294
rect 103542 140058 138986 140294
rect 139222 140058 139306 140294
rect 139542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 99266 136894
rect 99502 136658 99586 136894
rect 99822 136658 135266 136894
rect 135502 136658 135586 136894
rect 135822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 99266 136574
rect 99502 136338 99586 136574
rect 99822 136338 135266 136574
rect 135502 136338 135586 136574
rect 135822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 95546 133174
rect 95782 132938 95866 133174
rect 96102 132938 131546 133174
rect 131782 132938 131866 133174
rect 132102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 95546 132854
rect 95782 132618 95866 132854
rect 96102 132618 131546 132854
rect 131782 132618 131866 132854
rect 132102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 91826 129454
rect 92062 129218 92146 129454
rect 92382 129218 127826 129454
rect 128062 129218 128146 129454
rect 128382 129218 163826 129454
rect 164062 129218 164146 129454
rect 164382 129218 189610 129454
rect 189846 129218 220330 129454
rect 220566 129218 251050 129454
rect 251286 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 419610 129454
rect 419846 129218 450330 129454
rect 450566 129218 481050 129454
rect 481286 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 91826 129134
rect 92062 128898 92146 129134
rect 92382 128898 127826 129134
rect 128062 128898 128146 129134
rect 128382 128898 163826 129134
rect 164062 128898 164146 129134
rect 164382 128898 189610 129134
rect 189846 128898 220330 129134
rect 220566 128898 251050 129134
rect 251286 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 419610 129134
rect 419846 128898 450330 129134
rect 450566 128898 481050 129134
rect 481286 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 84986 122614
rect 85222 122378 85306 122614
rect 85542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 84986 122294
rect 85222 122058 85306 122294
rect 85542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 174250 111454
rect 174486 111218 204970 111454
rect 205206 111218 235690 111454
rect 235926 111218 266410 111454
rect 266646 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 404250 111454
rect 404486 111218 434970 111454
rect 435206 111218 465690 111454
rect 465926 111218 496410 111454
rect 496646 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 174250 111134
rect 174486 110898 204970 111134
rect 205206 110898 235690 111134
rect 235926 110898 266410 111134
rect 266646 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 404250 111134
rect 404486 110898 434970 111134
rect 435206 110898 465690 111134
rect 465926 110898 496410 111134
rect 496646 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 66986 104614
rect 67222 104378 67306 104614
rect 67542 104378 102986 104614
rect 103222 104378 103306 104614
rect 103542 104378 138986 104614
rect 139222 104378 139306 104614
rect 139542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 66986 104294
rect 67222 104058 67306 104294
rect 67542 104058 102986 104294
rect 103222 104058 103306 104294
rect 103542 104058 138986 104294
rect 139222 104058 139306 104294
rect 139542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 99266 100894
rect 99502 100658 99586 100894
rect 99822 100658 135266 100894
rect 135502 100658 135586 100894
rect 135822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 99266 100574
rect 99502 100338 99586 100574
rect 99822 100338 135266 100574
rect 135502 100338 135586 100574
rect 135822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 95546 97174
rect 95782 96938 95866 97174
rect 96102 96938 131546 97174
rect 131782 96938 131866 97174
rect 132102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 95546 96854
rect 95782 96618 95866 96854
rect 96102 96618 131546 96854
rect 131782 96618 131866 96854
rect 132102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 91826 93454
rect 92062 93218 92146 93454
rect 92382 93218 127826 93454
rect 128062 93218 128146 93454
rect 128382 93218 163826 93454
rect 164062 93218 164146 93454
rect 164382 93218 189610 93454
rect 189846 93218 220330 93454
rect 220566 93218 251050 93454
rect 251286 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 419610 93454
rect 419846 93218 450330 93454
rect 450566 93218 481050 93454
rect 481286 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 91826 93134
rect 92062 92898 92146 93134
rect 92382 92898 127826 93134
rect 128062 92898 128146 93134
rect 128382 92898 163826 93134
rect 164062 92898 164146 93134
rect 164382 92898 189610 93134
rect 189846 92898 220330 93134
rect 220566 92898 251050 93134
rect 251286 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 419610 93134
rect 419846 92898 450330 93134
rect 450566 92898 481050 93134
rect 481286 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 174250 75454
rect 174486 75218 204970 75454
rect 205206 75218 235690 75454
rect 235926 75218 266410 75454
rect 266646 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 404250 75454
rect 404486 75218 434970 75454
rect 435206 75218 465690 75454
rect 465926 75218 496410 75454
rect 496646 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 174250 75134
rect 174486 74898 204970 75134
rect 205206 74898 235690 75134
rect 235926 74898 266410 75134
rect 266646 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 404250 75134
rect 404486 74898 434970 75134
rect 435206 74898 465690 75134
rect 465926 74898 496410 75134
rect 496646 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 189610 57454
rect 189846 57218 220330 57454
rect 220566 57218 251050 57454
rect 251286 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 419610 57454
rect 419846 57218 450330 57454
rect 450566 57218 481050 57454
rect 481286 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 189610 57134
rect 189846 56898 220330 57134
rect 220566 56898 251050 57134
rect 251286 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 419610 57134
rect 419846 56898 450330 57134
rect 450566 56898 481050 57134
rect 481286 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 174250 39454
rect 174486 39218 204970 39454
rect 205206 39218 235690 39454
rect 235926 39218 266410 39454
rect 266646 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 404250 39454
rect 404486 39218 434970 39454
rect 435206 39218 465690 39454
rect 465926 39218 496410 39454
rect 496646 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 174250 39134
rect 174486 38898 204970 39134
rect 205206 38898 235690 39134
rect 235926 38898 266410 39134
rect 266646 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 404250 39134
rect 404486 38898 434970 39134
rect 435206 38898 465690 39134
rect 465926 38898 496410 39134
rect 496646 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Core  core
timestamp 0
transform 1 0 30000 0 1 300000
box 0 0 100000 100000
use sky130_sram_2kbyte_1rw1r_32x512_8  dmem
timestamp 0
transform 1 0 400000 0 1 500000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  imem
timestamp 0
transform 1 0 50000 0 1 500000
box 0 0 136620 83308
use Motor_Top  m1
timestamp 0
transform 1 0 440000 0 1 300000
box 0 0 110000 110000
use Motor_Top  m2
timestamp 0
transform 1 0 170000 0 1 30000
box 0 0 110000 110000
use Motor_Top  m3
timestamp 0
transform 1 0 400000 0 1 30000
box 0 0 110000 110000
use WB_InterConnect  wb_inter_connect
timestamp 0
transform 1 0 190000 0 1 200000
box 0 0 220000 220000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 28000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 142000 218414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 142000 254414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 142000 398414 198000 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 142000 470414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 142000 506414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 298000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 402000 74414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 402000 110414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 142000 182414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 422000 398414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 142000 434414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 412000 470414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 412000 506414 498000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 402000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 585308 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 585308 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 585308 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 585308 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 422000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 422000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 422000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 422000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 422000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 585308 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 585308 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 585308 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 585308 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 412000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 28000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 142000 222134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 142000 258134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 142000 402134 198000 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 142000 438134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 142000 474134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 142000 510134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 298000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 402000 78134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 402000 114134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 142000 186134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 422000 402134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 412000 438134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 412000 474134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 412000 510134 498000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 402000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 585308 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 585308 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 585308 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 585308 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 422000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 422000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 422000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 422000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 422000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 585308 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 585308 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 585308 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 585308 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 412000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 28000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 142000 189854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 142000 225854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 142000 261854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 142000 405854 198000 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 142000 441854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 142000 477854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 298000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 402000 81854 498000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 402000 117854 498000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 498000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 422000 405854 498000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 412000 441854 498000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 412000 477854 498000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 412000 513854 498000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 402000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 585308 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 585308 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 585308 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 422000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 422000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 422000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 422000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 422000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 422000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 585308 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 585308 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 585308 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 585308 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 412000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 28000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 142000 193574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 142000 229574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 142000 265574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 142000 409574 198000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 142000 445574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 142000 481574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 298000 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 402000 49574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 402000 85574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 402000 121574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 422000 409574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 412000 445574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 412000 481574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 412000 517574 498000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 585308 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 585308 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 585308 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 585308 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 422000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 422000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 422000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 422000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 422000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 422000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 585308 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 585308 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 585308 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 585308 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 28000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 142000 207854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 142000 243854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 142000 279854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 198000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 142000 459854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 142000 495854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 298000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 402000 63854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 402000 99854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 142000 171854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 142000 423854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 412000 459854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 412000 495854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 412000 531854 498000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 585308 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 585308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 585308 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 585308 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 422000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 422000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 422000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 422000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 422000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 422000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 585308 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 585308 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 585308 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 585308 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 28000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 142000 211574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 142000 247574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 198000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 142000 463574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 142000 499574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 298000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 402000 67574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 402000 103574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 142000 175574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 142000 427574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 412000 463574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 412000 499574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 412000 535574 498000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 402000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 585308 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 585308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 585308 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 585308 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 422000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 422000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 422000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 422000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 422000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 422000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 585308 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 585308 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 585308 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 585308 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 28000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 142000 200414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 142000 236414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 142000 272414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 198000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 142000 452414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 142000 488414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 298000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 402000 56414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 402000 92414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 402000 128414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 142000 416414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 412000 452414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 412000 488414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 412000 524414 498000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 585308 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 585308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 585308 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 585308 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 422000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 422000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 422000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 422000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 422000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 422000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 585308 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 585308 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 585308 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 585308 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 28000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 142000 204134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 142000 240134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 142000 276134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 198000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 142000 456134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 142000 492134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 298000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 402000 60134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 402000 96134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 402000 132134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 142000 168134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 142000 420134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 412000 456134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 412000 492134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 412000 528134 498000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 585308 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 585308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 585308 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 585308 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 422000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 422000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 422000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 422000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 422000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 422000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 585308 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 585308 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 585308 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 585308 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
