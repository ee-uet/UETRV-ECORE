VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Motor_Top
  CLASS BLOCK ;
  FOREIGN Motor_Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 500.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 0.000 9.110 4.000 ;
    END
  END clock
  PIN io_ba_match
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 10.920 500.000 11.520 ;
    END
  END io_ba_match
  PIN io_motor_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END io_motor_irq
  PIN io_pwm_high
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 496.000 14.170 500.000 ;
    END
  END io_pwm_high
  PIN io_pwm_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 496.000 41.770 500.000 ;
    END
  END io_pwm_low
  PIN io_qei_ch_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 33.360 500.000 33.960 ;
    END
  END io_qei_ch_a
  PIN io_qei_ch_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END io_qei_ch_b
  PIN io_wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END io_wbs_ack_o
  PIN io_wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 496.000 69.370 500.000 ;
    END
  END io_wbs_data_o[0]
  PIN io_wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 496.000 291.550 500.000 ;
    END
  END io_wbs_data_o[10]
  PIN io_wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END io_wbs_data_o[11]
  PIN io_wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_wbs_data_o[12]
  PIN io_wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END io_wbs_data_o[13]
  PIN io_wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 328.480 500.000 329.080 ;
    END
  END io_wbs_data_o[14]
  PIN io_wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 374.040 500.000 374.640 ;
    END
  END io_wbs_data_o[15]
  PIN io_wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END io_wbs_data_o[16]
  PIN io_wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 230.560 4.000 231.160 ;
    END
  END io_wbs_data_o[17]
  PIN io_wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END io_wbs_data_o[18]
  PIN io_wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END io_wbs_data_o[19]
  PIN io_wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END io_wbs_data_o[1]
  PIN io_wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 396.480 500.000 397.080 ;
    END
  END io_wbs_data_o[20]
  PIN io_wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END io_wbs_data_o[21]
  PIN io_wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 496.000 402.870 500.000 ;
    END
  END io_wbs_data_o[22]
  PIN io_wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 419.600 500.000 420.200 ;
    END
  END io_wbs_data_o[23]
  PIN io_wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 465.160 500.000 465.760 ;
    END
  END io_wbs_data_o[24]
  PIN io_wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END io_wbs_data_o[25]
  PIN io_wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END io_wbs_data_o[26]
  PIN io_wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END io_wbs_data_o[27]
  PIN io_wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END io_wbs_data_o[28]
  PIN io_wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END io_wbs_data_o[29]
  PIN io_wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 146.920 500.000 147.520 ;
    END
  END io_wbs_data_o[2]
  PIN io_wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END io_wbs_data_o[30]
  PIN io_wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 496.000 486.130 500.000 ;
    END
  END io_wbs_data_o[31]
  PIN io_wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END io_wbs_data_o[3]
  PIN io_wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END io_wbs_data_o[4]
  PIN io_wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 214.920 500.000 215.520 ;
    END
  END io_wbs_data_o[5]
  PIN io_wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 238.040 500.000 238.640 ;
    END
  END io_wbs_data_o[6]
  PIN io_wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END io_wbs_data_o[7]
  PIN io_wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 496.000 236.350 500.000 ;
    END
  END io_wbs_data_o[8]
  PIN io_wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 260.480 500.000 261.080 ;
    END
  END io_wbs_data_o[9]
  PIN io_wbs_m2s_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 55.800 500.000 56.400 ;
    END
  END io_wbs_m2s_addr[0]
  PIN io_wbs_m2s_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 282.920 500.000 283.520 ;
    END
  END io_wbs_m2s_addr[10]
  PIN io_wbs_m2s_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END io_wbs_m2s_addr[11]
  PIN io_wbs_m2s_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 496.000 319.610 500.000 ;
    END
  END io_wbs_m2s_addr[12]
  PIN io_wbs_m2s_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 306.040 500.000 306.640 ;
    END
  END io_wbs_m2s_addr[13]
  PIN io_wbs_m2s_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END io_wbs_m2s_addr[14]
  PIN io_wbs_m2s_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 496.000 347.210 500.000 ;
    END
  END io_wbs_m2s_addr[15]
  PIN io_wbs_m2s_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 101.360 500.000 101.960 ;
    END
  END io_wbs_m2s_addr[1]
  PIN io_wbs_m2s_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 169.360 500.000 169.960 ;
    END
  END io_wbs_m2s_addr[2]
  PIN io_wbs_m2s_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 192.480 500.000 193.080 ;
    END
  END io_wbs_m2s_addr[3]
  PIN io_wbs_m2s_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 496.000 152.630 500.000 ;
    END
  END io_wbs_m2s_addr[4]
  PIN io_wbs_m2s_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 496.000 180.690 500.000 ;
    END
  END io_wbs_m2s_addr[5]
  PIN io_wbs_m2s_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END io_wbs_m2s_addr[6]
  PIN io_wbs_m2s_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END io_wbs_m2s_addr[7]
  PIN io_wbs_m2s_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 496.000 263.950 500.000 ;
    END
  END io_wbs_m2s_addr[8]
  PIN io_wbs_m2s_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_wbs_m2s_addr[9]
  PIN io_wbs_m2s_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 78.920 500.000 79.520 ;
    END
  END io_wbs_m2s_data[0]
  PIN io_wbs_m2s_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END io_wbs_m2s_data[10]
  PIN io_wbs_m2s_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END io_wbs_m2s_data[11]
  PIN io_wbs_m2s_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END io_wbs_m2s_data[12]
  PIN io_wbs_m2s_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END io_wbs_m2s_data[13]
  PIN io_wbs_m2s_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 351.600 500.000 352.200 ;
    END
  END io_wbs_m2s_data[14]
  PIN io_wbs_m2s_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_wbs_m2s_data[15]
  PIN io_wbs_m2s_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END io_wbs_m2s_data[16]
  PIN io_wbs_m2s_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END io_wbs_m2s_data[17]
  PIN io_wbs_m2s_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 496.000 375.270 500.000 ;
    END
  END io_wbs_m2s_data[18]
  PIN io_wbs_m2s_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END io_wbs_m2s_data[19]
  PIN io_wbs_m2s_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 124.480 500.000 125.080 ;
    END
  END io_wbs_m2s_data[1]
  PIN io_wbs_m2s_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 286.320 4.000 286.920 ;
    END
  END io_wbs_m2s_data[20]
  PIN io_wbs_m2s_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END io_wbs_m2s_data[21]
  PIN io_wbs_m2s_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END io_wbs_m2s_data[22]
  PIN io_wbs_m2s_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 442.040 500.000 442.640 ;
    END
  END io_wbs_m2s_data[23]
  PIN io_wbs_m2s_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 496.000 430.470 500.000 ;
    END
  END io_wbs_m2s_data[24]
  PIN io_wbs_m2s_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 496.000 458.530 500.000 ;
    END
  END io_wbs_m2s_data[25]
  PIN io_wbs_m2s_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END io_wbs_m2s_data[26]
  PIN io_wbs_m2s_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END io_wbs_m2s_data[27]
  PIN io_wbs_m2s_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END io_wbs_m2s_data[28]
  PIN io_wbs_m2s_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END io_wbs_m2s_data[29]
  PIN io_wbs_m2s_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END io_wbs_m2s_data[2]
  PIN io_wbs_m2s_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 496.000 487.600 500.000 488.200 ;
    END
  END io_wbs_m2s_data[30]
  PIN io_wbs_m2s_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END io_wbs_m2s_data[31]
  PIN io_wbs_m2s_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 496.000 125.030 500.000 ;
    END
  END io_wbs_m2s_data[3]
  PIN io_wbs_m2s_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END io_wbs_m2s_data[4]
  PIN io_wbs_m2s_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 496.000 208.290 500.000 ;
    END
  END io_wbs_m2s_data[5]
  PIN io_wbs_m2s_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END io_wbs_m2s_data[6]
  PIN io_wbs_m2s_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END io_wbs_m2s_data[7]
  PIN io_wbs_m2s_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 0.000 223.010 4.000 ;
    END
  END io_wbs_m2s_data[8]
  PIN io_wbs_m2s_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END io_wbs_m2s_data[9]
  PIN io_wbs_m2s_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 496.000 97.430 500.000 ;
    END
  END io_wbs_m2s_sel[0]
  PIN io_wbs_m2s_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END io_wbs_m2s_sel[1]
  PIN io_wbs_m2s_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END io_wbs_m2s_sel[2]
  PIN io_wbs_m2s_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END io_wbs_m2s_sel[3]
  PIN io_wbs_m2s_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END io_wbs_m2s_stb
  PIN io_wbs_m2s_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END io_wbs_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 487.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 487.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 487.120 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 486.965 ;
      LAYER met1 ;
        RECT 5.520 10.640 494.040 487.120 ;
      LAYER met2 ;
        RECT 6.990 495.720 13.610 496.810 ;
        RECT 14.450 495.720 41.210 496.810 ;
        RECT 42.050 495.720 68.810 496.810 ;
        RECT 69.650 495.720 96.870 496.810 ;
        RECT 97.710 495.720 124.470 496.810 ;
        RECT 125.310 495.720 152.070 496.810 ;
        RECT 152.910 495.720 180.130 496.810 ;
        RECT 180.970 495.720 207.730 496.810 ;
        RECT 208.570 495.720 235.790 496.810 ;
        RECT 236.630 495.720 263.390 496.810 ;
        RECT 264.230 495.720 290.990 496.810 ;
        RECT 291.830 495.720 319.050 496.810 ;
        RECT 319.890 495.720 346.650 496.810 ;
        RECT 347.490 495.720 374.710 496.810 ;
        RECT 375.550 495.720 402.310 496.810 ;
        RECT 403.150 495.720 429.910 496.810 ;
        RECT 430.750 495.720 457.970 496.810 ;
        RECT 458.810 495.720 485.570 496.810 ;
        RECT 486.410 495.720 491.650 496.810 ;
        RECT 6.990 4.280 491.650 495.720 ;
        RECT 6.990 3.670 8.550 4.280 ;
        RECT 9.390 3.670 26.030 4.280 ;
        RECT 26.870 3.670 43.970 4.280 ;
        RECT 44.810 3.670 61.910 4.280 ;
        RECT 62.750 3.670 79.850 4.280 ;
        RECT 80.690 3.670 97.790 4.280 ;
        RECT 98.630 3.670 115.270 4.280 ;
        RECT 116.110 3.670 133.210 4.280 ;
        RECT 134.050 3.670 151.150 4.280 ;
        RECT 151.990 3.670 169.090 4.280 ;
        RECT 169.930 3.670 187.030 4.280 ;
        RECT 187.870 3.670 204.970 4.280 ;
        RECT 205.810 3.670 222.450 4.280 ;
        RECT 223.290 3.670 240.390 4.280 ;
        RECT 241.230 3.670 258.330 4.280 ;
        RECT 259.170 3.670 276.270 4.280 ;
        RECT 277.110 3.670 294.210 4.280 ;
        RECT 295.050 3.670 311.690 4.280 ;
        RECT 312.530 3.670 329.630 4.280 ;
        RECT 330.470 3.670 347.570 4.280 ;
        RECT 348.410 3.670 365.510 4.280 ;
        RECT 366.350 3.670 383.450 4.280 ;
        RECT 384.290 3.670 401.390 4.280 ;
        RECT 402.230 3.670 418.870 4.280 ;
        RECT 419.710 3.670 436.810 4.280 ;
        RECT 437.650 3.670 454.750 4.280 ;
        RECT 455.590 3.670 472.690 4.280 ;
        RECT 473.530 3.670 490.630 4.280 ;
        RECT 491.470 3.670 491.650 4.280 ;
      LAYER met3 ;
        RECT 4.400 489.240 496.000 490.105 ;
        RECT 4.000 488.600 496.000 489.240 ;
        RECT 4.000 487.200 495.600 488.600 ;
        RECT 4.000 472.280 496.000 487.200 ;
        RECT 4.400 470.880 496.000 472.280 ;
        RECT 4.000 466.160 496.000 470.880 ;
        RECT 4.000 464.760 495.600 466.160 ;
        RECT 4.000 453.920 496.000 464.760 ;
        RECT 4.400 452.520 496.000 453.920 ;
        RECT 4.000 443.040 496.000 452.520 ;
        RECT 4.000 441.640 495.600 443.040 ;
        RECT 4.000 435.560 496.000 441.640 ;
        RECT 4.400 434.160 496.000 435.560 ;
        RECT 4.000 420.600 496.000 434.160 ;
        RECT 4.000 419.200 495.600 420.600 ;
        RECT 4.000 416.520 496.000 419.200 ;
        RECT 4.400 415.120 496.000 416.520 ;
        RECT 4.000 398.160 496.000 415.120 ;
        RECT 4.400 397.480 496.000 398.160 ;
        RECT 4.400 396.760 495.600 397.480 ;
        RECT 4.000 396.080 495.600 396.760 ;
        RECT 4.000 379.800 496.000 396.080 ;
        RECT 4.400 378.400 496.000 379.800 ;
        RECT 4.000 375.040 496.000 378.400 ;
        RECT 4.000 373.640 495.600 375.040 ;
        RECT 4.000 361.440 496.000 373.640 ;
        RECT 4.400 360.040 496.000 361.440 ;
        RECT 4.000 352.600 496.000 360.040 ;
        RECT 4.000 351.200 495.600 352.600 ;
        RECT 4.000 343.080 496.000 351.200 ;
        RECT 4.400 341.680 496.000 343.080 ;
        RECT 4.000 329.480 496.000 341.680 ;
        RECT 4.000 328.080 495.600 329.480 ;
        RECT 4.000 324.040 496.000 328.080 ;
        RECT 4.400 322.640 496.000 324.040 ;
        RECT 4.000 307.040 496.000 322.640 ;
        RECT 4.000 305.680 495.600 307.040 ;
        RECT 4.400 305.640 495.600 305.680 ;
        RECT 4.400 304.280 496.000 305.640 ;
        RECT 4.000 287.320 496.000 304.280 ;
        RECT 4.400 285.920 496.000 287.320 ;
        RECT 4.000 283.920 496.000 285.920 ;
        RECT 4.000 282.520 495.600 283.920 ;
        RECT 4.000 268.960 496.000 282.520 ;
        RECT 4.400 267.560 496.000 268.960 ;
        RECT 4.000 261.480 496.000 267.560 ;
        RECT 4.000 260.080 495.600 261.480 ;
        RECT 4.000 249.920 496.000 260.080 ;
        RECT 4.400 248.520 496.000 249.920 ;
        RECT 4.000 239.040 496.000 248.520 ;
        RECT 4.000 237.640 495.600 239.040 ;
        RECT 4.000 231.560 496.000 237.640 ;
        RECT 4.400 230.160 496.000 231.560 ;
        RECT 4.000 215.920 496.000 230.160 ;
        RECT 4.000 214.520 495.600 215.920 ;
        RECT 4.000 213.200 496.000 214.520 ;
        RECT 4.400 211.800 496.000 213.200 ;
        RECT 4.000 194.840 496.000 211.800 ;
        RECT 4.400 193.480 496.000 194.840 ;
        RECT 4.400 193.440 495.600 193.480 ;
        RECT 4.000 192.080 495.600 193.440 ;
        RECT 4.000 176.480 496.000 192.080 ;
        RECT 4.400 175.080 496.000 176.480 ;
        RECT 4.000 170.360 496.000 175.080 ;
        RECT 4.000 168.960 495.600 170.360 ;
        RECT 4.000 157.440 496.000 168.960 ;
        RECT 4.400 156.040 496.000 157.440 ;
        RECT 4.000 147.920 496.000 156.040 ;
        RECT 4.000 146.520 495.600 147.920 ;
        RECT 4.000 139.080 496.000 146.520 ;
        RECT 4.400 137.680 496.000 139.080 ;
        RECT 4.000 125.480 496.000 137.680 ;
        RECT 4.000 124.080 495.600 125.480 ;
        RECT 4.000 120.720 496.000 124.080 ;
        RECT 4.400 119.320 496.000 120.720 ;
        RECT 4.000 102.360 496.000 119.320 ;
        RECT 4.400 100.960 495.600 102.360 ;
        RECT 4.000 83.320 496.000 100.960 ;
        RECT 4.400 81.920 496.000 83.320 ;
        RECT 4.000 79.920 496.000 81.920 ;
        RECT 4.000 78.520 495.600 79.920 ;
        RECT 4.000 64.960 496.000 78.520 ;
        RECT 4.400 63.560 496.000 64.960 ;
        RECT 4.000 56.800 496.000 63.560 ;
        RECT 4.000 55.400 495.600 56.800 ;
        RECT 4.000 46.600 496.000 55.400 ;
        RECT 4.400 45.200 496.000 46.600 ;
        RECT 4.000 34.360 496.000 45.200 ;
        RECT 4.000 32.960 495.600 34.360 ;
        RECT 4.000 28.240 496.000 32.960 ;
        RECT 4.400 26.840 496.000 28.240 ;
        RECT 4.000 11.920 496.000 26.840 ;
        RECT 4.000 10.520 495.600 11.920 ;
        RECT 4.000 9.880 496.000 10.520 ;
        RECT 4.400 9.015 496.000 9.880 ;
      LAYER met4 ;
        RECT 67.455 11.055 97.440 483.305 ;
        RECT 99.840 11.055 174.240 483.305 ;
        RECT 176.640 11.055 251.040 483.305 ;
        RECT 253.440 11.055 327.840 483.305 ;
        RECT 330.240 11.055 404.640 483.305 ;
        RECT 407.040 11.055 435.785 483.305 ;
  END
END Motor_Top
END LIBRARY

