* NGSPICE file created from Core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_4 abstract view
.subckt sky130_fd_sc_hd__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt Core clock io_dbus_addr[0] io_dbus_addr[10] io_dbus_addr[11] io_dbus_addr[12]
+ io_dbus_addr[13] io_dbus_addr[14] io_dbus_addr[15] io_dbus_addr[16] io_dbus_addr[17]
+ io_dbus_addr[18] io_dbus_addr[19] io_dbus_addr[1] io_dbus_addr[20] io_dbus_addr[21]
+ io_dbus_addr[22] io_dbus_addr[23] io_dbus_addr[24] io_dbus_addr[25] io_dbus_addr[26]
+ io_dbus_addr[27] io_dbus_addr[28] io_dbus_addr[29] io_dbus_addr[2] io_dbus_addr[30]
+ io_dbus_addr[31] io_dbus_addr[3] io_dbus_addr[4] io_dbus_addr[5] io_dbus_addr[6]
+ io_dbus_addr[7] io_dbus_addr[8] io_dbus_addr[9] io_dbus_ld_type[0] io_dbus_ld_type[1]
+ io_dbus_ld_type[2] io_dbus_rd_en io_dbus_rdata[0] io_dbus_rdata[10] io_dbus_rdata[11]
+ io_dbus_rdata[12] io_dbus_rdata[13] io_dbus_rdata[14] io_dbus_rdata[15] io_dbus_rdata[16]
+ io_dbus_rdata[17] io_dbus_rdata[18] io_dbus_rdata[19] io_dbus_rdata[1] io_dbus_rdata[20]
+ io_dbus_rdata[21] io_dbus_rdata[22] io_dbus_rdata[23] io_dbus_rdata[24] io_dbus_rdata[25]
+ io_dbus_rdata[26] io_dbus_rdata[27] io_dbus_rdata[28] io_dbus_rdata[29] io_dbus_rdata[2]
+ io_dbus_rdata[30] io_dbus_rdata[31] io_dbus_rdata[3] io_dbus_rdata[4] io_dbus_rdata[5]
+ io_dbus_rdata[6] io_dbus_rdata[7] io_dbus_rdata[8] io_dbus_rdata[9] io_dbus_st_type[0]
+ io_dbus_st_type[1] io_dbus_valid io_dbus_wdata[0] io_dbus_wdata[10] io_dbus_wdata[11]
+ io_dbus_wdata[12] io_dbus_wdata[13] io_dbus_wdata[14] io_dbus_wdata[15] io_dbus_wdata[16]
+ io_dbus_wdata[17] io_dbus_wdata[18] io_dbus_wdata[19] io_dbus_wdata[1] io_dbus_wdata[20]
+ io_dbus_wdata[21] io_dbus_wdata[22] io_dbus_wdata[23] io_dbus_wdata[24] io_dbus_wdata[25]
+ io_dbus_wdata[26] io_dbus_wdata[27] io_dbus_wdata[28] io_dbus_wdata[29] io_dbus_wdata[2]
+ io_dbus_wdata[30] io_dbus_wdata[31] io_dbus_wdata[3] io_dbus_wdata[4] io_dbus_wdata[5]
+ io_dbus_wdata[6] io_dbus_wdata[7] io_dbus_wdata[8] io_dbus_wdata[9] io_dbus_wr_en
+ io_ibus_addr[0] io_ibus_addr[10] io_ibus_addr[11] io_ibus_addr[12] io_ibus_addr[13]
+ io_ibus_addr[14] io_ibus_addr[15] io_ibus_addr[16] io_ibus_addr[17] io_ibus_addr[18]
+ io_ibus_addr[19] io_ibus_addr[1] io_ibus_addr[20] io_ibus_addr[21] io_ibus_addr[22]
+ io_ibus_addr[23] io_ibus_addr[24] io_ibus_addr[25] io_ibus_addr[26] io_ibus_addr[27]
+ io_ibus_addr[28] io_ibus_addr[29] io_ibus_addr[2] io_ibus_addr[30] io_ibus_addr[31]
+ io_ibus_addr[3] io_ibus_addr[4] io_ibus_addr[5] io_ibus_addr[6] io_ibus_addr[7]
+ io_ibus_addr[8] io_ibus_addr[9] io_ibus_inst[0] io_ibus_inst[10] io_ibus_inst[11]
+ io_ibus_inst[12] io_ibus_inst[13] io_ibus_inst[14] io_ibus_inst[15] io_ibus_inst[16]
+ io_ibus_inst[17] io_ibus_inst[18] io_ibus_inst[19] io_ibus_inst[1] io_ibus_inst[20]
+ io_ibus_inst[21] io_ibus_inst[22] io_ibus_inst[23] io_ibus_inst[24] io_ibus_inst[25]
+ io_ibus_inst[26] io_ibus_inst[27] io_ibus_inst[28] io_ibus_inst[29] io_ibus_inst[2]
+ io_ibus_inst[30] io_ibus_inst[31] io_ibus_inst[3] io_ibus_inst[4] io_ibus_inst[5]
+ io_ibus_inst[6] io_ibus_inst[7] io_ibus_inst[8] io_ibus_inst[9] io_ibus_valid io_irq_motor_irq
+ io_irq_spi_irq io_irq_uart_irq reset vccd1 vssd1
XFILLER_140_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17046__A1 _16932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__S0 _09955_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _09671_/A vssd1 vssd1 vccd1 vccd1 _09672_/A sky130_fd_sc_hd__clkbuf_4
X_18869_ _19286_/CLK _18869_/D vssd1 vssd1 vccd1 vccd1 _18869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09906__S0 _09904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11094__A1 _09477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09284__A2_N _12696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14446__A _14502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09105_ _09174_/A vssd1 vssd1 vccd1 vccd1 _09328_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10185__S _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14880__S _14882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16661__A _16806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12346__A1 _19419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17492__A _17716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _09941_/A _09935_/X _09937_/X _09740_/A vssd1 vssd1 vccd1 vccd1 _09938_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_89_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17037__A1 _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10204__S0 _09955_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09869_ _09931_/S vssd1 vssd1 vccd1 vccd1 _09930_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__A _15009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ _11900_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11903_/A sky130_fd_sc_hd__and2_2
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14120__S _14122_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12880_ _16845_/B _12560_/X _12562_/X _16431_/B _12879_/X vssd1 vssd1 vccd1 vccd1
+ _15479_/B sky130_fd_sc_hd__a221o_2
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11802_/A _11830_/X _11708_/A vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__o21a_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11045__A _19712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14550_ _14550_/A vssd1 vssd1 vccd1 vccd1 _14550_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11762_ _11762_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11788_/C sky130_fd_sc_hd__and2_1
XFILLER_14_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13501_ _13330_/X _18349_/Q _13503_/S vssd1 vssd1 vccd1 vccd1 _13502_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10832__A1 _09432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10713_ _18587_/Q _18858_/Q _19082_/Q _18826_/Q _09645_/S _09541_/A vssd1 vssd1 vccd1
+ vccd1 _10714_/B sky130_fd_sc_hd__mux4_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _13889_/X _18725_/Q _14489_/S vssd1 vssd1 vccd1 vccd1 _14482_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11693_ _15474_/A vssd1 vssd1 vccd1 vccd1 _16162_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_42_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _13586_/X _19382_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16221_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17760__A2 _17741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ _13432_/A vssd1 vssd1 vccd1 vccd1 _18320_/D sky130_fd_sc_hd__clkbuf_1
X_10644_ _10074_/X _10635_/X _10637_/Y _10643_/Y _09658_/X vssd1 vssd1 vccd1 vccd1
+ _10644_/X sky130_fd_sc_hd__o311a_4
XFILLER_155_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16151_ _16159_/C _16150_/Y _15482_/S vssd1 vssd1 vccd1 vccd1 _16151_/Y sky130_fd_sc_hd__a21oi_1
X_10575_ _10575_/A vssd1 vssd1 vccd1 vccd1 _10585_/A sky130_fd_sc_hd__clkbuf_2
X_13363_ _12861_/X _13370_/B _13362_/X _13051_/A vssd1 vssd1 vccd1 vccd1 _13363_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_158_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_127_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15102_ _15158_/A vssd1 vssd1 vccd1 vccd1 _15171_/S sky130_fd_sc_hd__buf_4
XFILLER_155_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12314_ _12314_/A _12314_/B vssd1 vssd1 vccd1 vccd1 _12314_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16082_ _12550_/X _16081_/Y _16082_/S vssd1 vssd1 vccd1 vccd1 _16082_/X sky130_fd_sc_hd__mux2_1
X_13294_ _14605_/A vssd1 vssd1 vccd1 vccd1 _13294_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16290__B _16290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15033_ _18954_/Q _15031_/X _15045_/S vssd1 vssd1 vccd1 vccd1 _15034_/A sky130_fd_sc_hd__mux2_1
X_12245_ _12245_/A vssd1 vssd1 vccd1 vccd1 _17835_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17276__A1 _17680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19841_ _19866_/CLK _19841_/D vssd1 vssd1 vccd1 vccd1 _19841_/Q sky130_fd_sc_hd__dfxtp_1
X_12176_ _19409_/Q _12176_/B vssd1 vssd1 vccd1 vccd1 _12177_/D sky130_fd_sc_hd__and2_1
XANTENNA__13419__B _13419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11127_ _18611_/Q _18946_/Q _11127_/S vssd1 vssd1 vccd1 vccd1 _11127_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10994__S1 _10934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16984_ _19647_/Q _16984_/B vssd1 vssd1 vccd1 vccd1 _16984_/X sky130_fd_sc_hd__or2_1
XFILLER_96_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19772_ _19775_/CLK _19772_/D vssd1 vssd1 vccd1 vccd1 _19772_/Q sky130_fd_sc_hd__dfxtp_1
X_18723_ _19311_/CLK _18723_/D vssd1 vssd1 vccd1 vccd1 _18723_/Q sky130_fd_sc_hd__dfxtp_1
X_15935_ _13525_/X _19301_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15936_/A sky130_fd_sc_hd__mux2_1
X_11058_ _19174_/Q _18788_/Q _19238_/Q _18357_/Q _11011_/X _11005_/X vssd1 vssd1 vccd1
+ vccd1 _11059_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13435__A _16619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10009_ _10014_/A _10009_/B vssd1 vssd1 vccd1 vccd1 _10009_/Y sky130_fd_sc_hd__nor2_1
X_18654_ _18824_/CLK _18654_/D vssd1 vssd1 vccd1 vccd1 _18654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15866_ _15866_/A vssd1 vssd1 vccd1 vccd1 _19270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17605_ _17605_/A _17605_/B vssd1 vssd1 vccd1 vccd1 _17605_/Y sky130_fd_sc_hd__nor2_1
X_14817_ _18860_/Q _13988_/X _14821_/S vssd1 vssd1 vccd1 vccd1 _14818_/A sky130_fd_sc_hd__mux2_1
X_18585_ _19081_/CLK _18585_/D vssd1 vssd1 vccd1 vccd1 _18585_/Q sky130_fd_sc_hd__dfxtp_1
X_15797_ _15797_/A vssd1 vssd1 vccd1 vccd1 _19239_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16746__A _16806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17536_ _11512_/B _17252_/X _17462_/X _17535_/Y vssd1 vssd1 vccd1 vccd1 _17536_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16539__B1 _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14748_ _14566_/X _18830_/Q _14748_/S vssd1 vssd1 vccd1 vccd1 _14749_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10284__C1 _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17467_ _17710_/S _17468_/B _17464_/X _17466_/X vssd1 vssd1 vccd1 vccd1 _17467_/X
+ sky130_fd_sc_hd__a211o_1
X_14679_ _14569_/X _18799_/Q _14687_/S vssd1 vssd1 vccd1 vccd1 _14680_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13170__A _15060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17751__A2 _17652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16418_ _19455_/Q _16415_/B _16417_/Y vssd1 vssd1 vccd1 vccd1 _19455_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19206_ _19302_/CLK _19206_/D vssd1 vssd1 vccd1 vccd1 _19206_/Q sky130_fd_sc_hd__dfxtp_1
X_17398_ _17395_/Y _17397_/Y _17572_/S vssd1 vssd1 vccd1 vccd1 _17398_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19137_ _19800_/CLK _19137_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
X_16349_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16388_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19068_ _19326_/CLK _19068_/D vssd1 vssd1 vccd1 vccd1 _19068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12328__A1 _12321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18019_ _19781_/Q _11915_/A _18027_/S vssd1 vssd1 vccd1 vccd1 _18020_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14205__S _14209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11000__A1 _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10354__A3 _10352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09723_ _10184_/A vssd1 vssd1 vccd1 vccd1 _10108_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09823__A _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10969__A _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15036__S _15045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09901__C1 _09964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09654_ _18415_/Q _18676_/Q _18575_/Q _18910_/Q _09538_/A _09547_/A vssd1 vssd1 vccd1
+ vccd1 _09654_/X sky130_fd_sc_hd__mux4_1
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09585_ _09600_/A vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12567__B2 _19345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17487__A _17731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ _19284_/Q _19122_/Q _18531_/Q _18301_/Q _09700_/A _10229_/X vssd1 vssd1 vccd1
+ vccd1 _10361_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10291_ _19318_/Q _18730_/Q _18767_/Q _18341_/Q _10260_/X _10263_/X vssd1 vssd1 vccd1
+ vccd1 _10291_/X sky130_fd_sc_hd__mux4_1
XFILLER_128_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12030_ _12030_/A vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__inv_2
XFILLER_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13954__S _13963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10976__S1 _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09733__A _09733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13981_ _14553_/A vssd1 vssd1 vccd1 vccd1 _13981_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ _15720_/A vssd1 vssd1 vccd1 vccd1 _19205_/D sky130_fd_sc_hd__clkbuf_1
X_12932_ _19629_/Q _12490_/A _12606_/Y _19559_/Q _12584_/Y vssd1 vssd1 vccd1 vccd1
+ _12932_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09594__S1 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15651_ _15708_/S vssd1 vssd1 vccd1 vccd1 _15660_/S sky130_fd_sc_hd__buf_2
XFILLER_73_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12863_ _12855_/X _12862_/X _12781_/A input26/X vssd1 vssd1 vccd1 vccd1 _15009_/A
+ sky130_fd_sc_hd__a2bb2o_2
XANTENNA__14785__S _14785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14615_/S sky130_fd_sc_hd__buf_4
X_18370_ _19315_/CLK _18370_/D vssd1 vssd1 vccd1 vccd1 _18370_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _11890_/B _12450_/B _11890_/C _18138_/A vssd1 vssd1 vccd1 vccd1 _17605_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_15582_ _15565_/X _15580_/X _15581_/Y _15549_/X _18272_/Q vssd1 vssd1 vccd1 vccd1
+ _15582_/X sky130_fd_sc_hd__a32o_2
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ _13065_/A vssd1 vssd1 vccd1 vccd1 _13144_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _12488_/B _17321_/B _17321_/C vssd1 vssd1 vccd1 vccd1 _17321_/X sky130_fd_sc_hd__and3b_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14533_ _14533_/A vssd1 vssd1 vccd1 vccd1 _18750_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _19629_/Q _19625_/Q _19620_/Q _11745_/D vssd1 vssd1 vccd1 vccd1 _11746_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17252_ _17252_/A vssd1 vssd1 vccd1 vccd1 _17252_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14464_ _14464_/A vssd1 vssd1 vccd1 vccd1 _18717_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11676_ _11676_/A _17480_/A vssd1 vssd1 vccd1 vccd1 _11730_/A sky130_fd_sc_hd__xnor2_2
XFILLER_174_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16203_ _16203_/A vssd1 vssd1 vccd1 vccd1 _19374_/D sky130_fd_sc_hd__clkbuf_1
X_13415_ _18253_/Q _13415_/B vssd1 vssd1 vccd1 vccd1 _13415_/X sky130_fd_sc_hd__or2_1
X_10627_ _10682_/A _10627_/B vssd1 vssd1 vccd1 vccd1 _10627_/Y sky130_fd_sc_hd__nor2_1
X_17183_ _17183_/A _17183_/B _17183_/C _17183_/D vssd1 vssd1 vccd1 vccd1 _17184_/B
+ sky130_fd_sc_hd__or4_1
X_14395_ _13870_/X _18687_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14396_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16134_ _16142_/C _16133_/Y _16109_/X vssd1 vssd1 vccd1 vccd1 _16134_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11230__A1 _11024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10664__S0 _10650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13346_ _12861_/X _13345_/X _12976_/A vssd1 vssd1 vccd1 vccd1 _13346_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15629__B hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10558_ _19312_/Q _18724_/Q _18761_/Q _18335_/Q _10763_/S _09590_/X vssd1 vssd1 vccd1
+ vccd1 _10559_/B sky130_fd_sc_hd__mux4_1
XFILLER_127_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16065_ _16073_/C _16065_/B vssd1 vssd1 vccd1 vccd1 _16065_/Y sky130_fd_sc_hd__nand2_1
X_13277_ _13277_/A vssd1 vssd1 vccd1 vccd1 _18308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10489_ _10485_/A _10486_/X _10488_/X vssd1 vssd1 vccd1 vccd1 _10489_/Y sky130_fd_sc_hd__o21ai_1
X_15016_ _15099_/S vssd1 vssd1 vccd1 vccd1 _15029_/S sky130_fd_sc_hd__buf_2
X_12228_ _19414_/Q _12228_/B vssd1 vssd1 vccd1 vccd1 _12271_/C sky130_fd_sc_hd__and2_1
XFILLER_69_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10967__S1 _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19824_ _19828_/CLK _19824_/D vssd1 vssd1 vccd1 vccd1 _19824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ _12159_/A _12159_/B vssd1 vssd1 vccd1 vccd1 _12209_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10741__B1 _09432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19755_ _19756_/CLK _19755_/D vssd1 vssd1 vccd1 vccd1 _19755_/Q sky130_fd_sc_hd__dfxtp_1
X_16967_ _16967_/A _16971_/B vssd1 vssd1 vccd1 vccd1 _16967_/X sky130_fd_sc_hd__or2_1
X_18706_ _19264_/CLK _18706_/D vssd1 vssd1 vccd1 vccd1 _18706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15918_ _19294_/Q _14611_/A _15920_/S vssd1 vssd1 vccd1 vccd1 _15919_/A sky130_fd_sc_hd__mux2_1
X_16898_ _16914_/A _16898_/B _16898_/C vssd1 vssd1 vccd1 vccd1 _19611_/D sky130_fd_sc_hd__nor3_1
X_19686_ _19693_/CLK _19686_/D vssd1 vssd1 vccd1 vccd1 _19686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15849_ _15849_/A vssd1 vssd1 vccd1 vccd1 _19263_/D sky130_fd_sc_hd__clkbuf_1
X_18637_ _19325_/CLK _18637_/D vssd1 vssd1 vccd1 vccd1 _18637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _18783_/Q vssd1 vssd1 vccd1 vccd1 _11001_/A sky130_fd_sc_hd__clkbuf_2
X_18568_ _19088_/CLK _18568_/D vssd1 vssd1 vccd1 vccd1 _18568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10257__C1 _09754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17519_ _17477_/X _17496_/X _17517_/Y _17518_/X _11683_/X vssd1 vssd1 vccd1 vccd1
+ _17519_/X sky130_fd_sc_hd__a32o_1
XFILLER_71_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18499_ _19091_/CLK _18499_/D vssd1 vssd1 vccd1 vccd1 _18499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12509__A _16622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11413__A _11413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10029__A _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17100__A _18071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11221__A1 _11075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12572__D_N _12571_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13774__S _13776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09553__A _09553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09706_ _10655_/A vssd1 vssd1 vccd1 vccd1 _09707_/A sky130_fd_sc_hd__buf_4
XFILLER_56_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09637_ _10579_/A vssd1 vssd1 vccd1 vccd1 _10704_/S sky130_fd_sc_hd__buf_2
XFILLER_167_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12237__B1 _19414_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09568_ _09557_/A _09567_/X _10296_/A vssd1 vssd1 vccd1 vccd1 _09568_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_169_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09653__A1 _09507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ _10633_/S vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__buf_2
XFILLER_169_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11530_ _11530_/A _11589_/A vssd1 vssd1 vccd1 vccd1 _11531_/A sky130_fd_sc_hd__nor2_1
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11461_ _11461_/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11461_/Y sky130_fd_sc_hd__nand2_1
XFILLER_139_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13200_ _19573_/Q _13006_/X _13199_/X _13012_/X vssd1 vssd1 vccd1 vccd1 _13200_/X
+ sky130_fd_sc_hd__a211o_1
X_10412_ _18929_/Q _18695_/Q _19377_/Q _19025_/Q _09681_/A _10312_/A vssd1 vssd1 vccd1
+ vccd1 _10412_/X sky130_fd_sc_hd__mux4_1
XFILLER_139_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17010__A _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09728__A _09728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14180_ _18601_/Q _14026_/X _14180_/S vssd1 vssd1 vccd1 vccd1 _14181_/A sky130_fd_sc_hd__mux2_1
X_11392_ _18943_/Q _18709_/Q _19391_/Q _19039_/Q _11388_/S _11389_/A vssd1 vssd1 vccd1
+ vccd1 _11393_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13131_ _13247_/S vssd1 vssd1 vccd1 vccd1 _13360_/S sky130_fd_sc_hd__clkbuf_2
X_10343_ _10342_/A _10340_/Y _10342_/Y _10378_/A vssd1 vssd1 vccd1 vccd1 _10343_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_125_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input55_A io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10274_ _10274_/A vssd1 vssd1 vccd1 vccd1 _10274_/X sky130_fd_sc_hd__clkbuf_4
X_13062_ _19720_/Q _15534_/B _13381_/S vssd1 vssd1 vccd1 vccd1 _13062_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13684__S _13686_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15465__A _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _19342_/Q _11859_/X _15488_/A vssd1 vssd1 vccd1 vccd1 _12013_/Y sky130_fd_sc_hd__o21ai_1
X_17870_ _17597_/A _17555_/X _17869_/X _17422_/A vssd1 vssd1 vccd1 vccd1 _17870_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16821_ _19580_/Q hold22/A _16821_/C vssd1 vssd1 vccd1 vccd1 _16824_/B sky130_fd_sc_hd__and3_1
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_181_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19305_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19540_ _19540_/CLK _19540_/D vssd1 vssd1 vccd1 vccd1 _19540_/Q sky130_fd_sc_hd__dfxtp_1
X_16752_ _19559_/Q _16752_/B _19557_/Q _16752_/D vssd1 vssd1 vccd1 vccd1 _16753_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_47_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13964_ _13964_/A vssd1 vssd1 vccd1 vccd1 _18517_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09567__S1 _10261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15703_ _15703_/A vssd1 vssd1 vccd1 vccd1 _19198_/D sky130_fd_sc_hd__clkbuf_1
X_12915_ _19144_/Q _12895_/X _12677_/X _19334_/Q _12914_/X vssd1 vssd1 vccd1 vccd1
+ _12915_/X sky130_fd_sc_hd__a221o_1
X_16683_ _19536_/Q _16687_/D _16682_/Y vssd1 vssd1 vccd1 vccd1 _19536_/D sky130_fd_sc_hd__o21a_1
X_19471_ _19471_/CLK _19471_/D vssd1 vssd1 vccd1 vccd1 _19471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_94_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13895_ _13895_/A vssd1 vssd1 vccd1 vccd1 _18497_/D sky130_fd_sc_hd__clkbuf_1
X_15634_ _15634_/A vssd1 vssd1 vccd1 vccd1 _19168_/D sky130_fd_sc_hd__clkbuf_1
X_18422_ _19239_/CLK _18422_/D vssd1 vssd1 vccd1 vccd1 _18422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12846_ _12861_/A vssd1 vssd1 vccd1 vccd1 _12848_/A sky130_fd_sc_hd__buf_2
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18353_ _19298_/CLK _18353_/D vssd1 vssd1 vccd1 vccd1 _18353_/Q sky130_fd_sc_hd__dfxtp_1
X_15565_ _15565_/A vssd1 vssd1 vccd1 vccd1 _15565_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ hold4/A _12773_/X _12422_/Y _12747_/A vssd1 vssd1 vccd1 vccd1 _18282_/D sky130_fd_sc_hd__a22o_1
XFILLER_159_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17304_ _17740_/A _17301_/X _17717_/S vssd1 vssd1 vccd1 vccd1 _17304_/X sky130_fd_sc_hd__mux2_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14516_/A vssd1 vssd1 vccd1 vccd1 _18741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11728_ _11728_/A _17252_/A vssd1 vssd1 vccd1 vccd1 _11729_/B sky130_fd_sc_hd__or2_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18284_ _19203_/CLK _18284_/D vssd1 vssd1 vccd1 vccd1 _18284_/Q sky130_fd_sc_hd__dfxtp_1
X_15496_ _19713_/Q _15495_/X _15516_/S vssd1 vssd1 vccd1 vccd1 _15496_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17235_ _17241_/A vssd1 vssd1 vccd1 vccd1 _17367_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__13859__S _13871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14447_ _14515_/S vssd1 vssd1 vccd1 vccd1 _14456_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_31_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11659_ _11698_/B vssd1 vssd1 vccd1 vccd1 _13430_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__16235__S _16235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11203__A1 _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17166_ _17166_/A _17166_/B _17166_/C _17166_/D vssd1 vssd1 vccd1 vccd1 _17185_/A
+ sky130_fd_sc_hd__or4_4
X_14378_ _13845_/X _18679_/Q _14384_/S vssd1 vssd1 vccd1 vccd1 _14379_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10411__C1 _09753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16117_ _16126_/C _16116_/Y _16109_/X vssd1 vssd1 vccd1 vccd1 _16117_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13329_ _15089_/A vssd1 vssd1 vccd1 vccd1 _14611_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17097_ _17097_/A vssd1 vssd1 vccd1 vccd1 _19694_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09357__B _17133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_134_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19799_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16048_ _15522_/X _16047_/Y _16052_/S vssd1 vssd1 vccd1 vccd1 _16048_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17890__A1 _17886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19807_ _19807_/CLK _19807_/D vssd1 vssd1 vccd1 vccd1 _19807_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09373__A _11307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_149_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19298_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_111_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17999_ _19772_/Q _19393_/Q _18005_/S vssd1 vssd1 vccd1 vccd1 _18000_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19738_ _19740_/CLK _19738_/D vssd1 vssd1 vccd1 vccd1 _19738_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__09558__S1 _10261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10312__A _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_145_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__C1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19669_ _19669_/CLK _19669_/D vssd1 vssd1 vccd1 vccd1 _19669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09422_ _11248_/A vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__buf_2
XFILLER_80_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16637__C _16659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11117__S1 _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _09339_/X _09352_/A _11647_/B _17127_/A _11652_/A vssd1 vssd1 vccd1 vccd1
+ _17112_/A sky130_fd_sc_hd__o221a_2
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _18142_/A _12696_/A _09283_/Y _19831_/Q vssd1 vssd1 vccd1 vccd1 _09284_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10796__A3 _10794_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10628__S0 _10055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15984__S _15992_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17330__B1 _09309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11053__S0 _10940_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12140__C _17779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10961_ _10961_/A _10961_/B vssd1 vssd1 vccd1 vccd1 _10961_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12700_ _12962_/A vssd1 vssd1 vccd1 vccd1 _12700_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15224__S _15228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13680_ _13294_/X _18411_/Q _13686_/S vssd1 vssd1 vccd1 vccd1 _13681_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10892_ _11138_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _10892_/X sky130_fd_sc_hd__or2_1
XFILLER_43_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12631_ _18163_/A vssd1 vssd1 vccd1 vccd1 _16341_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16844__A _18079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15350_ _19086_/Q _15044_/X _15350_/S vssd1 vssd1 vccd1 vccd1 _15351_/A sky130_fd_sc_hd__mux2_1
X_12562_ _13261_/A vssd1 vssd1 vccd1 vccd1 _12562_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14301_ _14369_/S vssd1 vssd1 vccd1 vccd1 _14310_/S sky130_fd_sc_hd__clkbuf_4
X_11513_ _11513_/A _11525_/A _11513_/C _17114_/C vssd1 vssd1 vccd1 vccd1 _17183_/B
+ sky130_fd_sc_hd__and4_1
X_15281_ _14569_/X _19055_/Q _15289_/S vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__mux2_1
X_12493_ _13389_/B _16939_/A vssd1 vssd1 vccd1 vccd1 _17028_/C sky130_fd_sc_hd__nor2_1
XANTENNA__10892__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17020_ _17020_/A _17024_/B vssd1 vssd1 vccd1 vccd1 _17020_/X sky130_fd_sc_hd__or2_1
XANTENNA__13186__A1 _15572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14232_ _14232_/A vssd1 vssd1 vccd1 vccd1 _18623_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09458__A _09981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19284_/CLK sky130_fd_sc_hd__clkbuf_16
X_11444_ _11448_/A _11451_/A _11448_/C _10495_/A vssd1 vssd1 vccd1 vccd1 _11444_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15894__S _15898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ _18593_/Q _14001_/X _14169_/S vssd1 vssd1 vccd1 vccd1 _14164_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16124__A1 _19351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11375_ _18512_/Q _19007_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _11375_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13114_ _13114_/A vssd1 vssd1 vccd1 vccd1 _13306_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10326_ _10406_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10326_/X sky130_fd_sc_hd__or2_1
XFILLER_153_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14094_ _13899_/X _18563_/Q _14096_/S vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__mux2_1
XFILLER_112_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17872__B2 _12317_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18971_ _19387_/CLK _18971_/D vssd1 vssd1 vccd1 vccd1 _18971_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output161_A _16302_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_66_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19491_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _17304_/X _17597_/X _17921_/X vssd1 vssd1 vccd1 vccd1 _17922_/X sky130_fd_sc_hd__a21o_1
X_13045_ input4/X _12974_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _13045_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10257_ _10249_/X _10252_/X _10254_/X _10256_/X _09754_/A vssd1 vssd1 vccd1 vccd1
+ _10257_/X sky130_fd_sc_hd__a221o_4
XFILLER_105_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12161__A2 _12468_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10188_ _10090_/X _10185_/X _10187_/X vssd1 vssd1 vccd1 vccd1 _10188_/X sky130_fd_sc_hd__a21o_1
X_17853_ _17856_/A _17856_/B _17896_/S vssd1 vssd1 vccd1 vccd1 _17853_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15635__B1 _13430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16804_ _19575_/Q _16802_/B _16764_/X vssd1 vssd1 vccd1 vccd1 _16804_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14996_ _14996_/A vssd1 vssd1 vccd1 vccd1 _14996_/X sky130_fd_sc_hd__clkbuf_2
X_17784_ _12123_/A _17737_/X _17783_/X _17761_/X vssd1 vssd1 vccd1 vccd1 _17784_/X
+ sky130_fd_sc_hd__o211a_4
XANTENNA__09314__B1 _11702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19523_ _19529_/CLK _19523_/D vssd1 vssd1 vccd1 vccd1 _19523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16735_ _16736_/B _16736_/C _19555_/Q vssd1 vssd1 vccd1 vccd1 _16737_/B sky130_fd_sc_hd__a21oi_1
X_13947_ _14715_/C _13947_/B _14372_/A vssd1 vssd1 vccd1 vccd1 _15854_/B sky130_fd_sc_hd__or3_4
XFILLER_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11121__B1 _09576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19454_ _19550_/CLK _19454_/D vssd1 vssd1 vccd1 vccd1 _19454_/Q sky130_fd_sc_hd__dfxtp_1
X_16666_ _16666_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16666_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11672__A1 _18114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ _13877_/X _18492_/Q _13887_/S vssd1 vssd1 vccd1 vccd1 _13879_/A sky130_fd_sc_hd__mux2_1
X_18405_ _18569_/CLK _18405_/D vssd1 vssd1 vccd1 vccd1 _18405_/Q sky130_fd_sc_hd__dfxtp_1
X_15617_ _15616_/X _19165_/Q _15627_/S vssd1 vssd1 vccd1 vccd1 _15618_/A sky130_fd_sc_hd__mux2_1
X_12829_ _12828_/X _18284_/Q _12887_/S vssd1 vssd1 vccd1 vccd1 _12830_/A sky130_fd_sc_hd__mux2_1
X_16597_ _16660_/A _16597_/B _16598_/B vssd1 vssd1 vccd1 vccd1 _19512_/D sky130_fd_sc_hd__nor3_1
XFILLER_62_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19385_ _19385_/CLK _19385_/D vssd1 vssd1 vccd1 vccd1 _19385_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16754__A _19553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15548_ _15607_/A hold10/A vssd1 vssd1 vccd1 vccd1 _15548_/Y sky130_fd_sc_hd__nand2_1
X_18336_ _19249_/CLK _18336_/D vssd1 vssd1 vccd1 vccd1 _18336_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18267_ _19725_/CLK _18267_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
X_15479_ _18255_/Q _15479_/B vssd1 vssd1 vccd1 vccd1 _15479_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_19_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19035_/CLK sky130_fd_sc_hd__clkbuf_16
X_17218_ _17218_/A vssd1 vssd1 vccd1 vccd1 _17709_/B sky130_fd_sc_hd__buf_2
XFILLER_162_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18198_ input38/X _18197_/X _18188_/X _18193_/X _12482_/A vssd1 vssd1 vccd1 vccd1
+ _18199_/B sky130_fd_sc_hd__a32o_1
XFILLER_144_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_71_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17149_ _17149_/A vssd1 vssd1 vccd1 vccd1 _17149_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11410__B _12482_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10307__A _10323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17863__A1 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ _09964_/Y _09966_/Y _09968_/Y _09970_/Y _09831_/A vssd1 vssd1 vccd1 vccd1
+ _09971_/X sky130_fd_sc_hd__o221a_2
XFILLER_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13618__A _19811_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15309__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__C1 _09658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15626__A0 _19736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11138__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10042__A _10042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09831__A _09831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17918__A2 _17232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12860__A0 _11168_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10010__S1 _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09405_ _09596_/A vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__buf_2
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15979__S _15981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09336_ _19865_/Q vssd1 vssd1 vccd1 vccd1 _18144_/A sky130_fd_sc_hd__buf_4
XFILLER_166_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13499__S _13503_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _12494_/A _09267_/B _18118_/A _09270_/B vssd1 vssd1 vccd1 vccd1 _13391_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_166_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13168__A1 input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _09194_/X _13944_/A _09196_/Y _09197_/X _19701_/Q vssd1 vssd1 vccd1 vccd1
+ _09198_/X sky130_fd_sc_hd__o221a_1
XFILLER_147_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12915__A1 _19144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12915__B2 _19334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11160_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _11160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_122_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12128__C1 _11686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10111_ _09667_/X _10101_/X _10110_/X _09758_/X _19730_/Q vssd1 vssd1 vccd1 vccd1
+ _11357_/A sky130_fd_sc_hd__a32o_4
X_11091_ _11026_/A _11090_/X _11042_/X vssd1 vssd1 vccd1 vccd1 _11091_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_136_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12432__A _12432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17606__A1 _17910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ _10042_/A _10042_/B vssd1 vssd1 vccd1 vccd1 _10042_/X sky130_fd_sc_hd__or2_1
XFILLER_102_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12151__B _19411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11048__A _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14850_ _18875_/Q _14036_/X _14854_/S vssd1 vssd1 vccd1 vccd1 _14851_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13801_ _13107_/X _18464_/Q _13809_/S vssd1 vssd1 vccd1 vccd1 _13802_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input18_A io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14781_ _14614_/X _18845_/Q _14781_/S vssd1 vssd1 vccd1 vccd1 _14782_/A sky130_fd_sc_hd__mux2_1
X_11993_ _16974_/A _11994_/C _19644_/Q vssd1 vssd1 vccd1 vccd1 _11993_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10887__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16520_ _19488_/Q _16520_/B _16915_/B vssd1 vssd1 vccd1 vccd1 _16521_/C sky130_fd_sc_hd__and3_1
X_13732_ _13138_/X _18434_/Q _13736_/S vssd1 vssd1 vccd1 vccd1 _13733_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10944_ _10937_/X _10941_/X _10942_/X _10951_/A _10943_/X vssd1 vssd1 vccd1 vccd1
+ _10949_/B sky130_fd_sc_hd__o221a_1
XANTENNA__16042__A0 _15515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16451_ _16450_/B _16450_/C _19467_/Q vssd1 vssd1 vccd1 vccd1 _16452_/C sky130_fd_sc_hd__a21oi_1
X_13663_ _13663_/A vssd1 vssd1 vccd1 vccd1 _18403_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14793__S _14799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ _11208_/A vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__buf_2
XFILLER_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15402_ _15459_/S vssd1 vssd1 vccd1 vccd1 _15411_/S sky130_fd_sc_hd__buf_2
XPHY_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12614_ _12714_/A _12614_/B vssd1 vssd1 vccd1 vccd1 _12614_/Y sky130_fd_sc_hd__nor2_1
X_19170_ _19203_/CLK _19170_/D vssd1 vssd1 vccd1 vccd1 _19170_/Q sky130_fd_sc_hd__dfxtp_1
X_16382_ _16390_/A _16387_/C vssd1 vssd1 vccd1 vccd1 _16382_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13594_ _13594_/A vssd1 vssd1 vccd1 vccd1 _18377_/D sky130_fd_sc_hd__clkbuf_1
X_18121_ _18121_/A vssd1 vssd1 vccd1 vccd1 _18135_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__17137__A3 _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15333_ _19078_/Q _15019_/X _15339_/S vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__mux2_1
X_12545_ _13400_/A vssd1 vssd1 vccd1 vccd1 _15613_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18052_ _18188_/A vssd1 vssd1 vccd1 vccd1 _18061_/S sky130_fd_sc_hd__clkbuf_2
X_15264_ _15264_/A vssd1 vssd1 vccd1 vccd1 _19047_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12476_ _12480_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _12476_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17003_ _19654_/Q _17011_/B vssd1 vssd1 vccd1 vccd1 _17003_/X sky130_fd_sc_hd__or2_1
XANTENNA__18098__A1 _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ _14215_/A vssd1 vssd1 vccd1 vccd1 _18615_/D sky130_fd_sc_hd__clkbuf_1
X_11427_ _11427_/A _11427_/B _11427_/C vssd1 vssd1 vccd1 vccd1 _11428_/B sky130_fd_sc_hd__nand3_1
X_15195_ _19017_/Q _15028_/X _15195_/S vssd1 vssd1 vccd1 vccd1 _15196_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10068__S1 _09507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14146_ _14146_/A vssd1 vssd1 vccd1 vccd1 _18585_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output86_A _12252_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11358_ _11433_/B vssd1 vssd1 vccd1 vccd1 _11358_/Y sky130_fd_sc_hd__inv_2
XFILLER_98_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10309_ _10361_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _10309_/X sky130_fd_sc_hd__or2_1
XANTENNA__13438__A _13494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14077_ _13873_/X _18555_/Q _14085_/S vssd1 vssd1 vccd1 vccd1 _14078_/A sky130_fd_sc_hd__mux2_1
X_18954_ _19006_/CLK _18954_/D vssd1 vssd1 vccd1 vccd1 _18954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11289_ _10895_/X _12450_/B _11016_/X _12448_/B _10987_/Y vssd1 vssd1 vccd1 vccd1
+ _11467_/B sky130_fd_sc_hd__o221ai_1
X_13028_ _13028_/A vssd1 vssd1 vccd1 vccd1 _18293_/D sky130_fd_sc_hd__clkbuf_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17905_ _19736_/Q _17831_/X _17904_/X vssd1 vssd1 vccd1 vccd1 _19736_/D sky130_fd_sc_hd__o21a_1
XFILLER_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18885_ _19365_/CLK _18885_/D vssd1 vssd1 vccd1 vccd1 _18885_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16749__A _19557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17836_ _17586_/X _17833_/Y _17835_/Y vssd1 vssd1 vccd1 vccd1 _17836_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09651__A _09651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17767_ _17406_/X _17764_/X _17766_/X _17537_/X vssd1 vssd1 vccd1 vccd1 _17767_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14979_ _14979_/A vssd1 vssd1 vccd1 vccd1 _18935_/D sky130_fd_sc_hd__clkbuf_1
X_19506_ _19540_/CLK _19506_/D vssd1 vssd1 vccd1 vccd1 _19506_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16718_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16718_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17698_ _17413_/A _17695_/X _17697_/Y _17494_/X vssd1 vssd1 vccd1 vccd1 _17698_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19437_ _19524_/CLK _19437_/D vssd1 vssd1 vccd1 vccd1 _19437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16649_ _19527_/Q _19526_/Q vssd1 vssd1 vccd1 vccd1 _16656_/C sky130_fd_sc_hd__and2_1
XFILLER_37_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19368_ _19369_/CLK _19368_/D vssd1 vssd1 vccd1 vccd1 _19368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09121_ _19847_/Q vssd1 vssd1 vccd1 vccd1 _09166_/A sky130_fd_sc_hd__inv_2
X_18319_ _19667_/CLK _18319_/D vssd1 vssd1 vccd1 vccd1 _18319_/Q sky130_fd_sc_hd__dfxtp_1
X_19299_ _19299_/CLK _19299_/D vssd1 vssd1 vccd1 vccd1 _19299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10620__A2 _10610_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15828__A _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10908__B1 _09561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15039__S _15045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13348__A _15092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _09954_/A vssd1 vssd1 vccd1 vccd1 _09956_/A sky130_fd_sc_hd__buf_2
XFILLER_103_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09885_ _10521_/A vssd1 vssd1 vccd1 vccd1 _09886_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_98_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11333__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14878__S _14882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16659__A _16659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09561__A _09561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16024__A0 _15495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16394__A _16549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13811__A _13822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10660_ _10660_/A vssd1 vssd1 vccd1 vccd1 _10660_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09319_ _14275_/A _15474_/A vssd1 vssd1 vccd1 vccd1 _18071_/S sky130_fd_sc_hd__or2_4
XANTENNA__11969__C _11969_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10591_ _19280_/Q _19118_/Q _18527_/Q _18297_/Q _10022_/X _10567_/X vssd1 vssd1 vccd1
+ vccd1 _10591_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14118__S _14118_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09462__C1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12427__A _17907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11331__A _11331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12330_ _12301_/X _12477_/B _12329_/Y vssd1 vssd1 vccd1 vccd1 _17878_/A sky130_fd_sc_hd__o21ai_4
XFILLER_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13957__S _13963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12261_ _12301_/A _12473_/B _12260_/Y vssd1 vssd1 vccd1 vccd1 _17845_/A sky130_fd_sc_hd__o21ai_4
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18114__A _18114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14000_ _14000_/A vssd1 vssd1 vccd1 vccd1 _18528_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13561__A1 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11212_ _11252_/A _11209_/X _11211_/X _11134_/X vssd1 vssd1 vccd1 vccd1 _11212_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_134_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12192_ _12423_/S vssd1 vssd1 vccd1 vccd1 _12404_/S sky130_fd_sc_hd__buf_2
XANTENNA__10375__A1 _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10381__S _10381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _11248_/A _11143_/B vssd1 vssd1 vccd1 vccd1 _11143_/X sky130_fd_sc_hd__or2_1
XFILLER_150_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10470__S1 _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput75 _11988_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_122_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput86 _12252_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[23] sky130_fd_sc_hd__buf_2
XFILLER_89_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput97 _11732_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[4] sky130_fd_sc_hd__buf_2
XFILLER_150_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15951_ _13547_/X _19308_/Q _15959_/S vssd1 vssd1 vccd1 vccd1 _15952_/A sky130_fd_sc_hd__mux2_1
X_11074_ _18485_/Q _18980_/Q _11074_/S vssd1 vssd1 vccd1 vccd1 _11074_/X sky130_fd_sc_hd__mux2_1
XFILLER_103_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09612__S0 _09599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14902_ _18898_/Q _14007_/X _14904_/S vssd1 vssd1 vccd1 vccd1 _14903_/A sky130_fd_sc_hd__mux2_1
X_10025_ _09557_/A _10021_/X _10024_/X vssd1 vssd1 vccd1 vccd1 _10025_/Y sky130_fd_sc_hd__o21ai_1
X_18670_ _18902_/CLK _18670_/D vssd1 vssd1 vccd1 vccd1 _18670_/Q sky130_fd_sc_hd__dfxtp_1
X_15882_ _15882_/A vssd1 vssd1 vccd1 vccd1 _19277_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16288__B _16288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17621_ _19714_/Q _17570_/X _17620_/X vssd1 vssd1 vccd1 vccd1 _19714_/D sky130_fd_sc_hd__o21a_1
XFILLER_76_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ _14833_/A vssd1 vssd1 vccd1 vccd1 _18867_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12824__A0 _09315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ _14589_/X _18837_/Q _14770_/S vssd1 vssd1 vccd1 vccd1 _14765_/A sky130_fd_sc_hd__mux2_1
X_17552_ _17576_/S _17552_/B vssd1 vssd1 vccd1 vccd1 _17552_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11976_ _17105_/A _12021_/A _12022_/A vssd1 vssd1 vccd1 vccd1 _11976_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16503_ _16541_/A _16503_/B _16503_/C vssd1 vssd1 vccd1 vccd1 _19485_/D sky130_fd_sc_hd__nor3_1
X_13715_ _13715_/A vssd1 vssd1 vccd1 vccd1 _18426_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17483_ _17483_/A vssd1 vssd1 vccd1 vccd1 _17483_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_17_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10927_ _19273_/Q _19111_/Q _18520_/Q _18290_/Q _10852_/S _10837_/A vssd1 vssd1 vccd1
+ vccd1 _10927_/X sky130_fd_sc_hd__mux4_1
XFILLER_45_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14695_ _14695_/A vssd1 vssd1 vccd1 vccd1 _18806_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17763__B1 _17762_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19222_ _19287_/CLK _19222_/D vssd1 vssd1 vccd1 vccd1 _19222_/Q sky130_fd_sc_hd__dfxtp_1
X_16434_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16470_/A sky130_fd_sc_hd__buf_2
X_13646_ _13646_/A vssd1 vssd1 vccd1 vccd1 _18395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10858_ _11111_/A vssd1 vssd1 vccd1 vccd1 _10977_/A sky130_fd_sc_hd__clkbuf_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16365_ _19437_/Q _16365_/B vssd1 vssd1 vccd1 vccd1 _16371_/C sky130_fd_sc_hd__and2_1
X_19153_ _19688_/CLK _19153_/D vssd1 vssd1 vccd1 vccd1 _19153_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13577_ _18372_/Q _13576_/X _13577_/S vssd1 vssd1 vccd1 vccd1 _13578_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ _10779_/A _10788_/X _09563_/A vssd1 vssd1 vccd1 vccd1 _10789_/Y sky130_fd_sc_hd__o21ai_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18104_ _18104_/A _18128_/B vssd1 vssd1 vccd1 vccd1 _18104_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10063__B1 _09640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15316_ _15316_/A vssd1 vssd1 vccd1 vccd1 _19071_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12528_ _13008_/A vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_172_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16296_ _16296_/A vssd1 vssd1 vccd1 vccd1 _19415_/D sky130_fd_sc_hd__clkbuf_1
X_19084_ _19086_/CLK _19084_/D vssd1 vssd1 vccd1 vccd1 _19084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12056__B _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15247_ _15315_/S vssd1 vssd1 vccd1 vccd1 _15256_/S sky130_fd_sc_hd__clkbuf_4
X_18035_ _18035_/A vssd1 vssd1 vccd1 vccd1 _19788_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12459_ _12459_/A _12461_/B vssd1 vssd1 vccd1 vccd1 _12459_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12355__A2 _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15178_ _19009_/Q _15003_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14129_ _14129_/A vssd1 vssd1 vccd1 vccd1 _18577_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10118__A1 _10174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18937_ _19391_/CLK _18937_/D vssd1 vssd1 vccd1 vccd1 _18937_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14698__S _14698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__B1 _09602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10213__S1 _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11866__A1 _11879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _09670_/A vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__buf_2
X_18868_ _19286_/CLK _18868_/D vssd1 vssd1 vccd1 vccd1 _18868_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09381__A _10031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17819_ _17820_/B _17819_/B vssd1 vssd1 vccd1 vccd1 _17823_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13068__B1 _13067_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18799_ _19249_/CLK _18799_/D vssd1 vssd1 vccd1 vccd1 _18799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11416__A _11416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09906__S1 _09905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15322__S _15328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17103__A _17163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_15_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19586_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09104_ _11525_/A vssd1 vssd1 vccd1 vccd1 _17120_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_164_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12594__A2 _12556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11229__S0 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10990__A _10990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17809__A1 _17810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__B1 _19392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11297__S _11297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15992__S _15992_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09937_ _10184_/A _09937_/B vssd1 vssd1 vccd1 vccd1 _09937_/X sky130_fd_sc_hd__or2_1
XFILLER_104_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10204__S1 _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ _09868_/A vssd1 vssd1 vccd1 vccd1 _09931_/S sky130_fd_sc_hd__clkbuf_4
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09799_ _10115_/A vssd1 vssd1 vccd1 vccd1 _09799_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_193_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11326__A _11331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ _11809_/A _11830_/B vssd1 vssd1 vccd1 vccd1 _11830_/X sky130_fd_sc_hd__and2b_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _11761_/A _17250_/A vssd1 vssd1 vccd1 vccd1 _11762_/B sky130_fd_sc_hd__or2_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18109__A _18109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14637__A _16301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13500_/A vssd1 vssd1 vccd1 vccd1 _18348_/D sky130_fd_sc_hd__clkbuf_1
X_10712_ _10773_/A _10712_/B vssd1 vssd1 vccd1 vccd1 _10712_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13541__A _15025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14502_/A vssd1 vssd1 vccd1 vccd1 _14489_/S sky130_fd_sc_hd__buf_4
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ _11686_/X _11688_/X _11689_/X _11691_/X vssd1 vssd1 vccd1 vccd1 _11692_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13431_ _13430_/X _18320_/Q _13431_/S vssd1 vssd1 vccd1 vccd1 _13432_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10643_ _10585_/A _10638_/X _10642_/X vssd1 vssd1 vccd1 vccd1 _10643_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09435__C1 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16150_ _19767_/Q _16150_/B vssd1 vssd1 vccd1 vccd1 _16150_/Y sky130_fd_sc_hd__nand2_1
X_13362_ _19769_/Q _13362_/B vssd1 vssd1 vccd1 vccd1 _13362_/X sky130_fd_sc_hd__or2_1
X_10574_ _09547_/X _10571_/Y _10573_/Y _09644_/A vssd1 vssd1 vccd1 vccd1 _10574_/X
+ sky130_fd_sc_hd__o211a_1
X_15101_ _15101_/A _15389_/B vssd1 vssd1 vccd1 vccd1 _15158_/A sky130_fd_sc_hd__nor2_2
XFILLER_10_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ _12265_/A _17845_/B _12288_/A vssd1 vssd1 vccd1 vccd1 _12314_/B sky130_fd_sc_hd__a21oi_1
X_16081_ _16091_/C _16081_/B vssd1 vssd1 vccd1 vccd1 _16081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13293_ _15083_/A vssd1 vssd1 vccd1 vccd1 _14605_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14731__A0 _14541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15032_ _15099_/S vssd1 vssd1 vccd1 vccd1 _15045_/S sky130_fd_sc_hd__buf_2
XFILLER_154_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09466__A _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12244_ _19794_/Q _11357_/A _12357_/S vssd1 vssd1 vccd1 vccd1 _12245_/A sky130_fd_sc_hd__mux2_4
XFILLER_142_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19840_ _19866_/CLK _19840_/D vssd1 vssd1 vccd1 vccd1 _19840_/Q sky130_fd_sc_hd__dfxtp_1
X_12175_ _12175_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12175_/Y sky130_fd_sc_hd__nand2_1
XFILLER_1_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11126_ _11138_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11126_/X sky130_fd_sc_hd__or2_1
XFILLER_95_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19771_ _19775_/CLK _19771_/D vssd1 vssd1 vccd1 vccd1 _19771_/Q sky130_fd_sc_hd__dfxtp_1
X_16983_ _17010_/A vssd1 vssd1 vccd1 vccd1 _16983_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_122_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13716__A _13762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18722_ _19310_/CLK _18722_/D vssd1 vssd1 vccd1 vccd1 _18722_/Q sky130_fd_sc_hd__dfxtp_1
X_15934_ _15934_/A vssd1 vssd1 vccd1 vccd1 _19300_/D sky130_fd_sc_hd__clkbuf_1
X_11057_ _09431_/A _11048_/X _11052_/X _11056_/X _10949_/A vssd1 vssd1 vccd1 vccd1
+ _11057_/X sky130_fd_sc_hd__a311o_1
XFILLER_77_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _19292_/Q _19130_/Q _18539_/Q _18309_/Q _09776_/A _10056_/A vssd1 vssd1 vccd1
+ vccd1 _10009_/B sky130_fd_sc_hd__mux4_1
X_18653_ _19271_/CLK _18653_/D vssd1 vssd1 vccd1 vccd1 _18653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15865_ _19270_/Q _14534_/A _15865_/S vssd1 vssd1 vccd1 vccd1 _15866_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17604_ _17812_/A vssd1 vssd1 vccd1 vccd1 _17910_/A sky130_fd_sc_hd__buf_2
XANTENNA__11236__A _19708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14816_ _14816_/A vssd1 vssd1 vccd1 vccd1 _18859_/D sky130_fd_sc_hd__clkbuf_1
X_18584_ _19365_/CLK _18584_/D vssd1 vssd1 vccd1 vccd1 _18584_/Q sky130_fd_sc_hd__dfxtp_1
X_15796_ _13531_/X _19239_/Q _15804_/S vssd1 vssd1 vccd1 vccd1 _15797_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17535_ _17765_/A _17535_/B vssd1 vssd1 vccd1 vccd1 _17535_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16539__A1 _16540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14747_ _14747_/A vssd1 vssd1 vccd1 vccd1 _18829_/D sky130_fd_sc_hd__clkbuf_1
X_11959_ _11959_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11960_/A sky130_fd_sc_hd__xnor2_1
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14678_ _14700_/A vssd1 vssd1 vccd1 vccd1 _14687_/S sky130_fd_sc_hd__buf_6
X_17466_ _17626_/A vssd1 vssd1 vccd1 vccd1 _17466_/X sky130_fd_sc_hd__buf_2
X_19205_ _19205_/CLK _19205_/D vssd1 vssd1 vccd1 vccd1 _19205_/Q sky130_fd_sc_hd__dfxtp_1
X_16417_ _19455_/Q _16415_/B _16402_/X vssd1 vssd1 vccd1 vccd1 _16417_/Y sky130_fd_sc_hd__a21oi_1
X_13629_ _12865_/X _18388_/Q _13631_/S vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16762__A _16762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17397_ _17512_/S _17236_/X _17396_/X vssd1 vssd1 vccd1 vccd1 _17397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_160_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19136_ _19786_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _19136_/Q sky130_fd_sc_hd__dfxtp_1
X_16348_ _16890_/A vssd1 vssd1 vccd1 vccd1 _16549_/A sky130_fd_sc_hd__buf_4
XFILLER_118_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13597__S _13609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ _18172_/A vssd1 vssd1 vccd1 vccd1 _18136_/A sky130_fd_sc_hd__buf_2
X_19067_ _19197_/CLK _19067_/D vssd1 vssd1 vccd1 vccd1 _19067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09376__A _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18018_ _18029_/A vssd1 vssd1 vccd1 vccd1 _18027_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_161_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09722_ _10200_/A vssd1 vssd1 vccd1 vccd1 _10184_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12530__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10198__S0 _09931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16002__A _16146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11303__A3 _18829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09653_ _09507_/A _09646_/Y _09651_/Y _10575_/A vssd1 vssd1 vccd1 vccd1 _09653_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09584_ _09705_/A vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__buf_2
XFILLER_83_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12264__A1 _10087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10985__A _19713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14891__S _14893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10290_ _10535_/A vssd1 vssd1 vccd1 vccd1 _10394_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12424__B _17232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17008__A _18097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13980_ _13980_/A vssd1 vssd1 vccd1 vccd1 _18522_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10189__S0 _09854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _19463_/Q vssd1 vssd1 vccd1 vccd1 _16440_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__A1 _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _15650_/A vssd1 vssd1 vccd1 vccd1 _19174_/D sky130_fd_sc_hd__clkbuf_1
X_12862_ _12891_/C _12858_/Y _12860_/X _12861_/X vssd1 vssd1 vccd1 vccd1 _12862_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_74_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11813_ _11813_/A vssd1 vssd1 vccd1 vccd1 _11890_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_14601_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14601_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15607_/A _18272_/Q vssd1 vssd1 vccd1 vccd1 _15581_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12255__A1 _19351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _18743_/Q vssd1 vssd1 vccd1 vccd1 _13065_/A sky130_fd_sc_hd__inv_2
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14532_ _14531_/X _18750_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14533_/A sky130_fd_sc_hd__mux2_1
X_17320_ _17462_/A _17316_/X _17317_/Y _17659_/A vssd1 vssd1 vccd1 vccd1 _17321_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _19630_/Q _19663_/Q vssd1 vssd1 vccd1 vccd1 _11745_/D sky130_fd_sc_hd__nand2_1
XFILLER_144_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14463_ _13864_/X _18717_/Q _14467_/S vssd1 vssd1 vccd1 vccd1 _14464_/A sky130_fd_sc_hd__mux2_1
X_17251_ _17563_/B _12309_/A _17251_/S vssd1 vssd1 vccd1 vccd1 _17251_/X sky130_fd_sc_hd__mux2_1
X_11675_ _11890_/B _12445_/B _11674_/X vssd1 vssd1 vccd1 vccd1 _17480_/A sky130_fd_sc_hd__o21a_1
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13414_ _13414_/A vssd1 vssd1 vccd1 vccd1 _18317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16202_ _13560_/X _19374_/Q _16202_/S vssd1 vssd1 vccd1 vccd1 _16203_/A sky130_fd_sc_hd__mux2_1
X_10626_ _18461_/Q _19052_/Q _19214_/Q _18429_/Q _10022_/X _10567_/X vssd1 vssd1 vccd1
+ vccd1 _10627_/B sky130_fd_sc_hd__mux4_1
X_17182_ _11566_/A _17105_/A _17122_/C _11510_/B vssd1 vssd1 vccd1 vccd1 _17183_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_168_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14394_ _14394_/A vssd1 vssd1 vccd1 vccd1 _18686_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16133_ _19764_/Q _16133_/B vssd1 vssd1 vccd1 vccd1 _16133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _19736_/Q _13344_/X _13345_/S vssd1 vssd1 vccd1 vccd1 _13345_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _10612_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10557_/X sky130_fd_sc_hd__or2_1
XFILLER_143_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12615__A _13400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14306__S _14310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__S1 _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13210__S _13252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16064_ _19752_/Q _16064_/B vssd1 vssd1 vccd1 vccd1 _16065_/B sky130_fd_sc_hd__nand2_1
XFILLER_142_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13276_ _13274_/X _18308_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _13277_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10488_ _09803_/A _10487_/X _10296_/A vssd1 vssd1 vccd1 vccd1 _10488_/X sky130_fd_sc_hd__o21a_1
XANTENNA__12334__B _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15015_ _15015_/A vssd1 vssd1 vccd1 vccd1 _15015_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_142_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12227_ _19414_/Q _12228_/B vssd1 vssd1 vccd1 vccd1 _12229_/B sky130_fd_sc_hd__nor2_1
XFILLER_97_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10135__A _11357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19823_ _19828_/CLK _19823_/D vssd1 vssd1 vccd1 vccd1 _19823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09924__A _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12158_ _19411_/Q _12093_/X _12154_/X _12157_/Y vssd1 vssd1 vccd1 vccd1 _16286_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15137__S _15145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11109_ _11042_/X _11101_/X _11104_/Y _11108_/Y _09553_/A vssd1 vssd1 vccd1 vccd1
+ _11109_/X sky130_fd_sc_hd__o311a_1
X_19754_ _19756_/CLK _19754_/D vssd1 vssd1 vccd1 vccd1 _19754_/Q sky130_fd_sc_hd__dfxtp_1
X_16966_ _15515_/X _16956_/X _16965_/X _16954_/X vssd1 vssd1 vccd1 vccd1 _19640_/D
+ sky130_fd_sc_hd__o211a_1
X_12089_ _12089_/A vssd1 vssd1 vccd1 vccd1 _12089_/X sky130_fd_sc_hd__buf_2
XFILLER_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18705_ _19387_/CLK _18705_/D vssd1 vssd1 vccd1 vccd1 _18705_/Q sky130_fd_sc_hd__dfxtp_1
X_15917_ _15917_/A vssd1 vssd1 vccd1 vccd1 _19293_/D sky130_fd_sc_hd__clkbuf_1
X_19685_ _19693_/CLK _19685_/D vssd1 vssd1 vccd1 vccd1 _19685_/Q sky130_fd_sc_hd__dfxtp_1
X_16897_ _16896_/B _16896_/C _19611_/Q vssd1 vssd1 vccd1 vccd1 _16898_/C sky130_fd_sc_hd__a21oi_1
XFILLER_49_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18636_ _19035_/CLK _18636_/D vssd1 vssd1 vccd1 vccd1 _18636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15848_ _13608_/X _19263_/Q _15848_/S vssd1 vssd1 vccd1 vccd1 _15849_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18567_ _19088_/CLK _18567_/D vssd1 vssd1 vccd1 vccd1 _18567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15779_ _15779_/A vssd1 vssd1 vccd1 vccd1 _19232_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17518_ _17596_/A vssd1 vssd1 vccd1 vccd1 _17518_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18498_ _19376_/CLK _18498_/D vssd1 vssd1 vccd1 vccd1 _18498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12509__B _12536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11413__B _12480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17449_ _17287_/X _17291_/X _17509_/S vssd1 vssd1 vccd1 vccd1 _17449_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16492__A _16549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10104__S0 _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__B1 _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10029__B _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19119_ _19119_/CLK _19119_/D vssd1 vssd1 vccd1 vccd1 _19119_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_141_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10407__S1 _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10193__C1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16999__A1 _15582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10732__A1 _10031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09705_ _09705_/A vssd1 vssd1 vccd1 vccd1 _10655_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13790__S _13798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09636_ _10773_/A vssd1 vssd1 vccd1 vccd1 _11331_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_66_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10591__S0 _10022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09567_ _19295_/Q _19133_/Q _18542_/Q _18312_/Q _10518_/S _10261_/A vssd1 vssd1 vccd1
+ vccd1 _09567_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09498_ _11318_/S vssd1 vssd1 vccd1 vccd1 _10633_/S sky130_fd_sc_hd__buf_4
XFILLER_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16923__A1 _16932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11460_ _11460_/A _11460_/B vssd1 vssd1 vccd1 vccd1 _11460_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _09728_/A _10404_/X _10406_/X _10410_/X _09753_/A vssd1 vssd1 vccd1 vccd1
+ _10411_/X sky130_fd_sc_hd__a311o_4
XFILLER_109_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ _11389_/A _11386_/Y _11389_/Y _11404_/A vssd1 vssd1 vccd1 vccd1 _11391_/X
+ sky130_fd_sc_hd__o211a_1
X_13130_ _13152_/C _13130_/B vssd1 vssd1 vccd1 vccd1 _13130_/Y sky130_fd_sc_hd__nor2_1
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ _16871_/A _12950_/X _12951_/X _16458_/A _13060_/X vssd1 vssd1 vccd1 vccd1
+ _15534_/B sky130_fd_sc_hd__a221o_2
X_10273_ _10342_/A _10269_/Y _10272_/Y _10439_/A vssd1 vssd1 vccd1 vccd1 _10273_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18122__A _18122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12012_ _11858_/S _12010_/Y _12066_/C _12068_/A vssd1 vssd1 vccd1 vccd1 _12012_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input48_A io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10723__A1 _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16820_ hold22/X _16821_/C _19580_/Q vssd1 vssd1 vccd1 vccd1 _16822_/B sky130_fd_sc_hd__a21oi_1
XFILLER_120_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17651__A2 _12773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16751_ _16799_/A _16751_/B _16758_/C vssd1 vssd1 vccd1 vccd1 _19559_/D sky130_fd_sc_hd__nor3_1
XANTENNA__13673__A0 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17680__B _17680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13963_ _18517_/Q _13962_/X _13963_/S vssd1 vssd1 vccd1 vccd1 _13964_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16577__A _16714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15702_ _14611_/X _19198_/Q _15704_/S vssd1 vssd1 vccd1 vccd1 _15703_/A sky130_fd_sc_hd__mux2_1
X_12914_ _19670_/Q _12817_/X _12680_/A _19637_/Q vssd1 vssd1 vccd1 vccd1 _12914_/X
+ sky130_fd_sc_hd__a22o_1
X_19470_ _19471_/CLK _19470_/D vssd1 vssd1 vccd1 vccd1 _19470_/Q sky130_fd_sc_hd__dfxtp_1
X_16682_ _16707_/A _16689_/D vssd1 vssd1 vccd1 vccd1 _16682_/Y sky130_fd_sc_hd__nor2_1
X_13894_ _13893_/X _18497_/Q _13903_/S vssd1 vssd1 vccd1 vccd1 _13895_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18421_ _19302_/CLK _18421_/D vssd1 vssd1 vccd1 vccd1 _18421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15633_ hold17/X _19168_/Q _15636_/S vssd1 vssd1 vccd1 vccd1 _15634_/A sky130_fd_sc_hd__mux2_1
X_12845_ _13113_/C _12845_/B vssd1 vssd1 vccd1 vccd1 _12845_/X sky130_fd_sc_hd__or2_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18352_ _19071_/CLK _18352_/D vssd1 vssd1 vccd1 vccd1 _18352_/Q sky130_fd_sc_hd__dfxtp_1
X_15564_ _15564_/A vssd1 vssd1 vccd1 vccd1 _19156_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ hold7/A _12773_/X _11413_/A _12747_/A vssd1 vssd1 vccd1 vccd1 _18281_/D sky130_fd_sc_hd__a22o_1
XANTENNA__10334__S0 _10215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17303_ _17535_/B vssd1 vssd1 vccd1 vccd1 _17717_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11728_/A _17252_/A vssd1 vssd1 vccd1 vccd1 _11729_/A sky130_fd_sc_hd__nand2_1
XFILLER_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14515_ _13940_/X _18741_/Q _14515_/S vssd1 vssd1 vccd1 vccd1 _14516_/A sky130_fd_sc_hd__mux2_1
X_15495_ _15478_/X _15493_/X _15494_/Y _13403_/X hold15/X vssd1 vssd1 vccd1 vccd1
+ _15495_/X sky130_fd_sc_hd__a32o_4
X_18283_ _19202_/CLK _18283_/D vssd1 vssd1 vccd1 vccd1 _18283_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15420__S _15422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17234_ _17305_/B vssd1 vssd1 vccd1 vccd1 _17234_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17201__A _17201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11658_ _19627_/Q _19622_/Q _11657_/Y _09295_/X vssd1 vssd1 vccd1 vccd1 _11696_/B
+ sky130_fd_sc_hd__a31o_1
X_14446_ _14502_/A vssd1 vssd1 vccd1 vccd1 _14515_/S sky130_fd_sc_hd__buf_6
XFILLER_30_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ _10614_/A _10606_/X _10608_/X _09450_/A vssd1 vssd1 vccd1 vccd1 _10609_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_7_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14377_ _14377_/A vssd1 vssd1 vccd1 vccd1 _18678_/D sky130_fd_sc_hd__clkbuf_1
X_17165_ _17165_/A _17165_/B vssd1 vssd1 vccd1 vccd1 _17166_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11589_ _11589_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _17109_/A sky130_fd_sc_hd__nor2_1
XFILLER_171_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13328_ _12855_/X _13314_/X _13317_/Y _13327_/X vssd1 vssd1 vccd1 vccd1 _15089_/A
+ sky130_fd_sc_hd__a22o_2
X_16116_ _19761_/Q _16116_/B vssd1 vssd1 vccd1 vccd1 _16116_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17096_ _19694_/Q _15631_/X _17098_/S vssd1 vssd1 vccd1 vccd1 _17097_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13259_ _19613_/Q vssd1 vssd1 vccd1 vccd1 _16904_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16047_ _16055_/C _16047_/B vssd1 vssd1 vccd1 vccd1 _16047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_170_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14560__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19806_ _19845_/CLK _19806_/D vssd1 vssd1 vccd1 vccd1 _19806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17998_ _17998_/A vssd1 vssd1 vccd1 vccd1 _19771_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19737_ _19775_/CLK _19737_/D vssd1 vssd1 vccd1 vccd1 _19737_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16949_ _16935_/A _16957_/B _16915_/A vssd1 vssd1 vccd1 vccd1 _16949_/X sky130_fd_sc_hd__a21o_1
XFILLER_93_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15391__A _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19668_ _19668_/CLK _19668_/D vssd1 vssd1 vccd1 vccd1 _19668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09421_ _18781_/Q vssd1 vssd1 vccd1 vccd1 _11248_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_92_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18619_ _18974_/CLK _18619_/D vssd1 vssd1 vccd1 vccd1 _18619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19599_ _19603_/CLK _19599_/D vssd1 vssd1 vccd1 vccd1 _19599_/Q sky130_fd_sc_hd__dfxtp_1
X_09352_ _09352_/A _11684_/C vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__or2_2
XFILLER_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09283_ _18142_/A _19585_/Q _19584_/Q vssd1 vssd1 vccd1 vccd1 _09283_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_166_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09829__A _09829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10628__S1 _11321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17765__B _17768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17330__B2 _12739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11053__S1 _11005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16397__A _16442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10960_ _18918_/Q _18684_/Q _19366_/Q _19014_/Q _09625_/A _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10961_/B sky130_fd_sc_hd__mux4_1
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11130__A1 _09416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14629__B _18207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09619_ _09644_/A _09619_/B vssd1 vssd1 vccd1 vccd1 _09619_/Y sky130_fd_sc_hd__nor2_1
X_10891_ _19273_/Q _19111_/Q _18520_/Q _18290_/Q _10878_/A _10817_/A vssd1 vssd1 vccd1
+ vccd1 _10892_/B sky130_fd_sc_hd__mux4_1
X_12630_ _16890_/A vssd1 vssd1 vccd1 vccd1 _18163_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12561_ _13356_/B vssd1 vssd1 vccd1 vccd1 _13261_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14645__A _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17021__A _18097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _11512_/A _11512_/B _11918_/B vssd1 vssd1 vccd1 vccd1 _17145_/D sky130_fd_sc_hd__and3_1
X_14300_ _14356_/A vssd1 vssd1 vccd1 vccd1 _14369_/S sky130_fd_sc_hd__buf_6
XANTENNA__09739__A _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15280_ _15302_/A vssd1 vssd1 vccd1 vccd1 _15289_/S sky130_fd_sc_hd__buf_6
X_12492_ _12543_/B _16624_/A _12548_/A vssd1 vssd1 vccd1 vccd1 _16939_/A sky130_fd_sc_hd__a21oi_2
XFILLER_141_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14231_ _18623_/Q _13994_/X _14231_/S vssd1 vssd1 vccd1 vccd1 _14232_/A sky130_fd_sc_hd__mux2_1
X_11443_ _11443_/A _11446_/A _11443_/C vssd1 vssd1 vccd1 vccd1 _11443_/Y sky130_fd_sc_hd__nand3_1
XFILLER_137_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12933__A2 _13008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14162_ _14162_/A vssd1 vssd1 vccd1 vccd1 _18592_/D sky130_fd_sc_hd__clkbuf_1
X_11374_ _18640_/Q _18975_/Q _11374_/S vssd1 vssd1 vccd1 vccd1 _11374_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13695__S _13703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13113_ _13127_/B _13113_/B _13113_/C vssd1 vssd1 vccd1 vccd1 _13113_/X sky130_fd_sc_hd__and3b_1
X_10325_ _19285_/Q _19123_/Q _18532_/Q _18302_/Q _09681_/A _10312_/A vssd1 vssd1 vccd1
+ vccd1 _10326_/B sky130_fd_sc_hd__mux4_1
X_14093_ _14093_/A vssd1 vssd1 vccd1 vccd1 _18562_/D sky130_fd_sc_hd__clkbuf_1
X_18970_ _19386_/CLK _18970_/D vssd1 vssd1 vccd1 vccd1 _18970_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15883__A1 _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _12426_/B _17589_/X _17919_/X _17920_/Y _17633_/A vssd1 vssd1 vccd1 vccd1
+ _17921_/X sky130_fd_sc_hd__a41o_1
X_13044_ _13041_/X _13043_/X _13113_/C vssd1 vssd1 vccd1 vccd1 _13044_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10256_ _10323_/A _10255_/X _09857_/A vssd1 vssd1 vccd1 vccd1 _10256_/X sky130_fd_sc_hd__o21a_1
XFILLER_106_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output154_A _16288_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ _17852_/A vssd1 vssd1 vccd1 vccd1 _17852_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10187_ _09690_/A _10186_/X _09866_/A vssd1 vssd1 vccd1 vccd1 _10187_/X sky130_fd_sc_hd__a21o_1
XFILLER_120_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15635__A1 _19738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16803_ _19574_/Q _16809_/D _16802_/Y vssd1 vssd1 vccd1 vccd1 _19574_/D sky130_fd_sc_hd__o21a_1
X_17783_ _17646_/X _17707_/X _17782_/Y _17386_/X vssd1 vssd1 vccd1 vccd1 _17783_/X
+ sky130_fd_sc_hd__a211o_1
X_14995_ _14995_/A vssd1 vssd1 vccd1 vccd1 _18943_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19522_ _19529_/CLK _19522_/D vssd1 vssd1 vccd1 vccd1 _19522_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16734_ _16736_/B _16736_/C _16733_/Y vssd1 vssd1 vccd1 vccd1 _19554_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13946_ _16619_/D _16622_/B _14642_/C vssd1 vssd1 vccd1 vccd1 _14372_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11121__A1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11121__B2 _11120_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19453_ _19524_/CLK _19453_/D vssd1 vssd1 vccd1 vccd1 _19453_/Q sky130_fd_sc_hd__dfxtp_1
X_16665_ _19531_/Q _16672_/D vssd1 vssd1 vccd1 vccd1 _16668_/B sky130_fd_sc_hd__and2_1
XFILLER_34_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13877_ _14557_/A vssd1 vssd1 vccd1 vccd1 _13877_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18404_ _19027_/CLK _18404_/D vssd1 vssd1 vccd1 vccd1 _18404_/Q sky130_fd_sc_hd__dfxtp_1
X_15616_ _19734_/Q _15615_/X _15626_/S vssd1 vssd1 vccd1 vccd1 _15616_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19384_ _19384_/CLK _19384_/D vssd1 vssd1 vccd1 vccd1 _19384_/Q sky130_fd_sc_hd__dfxtp_1
X_12828_ _14525_/A vssd1 vssd1 vccd1 vccd1 _12828_/X sky130_fd_sc_hd__clkbuf_1
X_16596_ _19512_/Q _19511_/Q _16596_/C vssd1 vssd1 vccd1 vccd1 _16598_/B sky130_fd_sc_hd__and3_1
X_18335_ _19312_/CLK _18335_/D vssd1 vssd1 vccd1 vccd1 _18335_/Q sky130_fd_sc_hd__dfxtp_1
X_15547_ _15613_/A vssd1 vssd1 vccd1 vccd1 _15607_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12773_/A vssd1 vssd1 vccd1 vccd1 _12759_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15150__S _15156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18266_ _19725_/CLK _18266_/D vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11898__B _17205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15478_ _15565_/A vssd1 vssd1 vccd1 vccd1 _15478_/X sky130_fd_sc_hd__clkbuf_2
X_17217_ _17213_/X _17216_/X _17336_/A vssd1 vssd1 vccd1 vccd1 _17217_/X sky130_fd_sc_hd__mux2_1
X_14429_ _14429_/A vssd1 vssd1 vccd1 vccd1 _18702_/D sky130_fd_sc_hd__clkbuf_1
X_18197_ _18197_/A vssd1 vssd1 vccd1 vccd1 _18197_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12075__A _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_14_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17148_ _17148_/A vssd1 vssd1 vccd1 vccd1 _19701_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_116_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _10205_/A _09969_/X _09909_/X vssd1 vssd1 vccd1 vccd1 _09970_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_157_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17079_ _19686_/Q _15588_/X _17083_/S vssd1 vssd1 vccd1 vccd1 _17080_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14290__A _14290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12803__A _16619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09384__A _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13618__B _14787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10323__A _10323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16929__B _16929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12860__A1 _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ _10889_/A vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__buf_2
XFILLER_38_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ _19859_/Q vssd1 vssd1 vccd1 vccd1 _18130_/A sky130_fd_sc_hd__buf_4
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09266_ _19823_/Q vssd1 vssd1 vccd1 vccd1 _18118_/A sky130_fd_sc_hd__inv_2
XFILLER_139_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15562__A0 _19725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_180_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19271_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17776__A _17779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ _19852_/Q _19812_/Q vssd1 vssd1 vccd1 vccd1 _09197_/X sky130_fd_sc_hd__and2_1
XFILLER_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14404__S _14406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10110_ _09730_/X _10103_/X _10105_/X _10109_/X _09754_/X vssd1 vssd1 vccd1 vccd1
+ _10110_/X sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_195_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19054_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _18453_/Q _19044_/Q _19206_/Q _18421_/Q _10969_/X _11100_/A vssd1 vssd1 vccd1
+ vccd1 _11090_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12432__B _12432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13340__A2 _12784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _19197_/Q _18811_/Q _19261_/Q _18380_/Q _09441_/X _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10042_/B sky130_fd_sc_hd__mux4_1
XFILLER_103_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13800_ _13822_/A vssd1 vssd1 vccd1 vccd1 _13809_/S sky130_fd_sc_hd__buf_6
XANTENNA__13544__A _15028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15235__S _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11992_ _19341_/Q _11766_/X _12037_/A _11991_/X _16109_/A vssd1 vssd1 vccd1 vccd1
+ _11992_/X sky130_fd_sc_hd__o221a_1
X_14780_ _14780_/A vssd1 vssd1 vccd1 vccd1 _18844_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ _13731_/A vssd1 vssd1 vccd1 vccd1 _18433_/D sky130_fd_sc_hd__clkbuf_1
X_10943_ _11007_/A vssd1 vssd1 vccd1 vccd1 _10943_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11064__A _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_133_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19756_/CLK sky130_fd_sc_hd__clkbuf_16
X_16450_ _19467_/Q _16450_/B _16450_/C vssd1 vssd1 vccd1 vccd1 _16452_/B sky130_fd_sc_hd__and3_1
XFILLER_16_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13662_ _13148_/X _18403_/Q _13664_/S vssd1 vssd1 vccd1 vccd1 _13663_/A sky130_fd_sc_hd__mux2_1
X_10874_ _11211_/A vssd1 vssd1 vccd1 vccd1 _11208_/A sky130_fd_sc_hd__buf_2
XFILLER_31_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15401_ _15401_/A vssd1 vssd1 vccd1 vccd1 _19108_/D sky130_fd_sc_hd__clkbuf_1
X_12613_ _12599_/X _12610_/X _12612_/X vssd1 vssd1 vccd1 vccd1 _12614_/B sky130_fd_sc_hd__a21oi_4
XPHY_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16381_ _19443_/Q _16381_/B vssd1 vssd1 vccd1 vccd1 _16387_/C sky130_fd_sc_hd__and2_1
X_13593_ _18377_/Q _13592_/X _13593_/S vssd1 vssd1 vccd1 vccd1 _13594_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14375__A _14443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18120_ _18134_/A vssd1 vssd1 vccd1 vccd1 _18120_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12544_ _13397_/A vssd1 vssd1 vccd1 vccd1 _12544_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09469__A _09469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15332_ _15332_/A vssd1 vssd1 vccd1 vccd1 _19077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_148_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19268_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_12_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18051_ _18051_/A vssd1 vssd1 vccd1 vccd1 _19795_/D sky130_fd_sc_hd__clkbuf_1
X_15263_ _14544_/X _19047_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15264_/A sky130_fd_sc_hd__mux2_1
X_12475_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12480_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16590__A _16812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17002_ _15588_/X _16997_/X _17001_/X _16995_/X vssd1 vssd1 vccd1 vccd1 _19653_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14214_ _18615_/Q _13969_/X _14220_/S vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__mux2_1
X_11426_ _11426_/A vssd1 vssd1 vccd1 vccd1 _11427_/C sky130_fd_sc_hd__inv_2
XFILLER_172_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18098__A2 _12694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15194_ _15194_/A vssd1 vssd1 vccd1 vccd1 _19016_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_137_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_188_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14145_ _18585_/Q _13975_/X _14147_/S vssd1 vssd1 vccd1 vccd1 _14146_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11357_ _11357_/A _12472_/B vssd1 vssd1 vccd1 vccd1 _11433_/B sky130_fd_sc_hd__nand2_1
XFILLER_141_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10308_ _18404_/Q _18665_/Q _18564_/Q _18899_/Q _09682_/A _09712_/A vssd1 vssd1 vccd1
+ vccd1 _10309_/B sky130_fd_sc_hd__mux4_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14076_ _14122_/S vssd1 vssd1 vccd1 vccd1 _14085_/S sky130_fd_sc_hd__buf_2
X_18953_ _19113_/CLK _18953_/D vssd1 vssd1 vccd1 vccd1 _18953_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output79_A _12092_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11288_ _11288_/A _12449_/B vssd1 vssd1 vccd1 vccd1 _11467_/A sky130_fd_sc_hd__nor2_1
XFILLER_112_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13027_ _13025_/X _18293_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13028_/A sky130_fd_sc_hd__mux2_1
X_17904_ _12389_/Y _17786_/A _17903_/X _12744_/A vssd1 vssd1 vccd1 vccd1 _17904_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10239_ _18597_/Q _18868_/Q _19092_/Q _18836_/Q _09700_/A _10238_/X vssd1 vssd1 vccd1
+ vccd1 _10239_/X sky130_fd_sc_hd__mux4_1
X_18884_ _19108_/CLK _18884_/D vssd1 vssd1 vccd1 vccd1 _18884_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10776__S0 _10785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17835_ _17835_/A _17835_/B vssd1 vssd1 vccd1 vccd1 _17835_/Y sky130_fd_sc_hd__nor2_1
XFILLER_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10696__A3 _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15145__S _15145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16281__A1 _12066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17766_ _17765_/A _17215_/X _17462_/X _17765_/Y vssd1 vssd1 vccd1 vccd1 _17766_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14978_ _18935_/Q vssd1 vssd1 vccd1 vccd1 _14979_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10797__B _12454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19505_ _19540_/CLK _19505_/D vssd1 vssd1 vccd1 vccd1 _19505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16717_ _19548_/Q _16722_/D _16716_/Y vssd1 vssd1 vccd1 vccd1 _19548_/D sky130_fd_sc_hd__o21a_1
X_13929_ _13928_/X _18508_/Q _13935_/S vssd1 vssd1 vccd1 vccd1 _13930_/A sky130_fd_sc_hd__mux2_1
X_17697_ _17490_/X _17694_/Y _17696_/Y vssd1 vssd1 vccd1 vccd1 _17697_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16033__A1 _19335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19436_ _19436_/CLK _19436_/D vssd1 vssd1 vccd1 vccd1 _19436_/Q sky130_fd_sc_hd__dfxtp_1
X_16648_ _19526_/Q _16644_/B _19527_/Q vssd1 vssd1 vccd1 vccd1 _16651_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19367_ _19367_/CLK _19367_/D vssd1 vssd1 vccd1 vccd1 _19367_/Q sky130_fd_sc_hd__dfxtp_1
X_16579_ _16610_/A _16584_/C vssd1 vssd1 vccd1 vccd1 _16579_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14285__A _14285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09120_ _09120_/A vssd1 vssd1 vccd1 vccd1 _17174_/A sky130_fd_sc_hd__clkbuf_4
X_18318_ _19635_/CLK _18318_/D vssd1 vssd1 vccd1 vccd1 _18318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19298_ _19298_/CLK _19298_/D vssd1 vssd1 vccd1 vccd1 _19298_/Q sky130_fd_sc_hd__dfxtp_1
X_18249_ _18249_/A vssd1 vssd1 vccd1 vccd1 _19866_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10620__A3 _10619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16931__C _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_171_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09953_ _09953_/A vssd1 vssd1 vccd1 vccd1 _09953_/Y sky130_fd_sc_hd__inv_2
XFILLER_131_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11149__A _11149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09884_ _10347_/A vssd1 vssd1 vccd1 vccd1 _10521_/A sky130_fd_sc_hd__buf_2
XFILLER_98_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11333__A1 _10639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10767__S0 _10030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_11_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19315_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16675__A _16812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_65_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19619_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09318_ _13391_/C vssd1 vssd1 vccd1 vccd1 _15474_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10590_ _10590_/A _10590_/B vssd1 vssd1 vccd1 vccd1 _10590_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09249_ _19832_/Q _19831_/Q vssd1 vssd1 vccd1 vccd1 _09253_/C sky130_fd_sc_hd__nand2_1
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _18130_/A _11516_/A _12302_/A vssd1 vssd1 vccd1 vccd1 _12260_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14642__B _18091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11211_ _11211_/A _11211_/B vssd1 vssd1 vccd1 vccd1 _11211_/X sky130_fd_sc_hd__or2_1
XFILLER_108_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14134__S _14136_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _17810_/A _12191_/B vssd1 vssd1 vccd1 vccd1 _12196_/A sky130_fd_sc_hd__xnor2_1
XFILLER_162_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11142_ _19268_/Q _19106_/Q _18515_/Q _18285_/Q _11123_/A _10933_/A vssd1 vssd1 vccd1
+ vccd1 _11143_/B sky130_fd_sc_hd__mux4_1
XANTENNA__13849__A0 _13848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput76 _12009_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[14] sky130_fd_sc_hd__buf_2
XANTENNA__11059__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 _12269_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[24] sky130_fd_sc_hd__buf_2
X_15950_ _15996_/S vssd1 vssd1 vccd1 vccd1 _15959_/S sky130_fd_sc_hd__buf_2
X_11073_ _18641_/Q vssd1 vssd1 vccd1 vccd1 _11074_/S sky130_fd_sc_hd__buf_4
Xoutput98 _11765_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18130__A _18130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09612__S1 _09419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ _14901_/A vssd1 vssd1 vccd1 vccd1 _18897_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09752__A _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input30_A io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10024_ _10590_/A _10023_/X _09640_/X vssd1 vssd1 vccd1 vccd1 _10024_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15881_ _19277_/Q _14557_/A _15887_/S vssd1 vssd1 vccd1 vccd1 _15882_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11875__A2 _11854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17620_ _11824_/Y _17786_/A _17608_/X _17619_/X _12773_/A vssd1 vssd1 vccd1 vccd1
+ _17620_/X sky130_fd_sc_hd__a221o_1
X_14832_ _18867_/Q _14010_/X _14832_/S vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_18_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19390_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13077__B2 _19342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17551_ _17364_/A _17357_/X _17609_/A vssd1 vssd1 vccd1 vccd1 _17551_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14763_ _14763_/A vssd1 vssd1 vccd1 vccd1 _18836_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11627__A2 _12443_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12824__A1 _13408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11975_ _11969_/C _11963_/X _11974_/X vssd1 vssd1 vccd1 vccd1 _11975_/X sky130_fd_sc_hd__o21a_2
XANTENNA__16015__A1 _19332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__S0 _11127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16502_ _16501_/B _16501_/C _19485_/Q vssd1 vssd1 vccd1 vccd1 _16503_/C sky130_fd_sc_hd__a21oi_1
XFILLER_72_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13714_ _12999_/X _18426_/Q _13714_/S vssd1 vssd1 vccd1 vccd1 _13715_/A sky130_fd_sc_hd__mux2_1
X_17482_ _17731_/S _17481_/X _17457_/X vssd1 vssd1 vccd1 vccd1 _17700_/A sky130_fd_sc_hd__o21ai_2
X_10926_ _10981_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10926_/Y sky130_fd_sc_hd__nor2_1
X_14694_ _14592_/X _18806_/Q _14698_/S vssd1 vssd1 vccd1 vccd1 _14695_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19221_ _19379_/CLK _19221_/D vssd1 vssd1 vccd1 vccd1 _19221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16433_ _16442_/A _16433_/B _16433_/C vssd1 vssd1 vccd1 vccd1 _19461_/D sky130_fd_sc_hd__nor3_1
XFILLER_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13645_ _13025_/X _18395_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13646_/A sky130_fd_sc_hd__mux2_1
X_10857_ _11228_/A vssd1 vssd1 vccd1 vccd1 _11111_/A sky130_fd_sc_hd__buf_2
XFILLER_60_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12618__A _13422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19152_ _19688_/CLK _19152_/D vssd1 vssd1 vccd1 vccd1 _19152_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16364_ _16388_/A _16364_/B _16365_/B vssd1 vssd1 vccd1 vccd1 _19436_/D sky130_fd_sc_hd__nor3_1
XFILLER_158_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13576_ _15060_/A vssd1 vssd1 vccd1 vccd1 _13576_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17515__A1 _17716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10788_ _18921_/Q _18687_/Q _19369_/Q _19017_/Q _09519_/A _09506_/A vssd1 vssd1 vccd1
+ vccd1 _10788_/X sky130_fd_sc_hd__mux4_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18103_ _19816_/Q _18086_/X _18102_/Y _18097_/X vssd1 vssd1 vccd1 vccd1 _19816_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10063__A1 _10680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__B1 _09469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ _14620_/X _19071_/Q _15315_/S vssd1 vssd1 vccd1 vccd1 _15316_/A sky130_fd_sc_hd__mux2_1
X_12527_ _12817_/A vssd1 vssd1 vccd1 vccd1 _13008_/A sky130_fd_sc_hd__buf_2
XFILLER_145_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19083_ _19374_/CLK _19083_/D vssd1 vssd1 vccd1 vccd1 _19083_/Q sky130_fd_sc_hd__dfxtp_1
X_16295_ _16298_/A _16295_/B vssd1 vssd1 vccd1 vccd1 _16296_/A sky130_fd_sc_hd__and2_1
XANTENNA__10138__A _10138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18034_ _19788_/Q _19409_/Q _18038_/S vssd1 vssd1 vccd1 vccd1 _18035_/A sky130_fd_sc_hd__mux2_1
X_15246_ _15302_/A vssd1 vssd1 vccd1 vccd1 _15315_/S sky130_fd_sc_hd__buf_6
X_12458_ _12458_/A vssd1 vssd1 vccd1 vccd1 _12458_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_172_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10572__S _10572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _11384_/Y _09835_/X _11398_/X _11408_/X vssd1 vssd1 vccd1 vccd1 _12482_/C
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__17818__A2 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15177_ _15177_/A vssd1 vssd1 vccd1 vccd1 _19008_/D sky130_fd_sc_hd__clkbuf_1
X_12389_ _12389_/A _12389_/B vssd1 vssd1 vccd1 vccd1 _12389_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__12760__B1 _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14128_ _18577_/Q _13943_/X _14136_/S vssd1 vssd1 vccd1 vccd1 _14129_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10771__C1 _09374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18936_ _19491_/CLK _18936_/D vssd1 vssd1 vccd1 vccd1 _18936_/Q sky130_fd_sc_hd__dfxtp_1
X_14059_ _13848_/X _18547_/Q _14063_/S vssd1 vssd1 vccd1 vccd1 _14060_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11315__A1 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A _11413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18867_ _19285_/CLK _18867_/D vssd1 vssd1 vccd1 vccd1 _18867_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold19_A hold19/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17818_ _10225_/Y _12727_/X _17817_/X vssd1 vssd1 vccd1 vccd1 _19728_/D sky130_fd_sc_hd__a21oi_1
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18798_ _19054_/CLK _18798_/D vssd1 vssd1 vccd1 vccd1 _18798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17749_ _17646_/X _17739_/X _17748_/X _17386_/X vssd1 vssd1 vccd1 vccd1 _17749_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11416__B _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17754__A1 _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19419_ _19699_/CLK _19419_/D vssd1 vssd1 vccd1 vccd1 _19419_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_74_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12528__A _13008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09103_ _09176_/A vssd1 vssd1 vccd1 vccd1 _11525_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15839__A _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11229__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14740__A1 _18826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__A1 _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14889__S _14893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17690__A0 _19718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09936_ _18409_/Q _18670_/Q _18569_/Q _18904_/Q _09868_/A _09713_/A vssd1 vssd1 vccd1
+ vccd1 _09937_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11306__A1 _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09572__A _09572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09867_ _09941_/A vssd1 vssd1 vccd1 vccd1 _10105_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_136_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ _11387_/A vssd1 vssd1 vccd1 vccd1 _11385_/S sky130_fd_sc_hd__buf_2
XANTENNA__09193__A_N _14297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11165__S0 _10964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13822__A _13822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11761_/A _17250_/A vssd1 vssd1 vccd1 vccd1 _11762_/A sky130_fd_sc_hd__nand2_1
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _18395_/Q _18656_/Q _18555_/Q _18890_/Q _11318_/S _09541_/A vssd1 vssd1 vccd1
+ vccd1 _10712_/B sky130_fd_sc_hd__mux4_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11691_ _12654_/B vssd1 vssd1 vccd1 vccd1 _11691_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11342__A _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13430_ _13430_/A _13430_/B vssd1 vssd1 vccd1 vccd1 _13430_/X sky130_fd_sc_hd__or2_1
X_10642_ _10639_/X _10641_/X _10074_/A vssd1 vssd1 vccd1 vccd1 _10642_/X sky130_fd_sc_hd__o21a_1
X_13361_ _19769_/Q _13362_/B vssd1 vssd1 vccd1 vccd1 _13370_/B sky130_fd_sc_hd__nand2_1
XFILLER_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _10693_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10573_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18125__A _18125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15100_ _15100_/A vssd1 vssd1 vccd1 vccd1 _18975_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12312_ _12312_/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12312_/Y sky130_fd_sc_hd__nor2_1
X_16080_ _19755_/Q _16080_/B vssd1 vssd1 vccd1 vccd1 _16081_/B sky130_fd_sc_hd__nand2_1
X_13292_ _13051_/X _13278_/X _13282_/Y _13291_/X vssd1 vssd1 vccd1 vccd1 _15083_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_166_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15031_ _15031_/A vssd1 vssd1 vccd1 vccd1 _15031_/X sky130_fd_sc_hd__clkbuf_2
X_12243_ _17835_/A _12243_/B vssd1 vssd1 vccd1 vccd1 _12248_/A sky130_fd_sc_hd__xnor2_1
XFILLER_163_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12742__B1 _11288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12174_ _12174_/A vssd1 vssd1 vccd1 vccd1 _12175_/B sky130_fd_sc_hd__clkinv_2
XANTENNA__14799__S _14799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__C _11560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11125_ _18914_/Q _18680_/Q _19362_/Q _19010_/Q _11173_/S _11124_/X vssd1 vssd1 vccd1
+ vccd1 _11126_/B sky130_fd_sc_hd__mux4_1
X_19770_ _19799_/CLK _19770_/D vssd1 vssd1 vccd1 vccd1 _19770_/Q sky130_fd_sc_hd__dfxtp_2
X_16982_ _15550_/X _16970_/X _16980_/X _16981_/X vssd1 vssd1 vccd1 vccd1 _19646_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18721_ _19310_/CLK _18721_/D vssd1 vssd1 vccd1 vccd1 _18721_/Q sky130_fd_sc_hd__dfxtp_1
X_11056_ _11064_/A _11053_/X _11055_/X _09447_/A vssd1 vssd1 vccd1 vccd1 _11056_/X
+ sky130_fd_sc_hd__o211a_1
X_15933_ _13522_/X _19300_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15934_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09910__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10007_ _10289_/A _10006_/X _09820_/A vssd1 vssd1 vccd1 vccd1 _10007_/Y sky130_fd_sc_hd__o21ai_1
X_18652_ _19305_/CLK _18652_/D vssd1 vssd1 vccd1 vccd1 _18652_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11517__A _17175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15864_ _15864_/A vssd1 vssd1 vccd1 vccd1 _19269_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17603_ _17603_/A vssd1 vssd1 vccd1 vccd1 _17812_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14815_ _18859_/Q _13985_/X _14821_/S vssd1 vssd1 vccd1 vccd1 _14816_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18583_ _19367_/CLK _18583_/D vssd1 vssd1 vccd1 vccd1 _18583_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15795_ _15852_/S vssd1 vssd1 vccd1 vccd1 _15804_/S sky130_fd_sc_hd__buf_2
XFILLER_92_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11156__S0 _09496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17534_ _17534_/A vssd1 vssd1 vccd1 vccd1 _17765_/A sky130_fd_sc_hd__clkbuf_2
X_14746_ _14563_/X _18829_/Q _14748_/S vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12273__A2 _12269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11958_ _11903_/A _11903_/B _11931_/A _11957_/Y vssd1 vssd1 vccd1 vccd1 _11959_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_33_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10284__A1 _09765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10909_ _11020_/A vssd1 vssd1 vccd1 vccd1 _10910_/A sky130_fd_sc_hd__clkbuf_4
X_17465_ _17659_/A vssd1 vssd1 vccd1 vccd1 _17626_/A sky130_fd_sc_hd__clkbuf_2
X_14677_ _14677_/A vssd1 vssd1 vccd1 vccd1 _18798_/D sky130_fd_sc_hd__clkbuf_1
X_11889_ _19401_/Q _11793_/X _11883_/X _11888_/Y vssd1 vssd1 vccd1 vccd1 _16262_/B
+ sky130_fd_sc_hd__o22a_1
X_19204_ _19300_/CLK _19204_/D vssd1 vssd1 vccd1 vccd1 _19204_/Q sky130_fd_sc_hd__dfxtp_1
X_16416_ _19454_/Q _16414_/B _16415_/Y vssd1 vssd1 vccd1 vccd1 _19454_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13628_ _13628_/A vssd1 vssd1 vccd1 vccd1 _18387_/D sky130_fd_sc_hd__clkbuf_1
X_17396_ _17396_/A _17396_/B vssd1 vssd1 vccd1 vccd1 _17396_/X sky130_fd_sc_hd__or2_1
XFILLER_34_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19135_ _19297_/CLK _19135_/D vssd1 vssd1 vccd1 vccd1 _19135_/Q sky130_fd_sc_hd__dfxtp_1
X_16347_ _16351_/B _16351_/C _16346_/Y vssd1 vssd1 vccd1 vccd1 _19432_/D sky130_fd_sc_hd__o21a_1
X_13559_ _13559_/A vssd1 vssd1 vccd1 vccd1 _18366_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16172__A0 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19066_ _19292_/CLK _19066_/D vssd1 vssd1 vccd1 vccd1 _19066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16278_ _16278_/A vssd1 vssd1 vccd1 vccd1 _16278_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_161_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18017_ _18017_/A vssd1 vssd1 vccd1 vccd1 _19780_/D sky130_fd_sc_hd__clkbuf_1
X_15229_ _15229_/A vssd1 vssd1 vccd1 vccd1 _19032_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12733__A0 _18254_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12811__A _13275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09721_ _10419_/A vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__buf_2
XFILLER_113_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18919_ _19076_/CLK _18919_/D vssd1 vssd1 vccd1 vccd1 _18919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12530__B _13391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10198__S1 _09871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09901__A1 _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09652_ _10773_/A vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10331__A _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09583_ _10769_/A vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11147__S0 _10962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17114__A _17114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17727__A1 _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17768__B _17768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_62_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__A _15044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12724__A0 _09194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10940__S _10940_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09919_ _18474_/Q _19065_/Q _19227_/Q _18442_/Q _09918_/X _09905_/X vssd1 vssd1 vccd1
+ vccd1 _09920_/B sky130_fd_sc_hd__mux4_1
XFILLER_101_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10189__S1 _09871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _19595_/Q vssd1 vssd1 vccd1 vccd1 _16854_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _12861_/A vssd1 vssd1 vccd1 vccd1 _12861_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14600_/A vssd1 vssd1 vccd1 vccd1 _18771_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15243__S _15243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11826_/A _11793_/X _11799_/Y _11811_/X vssd1 vssd1 vccd1 vccd1 _16255_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15580_ _18272_/Q _15580_/B vssd1 vssd1 vccd1 vccd1 _15580_/X sky130_fd_sc_hd__or2_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _09309_/X _13399_/B _13143_/S vssd1 vssd1 vccd1 vccd1 _12792_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09656__B1 _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14531_ _14531_/A vssd1 vssd1 vccd1 vccd1 _14531_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _13430_/A _11804_/B _11743_/C vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__and3b_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16926__C1 _16269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11072__A _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17250_ _17250_/A vssd1 vssd1 vccd1 vccd1 _17563_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13204__A1 _15580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14462_ _14462_/A vssd1 vssd1 vccd1 vccd1 _18716_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _11755_/A _11673_/X _11942_/A vssd1 vssd1 vccd1 vccd1 _11674_/X sky130_fd_sc_hd__a21o_2
XFILLER_30_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16201_ _16201_/A vssd1 vssd1 vccd1 vccd1 _19373_/D sky130_fd_sc_hd__clkbuf_1
X_13413_ _13412_/X _18317_/Q _13424_/S vssd1 vssd1 vccd1 vccd1 _13414_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15479__A _18255_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17181_ _17286_/S vssd1 vssd1 vccd1 vccd1 _17190_/A sky130_fd_sc_hd__clkbuf_2
X_10625_ _10682_/A _10624_/X _09630_/X vssd1 vssd1 vccd1 vccd1 _10625_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_167_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14393_ _13867_/X _18686_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14394_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18143__A1 _17125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11310__S0 _10660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09477__A _09477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16132_ _19764_/Q _16133_/B vssd1 vssd1 vccd1 vccd1 _16142_/C sky130_fd_sc_hd__or2_1
X_13344_ _19617_/Q _13260_/X _13261_/X _19485_/Q _13343_/X vssd1 vssd1 vccd1 vccd1
+ _13344_/X sky130_fd_sc_hd__a221o_4
X_10556_ _19184_/Q _18798_/Q _19248_/Q _18367_/Q _09415_/A _09443_/X vssd1 vssd1 vccd1
+ vccd1 _10557_/B sky130_fd_sc_hd__mux4_2
XFILLER_127_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12615__B _18254_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17694__A _17696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16063_ _19752_/Q _16064_/B vssd1 vssd1 vccd1 vccd1 _16073_/C sky130_fd_sc_hd__or2_1
X_10487_ _18593_/Q _18864_/Q _19088_/Q _18832_/Q _10520_/S _10347_/A vssd1 vssd1 vccd1
+ vccd1 _10487_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13275_ _13275_/A vssd1 vssd1 vccd1 vccd1 _13350_/S sky130_fd_sc_hd__buf_4
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15014_ _15014_/A vssd1 vssd1 vccd1 vccd1 _18948_/D sky130_fd_sc_hd__clkbuf_1
X_12226_ _19412_/Q _19413_/Q _12226_/C vssd1 vssd1 vccd1 vccd1 _12228_/B sky130_fd_sc_hd__and3_1
XFILLER_170_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10135__B _12472_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15418__S _15422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19822_ _19845_/CLK _19822_/D vssd1 vssd1 vccd1 vccd1 _19822_/Q sky130_fd_sc_hd__dfxtp_1
X_12157_ _11884_/X _12155_/Y _12205_/C _11835_/X vssd1 vssd1 vccd1 vccd1 _12157_/Y
+ sky130_fd_sc_hd__o31ai_1
XANTENNA__13727__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12631__A _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11108_ _11111_/A _11105_/X _11107_/X vssd1 vssd1 vccd1 vccd1 _11108_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16965_ _19640_/Q _16971_/B vssd1 vssd1 vccd1 vccd1 _16965_/X sky130_fd_sc_hd__or2_1
XFILLER_111_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12088_ _12088_/A _12120_/A vssd1 vssd1 vccd1 vccd1 _12091_/A sky130_fd_sc_hd__nor2_1
X_19753_ _19756_/CLK _19753_/D vssd1 vssd1 vccd1 vccd1 _19753_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11039_ _11219_/S vssd1 vssd1 vccd1 vccd1 _11265_/S sky130_fd_sc_hd__clkbuf_4
X_18704_ _19386_/CLK _18704_/D vssd1 vssd1 vccd1 vccd1 _18704_/Q sky130_fd_sc_hd__dfxtp_1
X_15916_ _19293_/Q _14608_/A _15920_/S vssd1 vssd1 vccd1 vccd1 _15917_/A sky130_fd_sc_hd__mux2_1
X_19684_ _19687_/CLK _19684_/D vssd1 vssd1 vccd1 vccd1 _19684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16896_ _19611_/Q _16896_/B _16896_/C vssd1 vssd1 vccd1 vccd1 _16898_/B sky130_fd_sc_hd__and3_1
X_18635_ _19386_/CLK _18635_/D vssd1 vssd1 vccd1 vccd1 _18635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15847_ _15847_/A vssd1 vssd1 vccd1 vccd1 _19262_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18566_ _19286_/CLK _18566_/D vssd1 vssd1 vccd1 vccd1 _18566_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ _13611_/X _19232_/Q _15780_/S vssd1 vssd1 vccd1 vccd1 _15779_/A sky130_fd_sc_hd__mux2_1
X_17517_ _17733_/A _17517_/B vssd1 vssd1 vccd1 vccd1 _17517_/Y sky130_fd_sc_hd__nand2_1
X_14729_ _14537_/X _18821_/Q _14737_/S vssd1 vssd1 vccd1 vccd1 _14730_/A sky130_fd_sc_hd__mux2_1
X_18497_ _19120_/CLK _18497_/D vssd1 vssd1 vccd1 vccd1 _18497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16773__A _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17448_ _17273_/X _17284_/X _17448_/S vssd1 vssd1 vccd1 vccd1 _17448_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17379_ _17379_/A vssd1 vssd1 vccd1 vccd1 _17379_/Y sky130_fd_sc_hd__inv_2
XFILLER_118_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12806__A _19811_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__S1 _10090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__S0 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19118_ _19280_/CLK _19118_/D vssd1 vssd1 vccd1 vccd1 _19118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09387__A _11297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19049_ _19243_/CLK _19049_/D vssd1 vssd1 vccd1 vccd1 _19049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11804__A_N _11743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15328__S _15328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13356__B _13356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09704_ _09743_/A vssd1 vssd1 vccd1 vccd1 _09704_/X sky130_fd_sc_hd__buf_2
XFILLER_114_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09850__A _09850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15959__A0 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ _10848_/A vssd1 vssd1 vccd1 vccd1 _10773_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10591__S1 _10567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09566_ _09803_/A _09566_/B vssd1 vssd1 vccd1 vccd1 _09566_/Y sky130_fd_sc_hd__nor2_1
XFILLER_130_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11604__B _11840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17779__A _17779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09497_ _10854_/S vssd1 vssd1 vccd1 vccd1 _11318_/S sky130_fd_sc_hd__buf_2
XANTENNA__11996__A1 _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _10404_/A _10407_/X _10409_/X _10243_/X vssd1 vssd1 vccd1 vccd1 _10410_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09297__A _19626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11390_ _11390_/A vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _18628_/Q _18963_/Q _10341_/S vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__mux2_1
XFILLER_164_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17884__B1 _17883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13060_ _19533_/Q _13004_/X _13054_/X _19501_/Q _13059_/X vssd1 vssd1 vccd1 vccd1
+ _13060_/X sky130_fd_sc_hd__a221o_2
XFILLER_151_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10272_ _10272_/A _10272_/B vssd1 vssd1 vccd1 vccd1 _10272_/Y sky130_fd_sc_hd__nand2_1
XFILLER_117_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11822__B_N _17247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ _12011_/A _19406_/Q _12011_/C vssd1 vssd1 vccd1 vccd1 _12066_/C sky130_fd_sc_hd__and3_1
XFILLER_133_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13547__A _15031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10670__S _10670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11920__A1 _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11381__C1 _09740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__B _17222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16750_ _19551_/Q _16750_/B _16750_/C _16750_/D vssd1 vssd1 vccd1 vccd1 _16758_/C
+ sky130_fd_sc_hd__and4_1
X_13962_ _14534_/A vssd1 vssd1 vccd1 vccd1 _13962_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_101_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15701_ _15701_/A vssd1 vssd1 vccd1 vccd1 _19197_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09760__A _09760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12913_ _19558_/Q vssd1 vssd1 vccd1 vccd1 _16752_/B sky130_fd_sc_hd__buf_2
X_16681_ _19536_/Q _19535_/Q _16681_/C _16681_/D vssd1 vssd1 vccd1 vccd1 _16689_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_111_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13893_ _14573_/A vssd1 vssd1 vccd1 vccd1 _13893_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18420_ _19205_/CLK _18420_/D vssd1 vssd1 vccd1 vccd1 _18420_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15632_ _19737_/Q _15631_/X _15632_/S vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__mux2_1
XFILLER_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _19709_/Q _13415_/B _13247_/S vssd1 vssd1 vccd1 vccd1 _12845_/B sky130_fd_sc_hd__mux2_1
XFILLER_62_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18351_ _19328_/CLK _18351_/D vssd1 vssd1 vccd1 vccd1 _18351_/Q sky130_fd_sc_hd__dfxtp_1
X_15563_ hold20/X _19156_/Q _15570_/S vssd1 vssd1 vccd1 vccd1 _15564_/A sky130_fd_sc_hd__mux2_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ _18280_/Q _12773_/X _11418_/A _12769_/X vssd1 vssd1 vccd1 vccd1 _18280_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16593__A _16890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17302_ _17391_/A vssd1 vssd1 vccd1 vccd1 _17535_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15178__A1 _15003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14514_/A vssd1 vssd1 vccd1 vccd1 _18740_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _19775_/Q _11070_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _17252_/A sky130_fd_sc_hd__mux2_4
X_18282_ _18282_/CLK _18282_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_2
X_15494_ _15494_/A hold15/A vssd1 vssd1 vccd1 vccd1 _15494_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17233_ _12487_/B _17251_/S _17232_/X vssd1 vssd1 vccd1 vccd1 _17305_/B sky130_fd_sc_hd__o21ai_4
XFILLER_70_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14445_ _15926_/B _15245_/B vssd1 vssd1 vccd1 vccd1 _14502_/A sky130_fd_sc_hd__nand2_4
X_11657_ _19628_/Q _19623_/Q vssd1 vssd1 vccd1 vccd1 _11657_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12626__A _18099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11739__A1 _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10098__S0 _10137_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10608_ _10617_/A _10608_/B vssd1 vssd1 vccd1 vccd1 _10608_/X sky130_fd_sc_hd__or2_1
X_17164_ _17164_/A vssd1 vssd1 vccd1 vccd1 _19706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14376_ _13837_/X _18678_/Q _14384_/S vssd1 vssd1 vccd1 vccd1 _14377_/A sky130_fd_sc_hd__mux2_1
X_11588_ _11525_/A _09158_/A _09211_/A _09176_/B _09169_/B vssd1 vssd1 vccd1 vccd1
+ _11591_/C sky130_fd_sc_hd__a41o_1
XANTENNA__10411__A1 _09728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16115_ _19761_/Q _16116_/B vssd1 vssd1 vccd1 vccd1 _16126_/C sky130_fd_sc_hd__or2_1
XANTENNA__17875__A0 _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13327_ _12861_/X _13326_/X _12976_/A vssd1 vssd1 vccd1 vccd1 _13327_/X sky130_fd_sc_hd__o21a_1
X_17095_ _17095_/A vssd1 vssd1 vccd1 vccd1 _19693_/D sky130_fd_sc_hd__clkbuf_1
X_10539_ _19722_/Q vssd1 vssd1 vccd1 vccd1 _10539_/Y sky130_fd_sc_hd__inv_2
XFILLER_142_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16046_ _19749_/Q _16046_/B vssd1 vssd1 vccd1 vccd1 _16047_/B sky130_fd_sc_hd__nand2_1
X_13258_ _13281_/B _13257_/Y _11499_/X vssd1 vssd1 vccd1 vccd1 _13258_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_142_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15148__S _15156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12209_ _12209_/A vssd1 vssd1 vccd1 vccd1 _12302_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13189_ _13177_/X _13187_/Y _13188_/Y vssd1 vssd1 vccd1 vccd1 _15063_/A sky130_fd_sc_hd__a21oi_4
X_19805_ _19845_/CLK _19805_/D vssd1 vssd1 vccd1 vccd1 _19805_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17997_ _19771_/Q _19392_/Q _18005_/S vssd1 vssd1 vccd1 vccd1 _17998_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16768__A _16778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13891__S _13903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16948_ _13418_/B _16943_/X _16947_/Y _16933_/X vssd1 vssd1 vccd1 vccd1 _19633_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19736_ _19736_/CLK _19736_/D vssd1 vssd1 vccd1 vccd1 _19736_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09670__A _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09963__S0 _10168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11675__B1 _11674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19667_ _19667_/CLK _19667_/D vssd1 vssd1 vccd1 vccd1 _19667_/Q sky130_fd_sc_hd__dfxtp_1
X_16879_ _19605_/Q _16879_/B _16879_/C vssd1 vssd1 vccd1 vccd1 _16881_/B sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_10_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14288__A _14288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13192__A _13275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09420_ _18941_/Q _18707_/Q _19389_/Q _19037_/Q _10496_/A _09671_/A vssd1 vssd1 vccd1
+ vccd1 _09420_/X sky130_fd_sc_hd__mux4_1
XFILLER_93_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18618_ _19081_/CLK _18618_/D vssd1 vssd1 vccd1 vccd1 _18618_/Q sky130_fd_sc_hd__dfxtp_1
X_19598_ _19598_/CLK _19598_/D vssd1 vssd1 vccd1 vccd1 _19598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _09351_/A _17126_/C _09350_/X vssd1 vssd1 vccd1 vccd1 _11684_/C sky130_fd_sc_hd__or3b_1
X_18549_ _19301_/CLK _18549_/D vssd1 vssd1 vccd1 vccd1 _18549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10325__S1 _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09282_ _19585_/Q vssd1 vssd1 vccd1 vccd1 _12696_/A sky130_fd_sc_hd__buf_2
XFILLER_166_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18207__B _18207_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12536__A _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14227__S _14231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10056__A _10056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15566__B _15566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12271__A _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09580__A _19736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10469__B2 _19723_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09618_ _19200_/Q _18814_/Q _19264_/Q _18383_/Q _09538_/A _09547_/A vssd1 vssd1 vccd1
+ vccd1 _09619_/B sky130_fd_sc_hd__mux4_1
X_10890_ _18456_/Q _19047_/Q _19209_/Q _18424_/Q _11049_/S _10817_/X vssd1 vssd1 vccd1
+ vccd1 _10890_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09549_ _10014_/A _09548_/X _09485_/A vssd1 vssd1 vccd1 vccd1 _09549_/X sky130_fd_sc_hd__o21a_1
XFILLER_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12560_ _13260_/A vssd1 vssd1 vccd1 vccd1 _12560_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _11511_/A _11511_/B vssd1 vssd1 vccd1 vccd1 _11512_/A sky130_fd_sc_hd__nor2_1
XFILLER_169_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ _12619_/A _16931_/A vssd1 vssd1 vccd1 vccd1 _13389_/B sky130_fd_sc_hd__or2_1
XFILLER_12_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13041__S _13143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14230_ _14230_/A vssd1 vssd1 vccd1 vccd1 _18622_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11442_ _11446_/A _11443_/C _11443_/A vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14161_ _18592_/Q _13997_/X _14169_/S vssd1 vssd1 vccd1 vccd1 _14162_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11373_ _11373_/A _11373_/B vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__or2_1
XFILLER_166_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10324_ _18468_/Q _19059_/Q _19221_/Q _18436_/Q _10367_/S _10314_/A vssd1 vssd1 vccd1
+ vccd1 _10324_/X sky130_fd_sc_hd__mux4_1
XANTENNA_input60_A io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13112_ _16069_/A _13095_/A _13083_/B _19755_/Q vssd1 vssd1 vccd1 vccd1 _13113_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_153_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14092_ _13896_/X _18562_/Q _14096_/S vssd1 vssd1 vccd1 vccd1 _14093_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10255_ _18469_/Q _19060_/Q _19222_/Q _18437_/Q _10247_/X _09712_/A vssd1 vssd1 vccd1
+ vccd1 _10255_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ _17920_/A _17920_/B vssd1 vssd1 vccd1 vccd1 _17920_/Y sky130_fd_sc_hd__nand2_1
X_13043_ _16055_/B _13064_/C vssd1 vssd1 vccd1 vccd1 _13043_/X sky130_fd_sc_hd__xor2_1
XFILLER_140_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17851_ _09972_/Y _12727_/X _17850_/X vssd1 vssd1 vccd1 vccd1 _19731_/D sky130_fd_sc_hd__a21oi_1
X_10186_ _18502_/Q _18997_/Q _10186_/S vssd1 vssd1 vccd1 vccd1 _10186_/X sky130_fd_sc_hd__mux2_1
X_16802_ _16840_/A _16802_/B vssd1 vssd1 vccd1 vccd1 _16802_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15635__A2 _16024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17782_ _17597_/X _17717_/X _17781_/X vssd1 vssd1 vccd1 vccd1 _17782_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_66_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14994_ _18943_/Q vssd1 vssd1 vccd1 vccd1 _14995_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_75_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18034__A0 _19788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16733_ _16736_/B _16736_/C _16718_/X vssd1 vssd1 vccd1 vccd1 _16733_/Y sky130_fd_sc_hd__a21oi_1
X_19521_ _19529_/CLK _19521_/D vssd1 vssd1 vccd1 vccd1 _19521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13945_ _18089_/A _14787_/B vssd1 vssd1 vccd1 vccd1 _15317_/A sky130_fd_sc_hd__or2_1
XFILLER_35_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19452_ _19550_/CLK _19452_/D vssd1 vssd1 vccd1 vccd1 _19452_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_184_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16664_ _16696_/A _16664_/B _16672_/D vssd1 vssd1 vccd1 vccd1 _19530_/D sky130_fd_sc_hd__nor3_1
X_13876_ _13876_/A vssd1 vssd1 vccd1 vccd1 _18491_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18403_ _19284_/CLK _18403_/D vssd1 vssd1 vccd1 vccd1 _18403_/Q sky130_fd_sc_hd__dfxtp_1
X_15615_ _15612_/X _18278_/Q _09234_/X _13398_/X _15614_/X vssd1 vssd1 vccd1 vccd1
+ _15615_/X sky130_fd_sc_hd__a32o_4
X_19383_ _19383_/CLK _19383_/D vssd1 vssd1 vccd1 vccd1 _19383_/Q sky130_fd_sc_hd__dfxtp_1
X_12827_ _15003_/A vssd1 vssd1 vccd1 vccd1 _14525_/A sky130_fd_sc_hd__clkbuf_2
X_16595_ _19511_/Q _16596_/C _19512_/Q vssd1 vssd1 vccd1 vccd1 _16597_/B sky130_fd_sc_hd__a21oi_1
XFILLER_90_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15431__S _15433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16754__C _16754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18334_ _19309_/CLK _18334_/D vssd1 vssd1 vccd1 vccd1 _18334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15546_ hold10/A _15546_/B vssd1 vssd1 vccd1 vccd1 _15546_/X sky130_fd_sc_hd__or2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12758_ _18268_/Q _12752_/X _11445_/A _12755_/X vssd1 vssd1 vccd1 vccd1 _18268_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11709_ _19634_/Q _11778_/B vssd1 vssd1 vccd1 vccd1 _11709_/X sky130_fd_sc_hd__and2_1
XFILLER_148_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18265_ _19201_/CLK _18265_/D vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_2
X_15477_ _15477_/A vssd1 vssd1 vccd1 vccd1 _19141_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12689_ _12544_/X _12687_/X _12688_/Y _12549_/X _18274_/Q vssd1 vssd1 vccd1 vccd1
+ _12689_/X sky130_fd_sc_hd__a32o_4
XANTENNA__12356__A _17886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17216_ _17722_/B _17215_/X _17261_/S vssd1 vssd1 vccd1 vccd1 _17216_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14428_ _13918_/X _18702_/Q _14428_/S vssd1 vssd1 vccd1 vccd1 _14429_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18196_ _18196_/A vssd1 vssd1 vccd1 vccd1 _19847_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17147_ _17160_/A _17147_/B vssd1 vssd1 vccd1 vccd1 _17148_/A sky130_fd_sc_hd__and2_1
X_14359_ _13925_/X _18672_/Q _14365_/S vssd1 vssd1 vccd1 vccd1 _14360_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10396__B1 _10297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09665__A _09665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17078_ _17078_/A vssd1 vssd1 vccd1 vccd1 _19685_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14290__B _18222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12137__A1 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16029_ _16039_/C _16029_/B vssd1 vssd1 vccd1 vccd1 _16029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_112_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10699__A1 _10074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16284__C1 _16280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18025__A0 _19784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19719_ _19736_/CLK _19719_/D vssd1 vssd1 vccd1 vccd1 _19719_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09403_ _11254_/A vssd1 vssd1 vccd1 vccd1 _10889_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ _19864_/Q _19863_/Q vssd1 vssd1 vccd1 vccd1 _11584_/B sky130_fd_sc_hd__or2_1
XFILLER_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17122__A _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12612__A2 _12586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09265_ _16625_/A _12508_/C _12606_/A vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__nor3_4
XFILLER_138_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15562__A1 _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09196_ _19852_/Q _19812_/Q vssd1 vssd1 vccd1 vccd1 _09196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_147_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17776__B _17779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13796__S _13798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15577__A _15603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16172__S _16180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09294__B _12621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10040_ _10040_/A _10040_/B _10040_/C vssd1 vssd1 vccd1 vccd1 _10040_/X sky130_fd_sc_hd__or3_4
XFILLER_114_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_49_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkbuf_2
XFILLER_76_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14420__S _14428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11991_ _11990_/X _11988_/Y _12100_/A vssd1 vssd1 vccd1 vccd1 _11991_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12300__A1 _19417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17731__S _17731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13730_ _13124_/X _18433_/Q _13736_/S vssd1 vssd1 vccd1 vccd1 _13731_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10942_ _18918_/Q _18684_/Q _19366_/Q _19014_/Q _11172_/S _11174_/A vssd1 vssd1 vccd1
+ vccd1 _10942_/X sky130_fd_sc_hd__mux4_1
XFILLER_72_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13661_ _13661_/A vssd1 vssd1 vccd1 vccd1 _18402_/D sky130_fd_sc_hd__clkbuf_1
X_10873_ _18488_/Q _18983_/Q _10873_/S vssd1 vssd1 vccd1 vccd1 _10873_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14656__A _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15400_ _19108_/Q _15012_/X _15400_/S vssd1 vssd1 vccd1 vccd1 _15401_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13560__A _15044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12612_ _19491_/Q _12586_/B _13261_/A _19459_/Q _12611_/X vssd1 vssd1 vccd1 vccd1
+ _12612_/X sky130_fd_sc_hd__a221o_2
X_16380_ _16388_/A _16380_/B _16381_/B vssd1 vssd1 vccd1 vccd1 _19442_/D sky130_fd_sc_hd__nor3_1
XPHY_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13592_ _15076_/A vssd1 vssd1 vccd1 vccd1 _13592_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15331_ _19077_/Q _15015_/X _15339_/S vssd1 vssd1 vccd1 vccd1 _15332_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12543_ _19700_/Q _12543_/B vssd1 vssd1 vccd1 vccd1 _13397_/A sky130_fd_sc_hd__and2b_2
XFILLER_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12176__A _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11080__A _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18050_ _19795_/Q _19416_/Q _18050_/S vssd1 vssd1 vccd1 vccd1 _18051_/A sky130_fd_sc_hd__mux2_1
X_15262_ _15262_/A vssd1 vssd1 vccd1 vccd1 _19046_/D sky130_fd_sc_hd__clkbuf_1
X_12474_ _12474_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _12474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17001_ _19653_/Q _17011_/B vssd1 vssd1 vccd1 vccd1 _17001_/X sky130_fd_sc_hd__or2_1
X_14213_ _14213_/A vssd1 vssd1 vccd1 vccd1 _18614_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11425_ _11433_/A _11431_/C _11423_/Y _11424_/Y vssd1 vssd1 vccd1 vccd1 _11428_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_126_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15193_ _19016_/Q _15025_/X _15195_/S vssd1 vssd1 vccd1 vccd1 _15194_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ _14144_/A vssd1 vssd1 vccd1 vccd1 _18584_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09485__A _09485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ _11439_/A _11441_/A _11439_/C _10304_/A _11355_/Y vssd1 vssd1 vccd1 vccd1
+ _11435_/C sky130_fd_sc_hd__a311o_1
XFILLER_153_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10307_ _10323_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10307_/X sky130_fd_sc_hd__or2_1
XFILLER_98_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14075_ _14075_/A vssd1 vssd1 vccd1 vccd1 _18554_/D sky130_fd_sc_hd__clkbuf_1
X_18952_ _19113_/CLK _18952_/D vssd1 vssd1 vccd1 vccd1 _18952_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11287_ _11464_/A _11285_/X _11465_/B vssd1 vssd1 vccd1 vccd1 _11287_/X sky130_fd_sc_hd__a21o_1
XFILLER_112_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13026_ _13387_/S vssd1 vssd1 vccd1 vccd1 _13091_/S sky130_fd_sc_hd__buf_2
X_17903_ _17852_/X _17459_/Y _17902_/X _17860_/X vssd1 vssd1 vccd1 vccd1 _17903_/X
+ sky130_fd_sc_hd__o211a_1
X_10238_ _10238_/A vssd1 vssd1 vccd1 vccd1 _10238_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_117_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11239__B _12443_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__B1 _19401_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18883_ _19108_/CLK _18883_/D vssd1 vssd1 vccd1 vccd1 _18883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10776__S1 _09506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16749__C _19553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10169_ _10169_/A _10169_/B vssd1 vssd1 vccd1 vccd1 _10169_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14330__S _14332_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17834_ _17832_/X _17833_/Y _17855_/S vssd1 vssd1 vccd1 vccd1 _17834_/X sky130_fd_sc_hd__mux2_1
XFILLER_120_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14977_ _14977_/A vssd1 vssd1 vccd1 vccd1 _18934_/D sky130_fd_sc_hd__clkbuf_1
X_17765_ _17765_/A _17768_/B vssd1 vssd1 vccd1 vccd1 _17765_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19504_ _19540_/CLK _19504_/D vssd1 vssd1 vccd1 vccd1 _19504_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15950__A _15996_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16716_ _16762_/A _16724_/D vssd1 vssd1 vccd1 vccd1 _16716_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13928_ _14608_/A vssd1 vssd1 vccd1 vccd1 _13928_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17696_ _17696_/A _17696_/B vssd1 vssd1 vccd1 vccd1 _17696_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19435_ _19524_/CLK _19435_/D vssd1 vssd1 vccd1 vccd1 _19435_/Q sky130_fd_sc_hd__dfxtp_1
X_16647_ _19526_/Q _16644_/B _16646_/Y vssd1 vssd1 vccd1 vccd1 _19526_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13859_ _13857_/X _18486_/Q _13871_/S vssd1 vssd1 vccd1 vccd1 _13860_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14566__A _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15161__S _15167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16578_ _19507_/Q _16578_/B vssd1 vssd1 vccd1 vccd1 _16584_/C sky130_fd_sc_hd__and2_1
XFILLER_37_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19366_ _19366_/CLK _19366_/D vssd1 vssd1 vccd1 vccd1 _19366_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__A1 _09390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18317_ _19667_/CLK _18317_/D vssd1 vssd1 vccd1 vccd1 _18317_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11702__B _12696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15529_ _15528_/X _19149_/Q _15544_/S vssd1 vssd1 vccd1 vccd1 _15530_/A sky130_fd_sc_hd__mux2_1
X_19297_ _19297_/CLK _19297_/D vssd1 vssd1 vccd1 vccd1 _19297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18248_ _18248_/A _18248_/B vssd1 vssd1 vccd1 vccd1 _18249_/A sky130_fd_sc_hd__and2_1
X_18179_ input64/X _18178_/X _18168_/X _18174_/X _19843_/Q vssd1 vssd1 vccd1 vccd1
+ _18180_/B sky130_fd_sc_hd__a32o_1
XFILLER_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14505__S _14511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10464__S0 _10499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09952_ _18505_/Q _19000_/Q _09952_/S vssd1 vssd1 vccd1 vccd1 _09953_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09883_ _09955_/S vssd1 vssd1 vccd1 vccd1 _10114_/S sky130_fd_sc_hd__clkbuf_4
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18220__B _18220_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10767__S1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14240__S _14242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14283__A1 input47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14283__B2 _18122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11286__A2_N _12447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15071__S _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _11551_/A _11551_/B vssd1 vssd1 vccd1 vccd1 _13391_/C sky130_fd_sc_hd__or2_1
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11612__B _17317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10509__A _10509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _19830_/Q _19829_/Q _19828_/Q _19827_/Q vssd1 vssd1 vccd1 vccd1 _16625_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_166_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_132_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14415__S _14417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _09179_/A _09208_/A vssd1 vssd1 vccd1 vccd1 _17145_/B sky130_fd_sc_hd__or2_2
XFILLER_31_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ _18450_/Q _19041_/Q _19203_/Q _18418_/Q _11065_/A _11124_/A vssd1 vssd1 vccd1
+ vccd1 _11211_/B sky130_fd_sc_hd__mux4_2
XANTENNA__10455__S0 _10499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12190_ _12305_/A _17802_/A _12164_/B vssd1 vssd1 vccd1 vccd1 _12191_/B sky130_fd_sc_hd__a21oi_1
XFILLER_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12443__B _12443_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _18451_/Q _19042_/Q _19204_/Q _18419_/Q _11050_/S _10934_/A vssd1 vssd1 vccd1
+ vccd1 _11141_/X sky130_fd_sc_hd__mux4_2
XFILLER_150_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11072_ _11072_/A _11072_/B vssd1 vssd1 vccd1 vccd1 _11072_/Y sky130_fd_sc_hd__nand2_1
Xoutput77 _12035_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[15] sky130_fd_sc_hd__buf_2
Xoutput88 _12291_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_95_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput99 _11796_/A vssd1 vssd1 vccd1 vccd1 io_dbus_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14900_ _18897_/Q _14004_/X _14904_/S vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10023_ _18603_/Q _18874_/Q _19098_/Q _18842_/Q _10022_/X _09651_/A vssd1 vssd1 vccd1
+ vccd1 _10023_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_1_clock clkbuf_1_0_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_103_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15880_ _15880_/A vssd1 vssd1 vccd1 vccd1 _19276_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14150__S _14158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14831_ _14831_/A vssd1 vssd1 vccd1 vccd1 _18866_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input23_A io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15471__B1 _13419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11075__A _11075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17550_ _17456_/X _17549_/Y _17550_/S vssd1 vssd1 vccd1 vccd1 _17657_/A sky130_fd_sc_hd__mux2_1
X_14762_ _14585_/X _18836_/Q _14770_/S vssd1 vssd1 vccd1 vccd1 _14763_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11974_ _11974_/A _12134_/A _11973_/X vssd1 vssd1 vccd1 vccd1 _11974_/X sky130_fd_sc_hd__or3b_1
XFILLER_16_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16501_ _19485_/Q _16501_/B _16501_/C vssd1 vssd1 vccd1 vccd1 _16503_/B sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_57_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13713_ _13713_/A vssd1 vssd1 vccd1 vccd1 _18425_/D sky130_fd_sc_hd__clkbuf_1
X_17481_ _17244_/X _17457_/B _17500_/S vssd1 vssd1 vccd1 vccd1 _17481_/X sky130_fd_sc_hd__mux2_1
X_10925_ _18456_/Q _19047_/Q _19209_/Q _18424_/Q _10862_/X _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10926_/B sky130_fd_sc_hd__mux4_1
X_14693_ _14693_/A vssd1 vssd1 vccd1 vccd1 _18805_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14386__A _14443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17763__A2 _17652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19220_ _19378_/CLK _19220_/D vssd1 vssd1 vccd1 vccd1 _19220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16432_ _16431_/B _16431_/C _19461_/Q vssd1 vssd1 vccd1 vccd1 _16433_/C sky130_fd_sc_hd__a21oi_1
XFILLER_108_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13644_ _13690_/S vssd1 vssd1 vccd1 vccd1 _13653_/S sky130_fd_sc_hd__buf_2
XFILLER_71_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10856_ _10968_/A vssd1 vssd1 vccd1 vccd1 _11228_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_72_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19151_ _19693_/CLK _19151_/D vssd1 vssd1 vccd1 vccd1 _19151_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _19436_/Q _19435_/Q _16363_/C vssd1 vssd1 vccd1 vccd1 _16365_/B sky130_fd_sc_hd__and3_1
XFILLER_9_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13575_/A vssd1 vssd1 vccd1 vccd1 _18371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10787_ _09651_/A _10784_/Y _10786_/Y _10575_/A vssd1 vssd1 vccd1 vccd1 _10787_/X
+ sky130_fd_sc_hd__o211a_1
X_18102_ _18102_/A _18128_/B vssd1 vssd1 vccd1 vccd1 _18102_/Y sky130_fd_sc_hd__nand2_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ _15314_/A vssd1 vssd1 vccd1 vccd1 _19070_/D sky130_fd_sc_hd__clkbuf_1
X_12526_ _13179_/A vssd1 vssd1 vccd1 vccd1 _12526_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19082_ _19085_/CLK _19082_/D vssd1 vssd1 vccd1 vccd1 _19082_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11260__A1 _09366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16294_ _16292_/Y _12134_/X _12232_/X _12236_/X _16293_/X vssd1 vssd1 vccd1 vccd1
+ _19414_/D sky130_fd_sc_hd__a221oi_1
XFILLER_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18033_ _18033_/A vssd1 vssd1 vccd1 vccd1 _19787_/D sky130_fd_sc_hd__clkbuf_1
X_15245_ _15710_/A _15245_/B vssd1 vssd1 vccd1 vccd1 _15302_/A sky130_fd_sc_hd__nand2_4
XFILLER_157_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12457_ _12462_/B _12457_/B vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__and2b_1
XANTENNA_output91_A _12369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11408_ _09831_/X _11407_/X _09762_/X vssd1 vssd1 vccd1 vccd1 _11408_/X sky130_fd_sc_hd__a21o_1
XFILLER_114_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15176_ _19008_/Q _14996_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15177_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12388_ _12388_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _12389_/B sky130_fd_sc_hd__nand2_2
XFILLER_153_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14127_ _14195_/S vssd1 vssd1 vccd1 vccd1 _14136_/S sky130_fd_sc_hd__buf_4
XFILLER_67_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _19720_/Q vssd1 vssd1 vccd1 vccd1 _11339_/Y sky130_fd_sc_hd__inv_2
XFILLER_114_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14058_ _14058_/A vssd1 vssd1 vccd1 vccd1 _18546_/D sky130_fd_sc_hd__clkbuf_1
X_18935_ _19391_/CLK _18935_/D vssd1 vssd1 vccd1 vccd1 _18935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15156__S _15156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13009_ _13009_/A vssd1 vssd1 vccd1 vccd1 _13009_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09662__B _12480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18866_ _19091_/CLK _18866_/D vssd1 vssd1 vccd1 vccd1 _18866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17817_ _12200_/A _17737_/X _17816_/X _17761_/X vssd1 vssd1 vccd1 vccd1 _17817_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18797_ _19247_/CLK _18797_/D vssd1 vssd1 vccd1 vccd1 _18797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12276__B1 _15632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17748_ _17419_/X _17741_/X _17747_/Y _17852_/A vssd1 vssd1 vccd1 vccd1 _17748_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10826__A1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17679_ _17710_/S _17676_/Y _17678_/X _17466_/X vssd1 vssd1 vccd1 vccd1 _17679_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14296__A _14296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17754__A2 _12089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19418_ _19802_/CLK _19418_/D vssd1 vssd1 vccd1 vccd1 _19418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_168_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_194_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19184_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10039__C1 _09989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12579__B2 _19346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19349_ _19349_/CLK _19349_/D vssd1 vssd1 vccd1 vccd1 _19349_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09102_ _11528_/B vssd1 vssd1 vccd1 vccd1 _09176_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15517__A1 _19147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10685__S0 _10022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__S _10763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12544__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15855__A _15911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_132_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _18282_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_171_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09935_ _18601_/Q _18872_/Q _19096_/Q _18840_/Q _10137_/S _10090_/A vssd1 vssd1 vccd1
+ vccd1 _09935_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17690__A1 _17688_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10999__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09866_ _09866_/A vssd1 vssd1 vccd1 vccd1 _09941_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_147_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19267_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09797_ _11389_/A _09784_/Y _09788_/Y _09817_/A vssd1 vssd1 vccd1 vccd1 _09797_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_93_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_81_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12019__B1 _12014_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10710_ _10705_/X _10707_/Y _10074_/A _10709_/Y vssd1 vssd1 vccd1 vccd1 _10710_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ _12184_/A vssd1 vssd1 vccd1 vccd1 _12654_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10641_ _18589_/Q _18860_/Q _19084_/Q _18828_/Q _09519_/A _10705_/A vssd1 vssd1 vccd1
+ vccd1 _10641_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11342__B _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ _19737_/Q _13359_/X _13360_/S vssd1 vssd1 vccd1 vccd1 _13360_/X sky130_fd_sc_hd__mux2_1
XFILLER_166_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10572_ _18623_/Q _18958_/Q _10572_/S vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__mux2_1
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12311_ _12311_/A vssd1 vssd1 vccd1 vccd1 _12347_/A sky130_fd_sc_hd__inv_2
XFILLER_158_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13291_ _12861_/X _13290_/X _12831_/X vssd1 vssd1 vccd1 vccd1 _13291_/X sky130_fd_sc_hd__o21a_1
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12454__A _12454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15030_ _15030_/A vssd1 vssd1 vccd1 vccd1 _18953_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10428__S0 _10381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ _17305_/A _12242_/B vssd1 vssd1 vccd1 vccd1 _12243_/B sky130_fd_sc_hd__or2_1
XFILLER_107_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10202__C1 _09754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12742__A1 hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12173_ _12173_/A _12173_/B vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__xnor2_2
XFILLER_150_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11124_ _11124_/A vssd1 vssd1 vccd1 vccd1 _11124_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__17681__A1 _17910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16981_ _16981_/A vssd1 vssd1 vccd1 vccd1 _16981_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18720_ _19370_/CLK _18720_/D vssd1 vssd1 vccd1 vccd1 _18720_/Q sky130_fd_sc_hd__dfxtp_1
X_11055_ _11195_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11055_/X sky130_fd_sc_hd__or2_1
X_15932_ _15932_/A vssd1 vssd1 vccd1 vccd1 _19299_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10006_ _19324_/Q _18736_/Q _18773_/Q _18347_/Q _09539_/A _09543_/A vssd1 vssd1 vccd1
+ vccd1 _10006_/X sky130_fd_sc_hd__mux4_1
X_15863_ _19269_/Q _14531_/A _15865_/S vssd1 vssd1 vccd1 vccd1 _15864_/A sky130_fd_sc_hd__mux2_1
X_18651_ _19271_/CLK _18651_/D vssd1 vssd1 vccd1 vccd1 _18651_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10600__S0 _10546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15704__S _15704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17602_ _17600_/X _17601_/Y _17744_/S vssd1 vssd1 vccd1 vccd1 _17602_/X sky130_fd_sc_hd__mux2_1
X_14814_ _14814_/A vssd1 vssd1 vccd1 vccd1 _18858_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15794_ _15794_/A vssd1 vssd1 vccd1 vccd1 _19238_/D sky130_fd_sc_hd__clkbuf_1
X_18582_ _19365_/CLK _18582_/D vssd1 vssd1 vccd1 vccd1 _18582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11156__S1 _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17533_ _17535_/B _17252_/X vssd1 vssd1 vccd1 vccd1 _17533_/X sky130_fd_sc_hd__or2b_1
X_14745_ _14745_/A vssd1 vssd1 vccd1 vccd1 _18828_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11957_ _11900_/A _11927_/A _11929_/B vssd1 vssd1 vccd1 vccd1 _11957_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12629__A _16245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17464_ _17907_/A _17461_/A _17462_/X _17463_/X vssd1 vssd1 vccd1 vccd1 _17464_/X
+ sky130_fd_sc_hd__o211a_1
X_10908_ _10961_/A _10907_/X _09561_/A vssd1 vssd1 vccd1 vccd1 _10908_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14676_ _14566_/X _18798_/Q _14676_/S vssd1 vssd1 vccd1 vccd1 _14677_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11481__B2 _11492_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ _11884_/X _11885_/Y _11939_/C _11962_/A vssd1 vssd1 vccd1 vccd1 _11888_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_60_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16415_ _16427_/A _16415_/B vssd1 vssd1 vccd1 vccd1 _16415_/Y sky130_fd_sc_hd__nor2_1
X_19203_ _19203_/CLK _19203_/D vssd1 vssd1 vccd1 vccd1 _19203_/Q sky130_fd_sc_hd__dfxtp_1
X_13627_ _12851_/X _18387_/Q _13631_/S vssd1 vssd1 vccd1 vccd1 _13628_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17395_ _17396_/B vssd1 vssd1 vccd1 vccd1 _17395_/Y sky130_fd_sc_hd__clkinv_2
X_10839_ _10839_/A _10839_/B vssd1 vssd1 vccd1 vccd1 _10839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16346_ _16351_/B _16351_/C _16293_/X vssd1 vssd1 vccd1 vccd1 _16346_/Y sky130_fd_sc_hd__a21oi_1
X_19134_ _19328_/CLK _19134_/D vssd1 vssd1 vccd1 vccd1 _19134_/Q sky130_fd_sc_hd__dfxtp_1
X_13558_ _18366_/Q _13557_/X _13561_/S vssd1 vssd1 vccd1 vccd1 _13559_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12509_ _16622_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _13054_/A sky130_fd_sc_hd__nor2_2
XFILLER_121_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19065_ _19291_/CLK _19065_/D vssd1 vssd1 vccd1 vccd1 _19065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16277_ _16277_/A vssd1 vssd1 vccd1 vccd1 _19407_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14055__S _14063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13489_ _13489_/A vssd1 vssd1 vccd1 vccd1 _18343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15228_ _19032_/Q _15076_/X _15228_/S vssd1 vssd1 vccd1 vccd1 _15229_/A sky130_fd_sc_hd__mux2_1
X_18016_ _19780_/Q _19401_/Q _18016_/S vssd1 vssd1 vccd1 vccd1 _18017_/A sky130_fd_sc_hd__mux2_1
XFILLER_161_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13894__S _13903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15159_ _19001_/Q _15079_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15160_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09673__A _10229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19541_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09720_ _10461_/A vssd1 vssd1 vccd1 vccd1 _10419_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_80_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18918_ _19366_/CLK _18918_/D vssd1 vssd1 vccd1 vccd1 _18918_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09651_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09651_/Y sky130_fd_sc_hd__nand2_1
XFILLER_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18849_ _19712_/CLK _18849_/D vssd1 vssd1 vccd1 vccd1 _18849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09582_ _10823_/A vssd1 vssd1 vccd1 vccd1 _10769_/A sky130_fd_sc_hd__buf_2
XFILLER_83_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11147__S1 _11075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17727__A2 _17722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10658__S0 _10650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A _10670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10432__C1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16163__A1 _19358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12274__A _19352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19325_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_128_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16180__S _16180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09583__A _10769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11618__A _11618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ _10166_/S vssd1 vssd1 vccd1 vccd1 _09918_/X sky130_fd_sc_hd__buf_2
XFILLER_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09849_ _10546_/S vssd1 vssd1 vccd1 vccd1 _09850_/A sky130_fd_sc_hd__clkbuf_4
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17305__A _17305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12860_ _11168_/Y _12614_/B _13345_/S vssd1 vssd1 vccd1 vccd1 _12860_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11773_/X _11810_/X _11623_/X vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__a21o_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09656__A1 _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12791_ _13114_/A vssd1 vssd1 vccd1 vccd1 _13143_/S sky130_fd_sc_hd__buf_2
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14530_ _14530_/A vssd1 vssd1 vccd1 vccd1 _18749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _19634_/Q _11705_/B _11706_/X vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__a21bo_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14461_ _13861_/X _18716_/Q _14467_/S vssd1 vssd1 vccd1 vccd1 _14462_/A sky130_fd_sc_hd__mux2_1
XFILLER_53_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12883__S _13144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11673_ _19845_/Q _11672_/X _11721_/S vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__mux2_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18136__A _18136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16200_ _13557_/X _19373_/Q _16202_/S vssd1 vssd1 vccd1 vccd1 _16201_/A sky130_fd_sc_hd__mux2_1
X_13412_ _11705_/B _13410_/X _15482_/S vssd1 vssd1 vccd1 vccd1 _13412_/X sky130_fd_sc_hd__mux2_1
X_17180_ _17274_/A vssd1 vssd1 vccd1 vccd1 _17286_/S sky130_fd_sc_hd__clkbuf_2
X_10624_ _19310_/Q _18722_/Q _18759_/Q _18333_/Q _10055_/S _11321_/A vssd1 vssd1 vccd1
+ vccd1 _10624_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15479__B _15479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14392_ _14392_/A vssd1 vssd1 vccd1 vccd1 _18685_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18143__A2 _18091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ _16131_/A vssd1 vssd1 vccd1 vccd1 _19352_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11310__S1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13343_ _16724_/C _12583_/X _12635_/X _19517_/Q _13342_/X vssd1 vssd1 vccd1 vccd1
+ _13343_/X sky130_fd_sc_hd__a221o_1
XFILLER_128_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ _09995_/X _10544_/X _10549_/X _10554_/X _10040_/A vssd1 vssd1 vccd1 vccd1
+ _10555_/X sky130_fd_sc_hd__a311o_4
XFILLER_154_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16062_ _16062_/A vssd1 vssd1 vccd1 vccd1 _19340_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17694__B _17696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ _14601_/A vssd1 vssd1 vccd1 vccd1 _13274_/X sky130_fd_sc_hd__clkbuf_1
X_10486_ _18401_/Q _18662_/Q _18561_/Q _18896_/Q _10274_/A _10348_/A vssd1 vssd1 vccd1
+ vccd1 _10486_/X sky130_fd_sc_hd__mux4_1
X_15013_ _18948_/Q _15012_/X _15013_/S vssd1 vssd1 vccd1 vccd1 _15014_/A sky130_fd_sc_hd__mux2_1
X_12225_ _12435_/A _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/Y sky130_fd_sc_hd__nand2_1
XFILLER_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14603__S _14615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19821_ _19845_/CLK _19821_/D vssd1 vssd1 vccd1 vccd1 _19821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12156_ _19650_/Q _19649_/Q _12156_/C vssd1 vssd1 vccd1 vccd1 _12205_/C sky130_fd_sc_hd__and3_1
XFILLER_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11107_ _09531_/A _11106_/X _11042_/A vssd1 vssd1 vccd1 vccd1 _11107_/X sky130_fd_sc_hd__o21a_1
X_19752_ _19756_/CLK _19752_/D vssd1 vssd1 vccd1 vccd1 _19752_/Q sky130_fd_sc_hd__dfxtp_1
X_16964_ _15509_/X _16956_/X _16963_/X _16954_/X vssd1 vssd1 vccd1 vccd1 _19639_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12087_ _12087_/A _17215_/A vssd1 vssd1 vccd1 vccd1 _12120_/A sky130_fd_sc_hd__nor2_1
X_18703_ _19385_/CLK _18703_/D vssd1 vssd1 vccd1 vccd1 _18703_/Q sky130_fd_sc_hd__dfxtp_1
X_11038_ _18582_/Q _18853_/Q _19077_/Q _18821_/Q _09496_/A _11100_/A vssd1 vssd1 vccd1
+ vccd1 _11038_/X sky130_fd_sc_hd__mux4_1
X_15915_ _15915_/A vssd1 vssd1 vccd1 vccd1 _19292_/D sky130_fd_sc_hd__clkbuf_1
X_19683_ _19688_/CLK _19683_/D vssd1 vssd1 vccd1 vccd1 _19683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16895_ _16896_/B _16896_/C _16894_/Y vssd1 vssd1 vccd1 vccd1 _19610_/D sky130_fd_sc_hd__o21a_1
XFILLER_37_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18634_ _19197_/CLK _18634_/D vssd1 vssd1 vccd1 vccd1 _18634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17215__A _17215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15846_ _13605_/X _19262_/Q _15848_/S vssd1 vssd1 vccd1 vccd1 _15847_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18565_ _18569_/CLK _18565_/D vssd1 vssd1 vccd1 vccd1 _18565_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12989_ _19433_/Q _13005_/A _12988_/X vssd1 vssd1 vccd1 vccd1 _12989_/X sky130_fd_sc_hd__o21a_1
X_15777_ _15777_/A vssd1 vssd1 vccd1 vccd1 _19231_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17516_ _17505_/Y _17515_/Y _17648_/S vssd1 vssd1 vccd1 vccd1 _17517_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10888__S0 _11172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14728_ _14785_/S vssd1 vssd1 vccd1 vccd1 _14737_/S sky130_fd_sc_hd__buf_2
XANTENNA__16917__B1 _16344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18496_ _19119_/CLK _18496_/D vssd1 vssd1 vccd1 vccd1 _18496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17447_ _17445_/X _17446_/X _17609_/A vssd1 vssd1 vccd1 vccd1 _17654_/B sky130_fd_sc_hd__mux2_1
X_14659_ _14541_/X _18790_/Q _14665_/S vssd1 vssd1 vccd1 vccd1 _14660_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09668__A _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17378_ _17552_/B _17377_/X _17613_/A vssd1 vssd1 vccd1 vccd1 _17379_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12806__B _14297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19117_ _19373_/CLK _19117_/D vssd1 vssd1 vccd1 vccd1 _19117_/Q sky130_fd_sc_hd__dfxtp_1
X_16329_ _16331_/B _16331_/C _16328_/Y vssd1 vssd1 vccd1 vccd1 _19426_/D sky130_fd_sc_hd__o21a_1
XFILLER_119_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17885__A _17886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12094__A _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19048_ _19243_/CLK _19048_/D vssd1 vssd1 vccd1 vccd1 _19048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_179_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12706__A1 _12696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14513__S _14515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10193__A1 _09844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10342__A _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09703_ _10094_/S vssd1 vssd1 vccd1 vccd1 _09743_/A sky130_fd_sc_hd__buf_2
XFILLER_96_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15344__S _15350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17125__A _17125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ _10682_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09565_ _18478_/Q _19069_/Q _19231_/Q _18446_/Q _10479_/S _09768_/A vssd1 vssd1 vccd1
+ vccd1 _09566_/B sky130_fd_sc_hd__mux4_1
XFILLER_43_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14631__A1 input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14631__B2 _18112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__S0 _11172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11604__C _11668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ _09496_/A vssd1 vssd1 vccd1 vccd1 _10854_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__17779__B _17779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16136__A1 _19353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11620__B _18087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17795__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ _10340_/A vssd1 vssd1 vccd1 vccd1 _10340_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17884__A1 _19734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10271_ _18629_/Q _18964_/Q _10381_/S vssd1 vssd1 vccd1 vccd1 _10272_/B sky130_fd_sc_hd__mux2_1
X_12010_ _12011_/A _12011_/C _19406_/Q vssd1 vssd1 vccd1 vccd1 _12010_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17636__A1 _11855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10803__S0 _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13039__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13961_ _13961_/A vssd1 vssd1 vccd1 vccd1 _18516_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09877__A1 _09667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09877__B2 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15254__S _15256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13563__A _15047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12912_ _16021_/B _12928_/C vssd1 vssd1 vccd1 vccd1 _12912_/X sky130_fd_sc_hd__xor2_1
XANTENNA__18061__A1 _12391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15700_ _14608_/X _19197_/Q _15704_/S vssd1 vssd1 vccd1 vccd1 _15701_/A sky130_fd_sc_hd__mux2_1
X_16680_ _16696_/A _16680_/B _16687_/D vssd1 vssd1 vccd1 vccd1 _19535_/D sky130_fd_sc_hd__nor3_1
X_13892_ _13892_/A vssd1 vssd1 vccd1 vccd1 _18496_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15631_ _15612_/X hold7/X _09234_/X _15630_/X vssd1 vssd1 vccd1 vccd1 _15631_/X sky130_fd_sc_hd__a31o_4
X_12843_ _18745_/Q vssd1 vssd1 vccd1 vccd1 _13247_/S sky130_fd_sc_hd__buf_2
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_opt_4_0_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15562_ _19725_/Q _12593_/B _15569_/S vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__mux2_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18350_ _19197_/CLK _18350_/D vssd1 vssd1 vccd1 vccd1 _18350_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _18279_/Q _12773_/X _11416_/A _12769_/X vssd1 vssd1 vccd1 vccd1 _18279_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_6_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_17301_ _17281_/X _17298_/X _17653_/A vssd1 vssd1 vccd1 vccd1 _17301_/X sky130_fd_sc_hd__mux2_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _13937_/X _18740_/Q _14515_/S vssd1 vssd1 vccd1 vccd1 _14514_/A sky130_fd_sc_hd__mux2_1
X_11725_ _11725_/A _17391_/A vssd1 vssd1 vccd1 vccd1 _11728_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10644__C1 _09658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15493_ hold15/A _15493_/B vssd1 vssd1 vccd1 vccd1 _15493_/X sky130_fd_sc_hd__or2_1
XANTENNA__17322__C_N _17319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18281_ _18282_/CLK _18281_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_2
XFILLER_30_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17232_ _17232_/A _17240_/S vssd1 vssd1 vccd1 vccd1 _17232_/X sky130_fd_sc_hd__or2b_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09488__A _11232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14444_ _14444_/A vssd1 vssd1 vccd1 vccd1 _18709_/D sky130_fd_sc_hd__clkbuf_1
X_11656_ _11644_/Y _11651_/X _11655_/Y vssd1 vssd1 vccd1 vccd1 _11656_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10607_ _18397_/Q _18658_/Q _18557_/Q _18892_/Q _10670_/S _09590_/A vssd1 vssd1 vccd1
+ vccd1 _10608_/B sky130_fd_sc_hd__mux4_1
X_17163_ _17163_/A _17163_/B vssd1 vssd1 vccd1 vccd1 _17164_/A sky130_fd_sc_hd__and2_1
XANTENNA__10098__S1 _09714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14375_ _14443_/S vssd1 vssd1 vccd1 vccd1 _14384_/S sky130_fd_sc_hd__buf_2
X_11587_ _11587_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _11591_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16114_ _16114_/A vssd1 vssd1 vccd1 vccd1 _16114_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13326_ _19735_/Q _13325_/X _13345_/S vssd1 vssd1 vccd1 vccd1 _13326_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17094_ _19693_/Q _15625_/X _17094_/S vssd1 vssd1 vccd1 vccd1 _17095_/A sky130_fd_sc_hd__mux2_1
X_10538_ _10531_/Y _10533_/Y _10535_/Y _10537_/Y _09830_/A vssd1 vssd1 vccd1 vccd1
+ _10538_/X sky130_fd_sc_hd__o221a_4
XFILLER_170_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_180_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15429__S _15433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16045_ _19749_/Q _16046_/B vssd1 vssd1 vccd1 vccd1 _16055_/C sky130_fd_sc_hd__or2_2
XANTENNA__13738__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11047__S0 _11196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13257_ _13245_/A _13256_/C _19764_/Q vssd1 vssd1 vccd1 vccd1 _13257_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_170_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10469_ _09666_/A _10459_/X _10468_/X _09757_/A _19723_/Q vssd1 vssd1 vccd1 vccd1
+ _10494_/A sky130_fd_sc_hd__a32o_4
XANTENNA__16114__A _16114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17627__A1 _17630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12208_ _12208_/A vssd1 vssd1 vccd1 vccd1 _12301_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13188_ input13/X _13166_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _13188_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_9_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19804_ _19845_/CLK _19804_/D vssd1 vssd1 vccd1 vccd1 _19804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12139_ _17790_/A vssd1 vssd1 vccd1 vccd1 _12142_/A sky130_fd_sc_hd__inv_2
XANTENNA__10162__A _10174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17996_ _18029_/A vssd1 vssd1 vccd1 vccd1 _18005_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__14310__A0 _13854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19735_ _19780_/CLK _19735_/D vssd1 vssd1 vccd1 vccd1 _19735_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_84_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16947_ _16947_/A _16970_/A vssd1 vssd1 vccd1 vccd1 _16947_/Y sky130_fd_sc_hd__nand2_1
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11675__A1 _11890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19666_ _19668_/CLK _19666_/D vssd1 vssd1 vccd1 vccd1 _19666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16878_ _16879_/B _16879_/C _16877_/Y vssd1 vssd1 vccd1 vccd1 _19604_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18617_ _19367_/CLK _18617_/D vssd1 vssd1 vccd1 vccd1 _18617_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15829_ _13579_/X _19254_/Q _15837_/S vssd1 vssd1 vccd1 vccd1 _15830_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19597_ _19598_/CLK _19597_/D vssd1 vssd1 vccd1 vccd1 _19597_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12089__A _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09350_ _17125_/A _18140_/A _18122_/A vssd1 vssd1 vccd1 vccd1 _09350_/X sky130_fd_sc_hd__and3_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18548_ _19205_/CLK _18548_/D vssd1 vssd1 vccd1 vccd1 _18548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10635__C1 _11331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09281_ _19832_/Q vssd1 vssd1 vccd1 vccd1 _18142_/A sky130_fd_sc_hd__inv_2
XFILLER_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18479_ _19264_/CLK _18479_/D vssd1 vssd1 vccd1 vccd1 _18479_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13412__S _15482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12536__B _12536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__S0 _09496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13352__A1 input24/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12271__B _19416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11902__A2 _11854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A _19710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09861__A _10197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15074__S _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10469__A2 _10459_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10013__S1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__B1 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09617_ _09617_/A vssd1 vssd1 vccd1 vccd1 _09617_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_71_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09548_ _18414_/Q _18675_/Q _18574_/Q _18909_/Q _09539_/A _09547_/X vssd1 vssd1 vccd1
+ vccd1 _09548_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09479_ _18644_/Q vssd1 vssd1 vccd1 vccd1 _10914_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12727__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15103__A _15171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11510_ _17166_/A _11510_/B vssd1 vssd1 vccd1 vccd1 _17145_/C sky130_fd_sc_hd__nor2_1
XFILLER_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12490_ _12490_/A vssd1 vssd1 vccd1 vccd1 _16931_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12918__B2 _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _11441_/A _11441_/B vssd1 vssd1 vccd1 vccd1 _11441_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14160_ _14182_/A vssd1 vssd1 vccd1 vccd1 _14169_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_164_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11372_ _18943_/Q _18709_/Q _19391_/Q _19039_/Q _11375_/S _09715_/X vssd1 vssd1 vccd1
+ vccd1 _11373_/B sky130_fd_sc_hd__mux4_1
XFILLER_165_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13111_ _19754_/Q _19755_/Q _13111_/C vssd1 vssd1 vccd1 vccd1 _13127_/B sky130_fd_sc_hd__and3_1
X_10323_ _10323_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10323_/X sky130_fd_sc_hd__or2_1
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14091_ _14091_/A vssd1 vssd1 vccd1 vccd1 _18561_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12462__A _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input53_A io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13042_ _19751_/Q vssd1 vssd1 vccd1 vccd1 _16055_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10254_ _10361_/A _10254_/B vssd1 vssd1 vccd1 vccd1 _10254_/X sky130_fd_sc_hd__or2_1
XFILLER_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13992__S _13995_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17850_ _12269_/A _17737_/A _17849_/Y _17761_/X vssd1 vssd1 vccd1 vccd1 _17850_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_78_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10185_ _18630_/Q _18965_/Q _10185_/S vssd1 vssd1 vccd1 vccd1 _10185_/X sky130_fd_sc_hd__mux2_1
XFILLER_78_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16801_ _19574_/Q _16809_/D vssd1 vssd1 vccd1 vccd1 _16802_/B sky130_fd_sc_hd__and2_1
XANTENNA__09771__A _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17781_ _17673_/A _17778_/X _17780_/X _17633_/A vssd1 vssd1 vccd1 vccd1 _17781_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_120_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14993_ _14993_/A vssd1 vssd1 vccd1 vccd1 _18942_/D sky130_fd_sc_hd__clkbuf_1
X_19520_ _19529_/CLK _19520_/D vssd1 vssd1 vccd1 vccd1 _19520_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13293__A _15083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18034__A1 _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ _16737_/A _16732_/B _16736_/C vssd1 vssd1 vccd1 vccd1 _19553_/D sky130_fd_sc_hd__nor3_1
XFILLER_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13944_ _13944_/A vssd1 vssd1 vccd1 vccd1 _18089_/A sky130_fd_sc_hd__buf_6
XFILLER_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_127_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19451_ _19524_/CLK _19451_/D vssd1 vssd1 vccd1 vccd1 _19451_/Q sky130_fd_sc_hd__dfxtp_1
X_16663_ _19530_/Q _19529_/Q _19528_/Q _16663_/D vssd1 vssd1 vccd1 vccd1 _16672_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13875_ _13873_/X _18491_/Q _13887_/S vssd1 vssd1 vccd1 vccd1 _13876_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18402_ _19377_/CLK _18402_/D vssd1 vssd1 vccd1 vccd1 _18402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15614_ _13306_/B _15613_/Y _18278_/Q vssd1 vssd1 vccd1 vccd1 _15614_/X sky130_fd_sc_hd__mux2_1
X_12826_ input12/X _12781_/X _12825_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _15003_/A
+ sky130_fd_sc_hd__a22o_1
X_19382_ _19382_/CLK _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Q sky130_fd_sc_hd__dfxtp_1
X_16594_ _16806_/A vssd1 vssd1 vccd1 vccd1 _16660_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18333_ _19248_/CLK _18333_/D vssd1 vssd1 vccd1 vccd1 _18333_/Q sky130_fd_sc_hd__dfxtp_1
X_15545_ _15545_/A vssd1 vssd1 vccd1 vccd1 _19152_/D sky130_fd_sc_hd__clkbuf_1
X_12757_ hold8/A _12752_/X _10494_/A _12755_/X vssd1 vssd1 vccd1 vccd1 _18267_/D sky130_fd_sc_hd__a22o_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14328__S _14332_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16109__A _16109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11708_ _11708_/A vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__inv_2
XFILLER_148_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15476_ _15475_/X _19141_/Q _15483_/S vssd1 vssd1 vccd1 vccd1 _15477_/A sky130_fd_sc_hd__mux2_1
X_18264_ _19201_/CLK _18264_/D vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_2
XFILLER_129_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12688_ _12713_/A _18274_/Q vssd1 vssd1 vccd1 vccd1 _12688_/Y sky130_fd_sc_hd__nand2_1
XFILLER_147_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14427_ _14427_/A vssd1 vssd1 vccd1 vccd1 _18701_/D sky130_fd_sc_hd__clkbuf_1
X_17215_ _17215_/A vssd1 vssd1 vccd1 vccd1 _17215_/X sky130_fd_sc_hd__buf_2
X_11639_ _11639_/A vssd1 vssd1 vccd1 vccd1 _11644_/B sky130_fd_sc_hd__clkinv_4
X_18195_ _18231_/A _18195_/B vssd1 vssd1 vccd1 vccd1 _18196_/A sky130_fd_sc_hd__and2_1
XFILLER_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09946__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17146_ _19701_/Q _17140_/A _17145_/Y _18099_/A vssd1 vssd1 vccd1 vccd1 _17147_/B
+ sky130_fd_sc_hd__a22o_1
X_14358_ _14358_/A vssd1 vssd1 vccd1 vccd1 _18671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10396__A1 _10378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13309_ _12798_/X _13297_/Y _13308_/X vssd1 vssd1 vccd1 vccd1 _15086_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__15159__S _15167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17077_ _19685_/Q _15582_/X _17083_/S vssd1 vssd1 vccd1 vccd1 _17078_/A sky130_fd_sc_hd__mux2_1
X_14289_ input49/X _14282_/X _14277_/X _14278_/X _18127_/A vssd1 vssd1 vccd1 vccd1
+ _18222_/B sky130_fd_sc_hd__a32o_2
XFILLER_115_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14063__S _14063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16028_ _19746_/Q _16028_/B vssd1 vssd1 vccd1 vccd1 _16029_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09633__S0 _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17979_ _13245_/A _19795_/Q _17979_/S vssd1 vssd1 vccd1 vccd1 _17980_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18025__A1 _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19718_ _19736_/CLK _19718_/D vssd1 vssd1 vccd1 vccd1 _19718_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__16036__A0 _15509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19649_ _19649_/CLK _19649_/D vssd1 vssd1 vccd1 vccd1 _19649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09402_ _11211_/A vssd1 vssd1 vccd1 vccd1 _11254_/A sky130_fd_sc_hd__buf_2
XFILLER_77_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18218__B _18218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09333_ _09351_/A vssd1 vssd1 vccd1 vccd1 _17126_/B sky130_fd_sc_hd__inv_2
XANTENNA__13270__A0 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14238__S _14242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _09270_/A vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11281__C1 _10929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09195_ _19811_/Q vssd1 vssd1 vccd1 vccd1 _13944_/A sky130_fd_sc_hd__inv_2
XANTENNA__10067__A _10684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18234__A _18234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09856__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10387__A1 _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09872__S0 _09930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12128__A2 _12123_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14701__S _14709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18016__A1 _19401_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11990_ _12011_/A _12011_/C vssd1 vssd1 vccd1 vccd1 _11990_/X sky130_fd_sc_hd__xor2_1
XFILLER_21_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10941_ _09393_/A _10940_/X _10807_/A vssd1 vssd1 vccd1 vccd1 _10941_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17775__A0 _17779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13660_ _13138_/X _18402_/Q _13664_/S vssd1 vssd1 vccd1 vccd1 _13661_/A sky130_fd_sc_hd__mux2_1
X_10872_ _18616_/Q _18951_/Q _10872_/S vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__mux2_1
XFILLER_72_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12611_ _19591_/Q _12697_/A _13004_/A _19523_/Q vssd1 vssd1 vccd1 vccd1 _12611_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13591_ _13591_/A vssd1 vssd1 vccd1 vccd1 _18376_/D sky130_fd_sc_hd__clkbuf_1
XPHY_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15330_ _15387_/S vssd1 vssd1 vccd1 vccd1 _15339_/S sky130_fd_sc_hd__buf_2
XANTENNA__10075__B1 _10074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12542_ hold8/A _12542_/B _12542_/C vssd1 vssd1 vccd1 vccd1 _12542_/X sky130_fd_sc_hd__or3_1
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15261_ _14541_/X _19046_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15262_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13013__B1 _13011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ _12474_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _12473_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18144__A _18144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17000_ _17013_/A vssd1 vssd1 vccd1 vccd1 _17011_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_126_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14212_ _18614_/Q _13965_/X _14220_/S vssd1 vssd1 vccd1 vccd1 _14213_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09766__A _09909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11424_ _11424_/A vssd1 vssd1 vccd1 vccd1 _11424_/Y sky130_fd_sc_hd__inv_2
XFILLER_137_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15192_ _15192_/A vssd1 vssd1 vccd1 vccd1 _19015_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14143_ _18584_/Q _13972_/X _14147_/S vssd1 vssd1 vccd1 vccd1 _14144_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_53_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11355_ _11437_/B vssd1 vssd1 vccd1 vccd1 _11355_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10705__A _10705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12119__A2 _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10306_ _18596_/Q _18867_/Q _19091_/Q _18835_/Q _09682_/A _09712_/A vssd1 vssd1 vccd1
+ vccd1 _10307_/B sky130_fd_sc_hd__mux4_1
X_14074_ _13870_/X _18554_/Q _14074_/S vssd1 vssd1 vccd1 vccd1 _14075_/A sky130_fd_sc_hd__mux2_1
X_18951_ _19329_/CLK _18951_/D vssd1 vssd1 vccd1 vccd1 _18951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11286_ _11070_/X _12447_/B _11192_/Y _12445_/B vssd1 vssd1 vccd1 vccd1 _11465_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_13025_ _14553_/A vssd1 vssd1 vccd1 vccd1 _13025_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17902_ _17478_/X _17454_/X _17901_/X _17646_/A vssd1 vssd1 vccd1 vccd1 _17902_/X
+ sky130_fd_sc_hd__a211o_1
X_10237_ _10250_/A vssd1 vssd1 vccd1 vccd1 _10237_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11878__A1 _11879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18882_ _19268_/CLK _18882_/D vssd1 vssd1 vccd1 vccd1 _18882_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17833_ _17835_/A _17835_/B vssd1 vssd1 vccd1 vccd1 _17833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10168_ _18631_/Q _18966_/Q _10168_/S vssd1 vssd1 vccd1 vccd1 _10169_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17764_ _17768_/B _17215_/X vssd1 vssd1 vccd1 vccd1 _17764_/X sky130_fd_sc_hd__or2b_1
X_14976_ _18934_/Q vssd1 vssd1 vccd1 vccd1 _14977_/A sky130_fd_sc_hd__clkbuf_1
X_10099_ _10108_/A _10099_/B vssd1 vssd1 vccd1 vccd1 _10099_/X sky130_fd_sc_hd__or2_1
XANTENNA__16018__A0 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19503_ _19540_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _19503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16715_ _19548_/Q _19547_/Q _16715_/C _16715_/D vssd1 vssd1 vccd1 vccd1 _16724_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13927_ _13927_/A vssd1 vssd1 vccd1 vccd1 _18507_/D sky130_fd_sc_hd__clkbuf_1
X_17695_ _17693_/X _17694_/Y _17898_/S vssd1 vssd1 vccd1 vccd1 _17695_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15442__S _15444_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19434_ _19583_/CLK _19434_/D vssd1 vssd1 vccd1 vccd1 _19434_/Q sky130_fd_sc_hd__dfxtp_1
X_16646_ _19526_/Q _16644_/B _16590_/X vssd1 vssd1 vccd1 vccd1 _16646_/Y sky130_fd_sc_hd__a21oi_1
X_13858_ _13941_/S vssd1 vssd1 vccd1 vccd1 _13871_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_16_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12809_ _14642_/D _14197_/B vssd1 vssd1 vccd1 vccd1 _13947_/B sky130_fd_sc_hd__nand2_1
XFILLER_16_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19365_ _19365_/CLK _19365_/D vssd1 vssd1 vccd1 vccd1 _19365_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12055__A1 _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16577_ _16714_/A vssd1 vssd1 vccd1 vccd1 _16610_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13789_ _13835_/S vssd1 vssd1 vccd1 vccd1 _13798_/S sky130_fd_sc_hd__buf_2
XFILLER_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ _19663_/CLK _18316_/D vssd1 vssd1 vccd1 vccd1 _18316_/Q sky130_fd_sc_hd__dfxtp_1
X_15528_ _19718_/Q _12651_/X _15543_/S vssd1 vssd1 vccd1 vccd1 _15528_/X sky130_fd_sc_hd__mux2_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_19296_ _19296_/CLK _19296_/D vssd1 vssd1 vccd1 vccd1 _19296_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10161__S0 _09904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__B _17215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13897__S _13903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18247_ input58/X _14274_/X _14277_/X _18234_/X _18146_/A vssd1 vssd1 vccd1 vccd1
+ _18248_/B sky130_fd_sc_hd__a32o_1
XFILLER_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15459_ _19135_/Q _15098_/X _15459_/S vssd1 vssd1 vccd1 vccd1 _15460_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11015__C1 _09465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13555__A1 _13554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09676__A _09676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18178_ _18197_/A vssd1 vssd1 vccd1 vccd1 _18178_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17129_ _11585_/C _09096_/Y _11511_/A _17176_/B _17128_/X vssd1 vssd1 vccd1 vccd1
+ _17130_/D sky130_fd_sc_hd__a2111o_1
XFILLER_144_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10464__S1 _10229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09951_ _10205_/A _09951_/B vssd1 vssd1 vccd1 vccd1 _09951_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09882_ _09952_/S vssd1 vssd1 vccd1 vccd1 _09955_/S sky130_fd_sc_hd__buf_2
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12818__B1 _12704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17133__A _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12046__A1 _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09316_ _11743_/C _11804_/B vssd1 vssd1 vccd1 vccd1 _11551_/B sky130_fd_sc_hd__or2b_2
XFILLER_90_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10152__S0 _09931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ _19833_/Q vssd1 vssd1 vccd1 vccd1 _16623_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13600__S _13609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09178_ _17753_/A _09213_/A vssd1 vssd1 vccd1 vccd1 _17184_/A sky130_fd_sc_hd__nand2_1
XFILLER_147_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10455__S1 _10229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _11254_/A _11140_/B vssd1 vssd1 vccd1 vccd1 _11140_/X sky130_fd_sc_hd__or2_1
Xclkbuf_4_5_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_1_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11071_ _18613_/Q _18948_/Q _11071_/S vssd1 vssd1 vccd1 vccd1 _11072_/B sky130_fd_sc_hd__mux2_1
Xoutput78 _12063_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[16] sky130_fd_sc_hd__buf_2
XANTENNA__14431__S _14439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput89 _12317_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[26] sky130_fd_sc_hd__buf_2
XFILLER_163_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10022_ _10631_/S vssd1 vssd1 vccd1 vccd1 _10022_/X sky130_fd_sc_hd__buf_4
XFILLER_88_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14830_ _18866_/Q _14007_/X _14832_/S vssd1 vssd1 vccd1 vccd1 _14831_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10260__A _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15471__A1 _11120_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input16_A io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14770_/S sky130_fd_sc_hd__buf_4
X_11973_ _11794_/X _11968_/Y _11971_/X _11972_/Y vssd1 vssd1 vccd1 vccd1 _11973_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_17_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14667__A _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16500_ _16501_/B _16501_/C _16499_/Y vssd1 vssd1 vccd1 vccd1 _19484_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13712_ _12981_/X _18425_/Q _13714_/S vssd1 vssd1 vccd1 vccd1 _13713_/A sky130_fd_sc_hd__mux2_1
X_10924_ _10981_/A _10923_/X _09561_/A vssd1 vssd1 vccd1 vccd1 _10924_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_44_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14692_ _14589_/X _18805_/Q _14698_/S vssd1 vssd1 vccd1 vccd1 _14693_/A sky130_fd_sc_hd__mux2_1
X_17480_ _17480_/A vssd1 vssd1 vccd1 vccd1 _17731_/S sky130_fd_sc_hd__buf_2
XFILLER_45_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10391__S0 _10260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16431_ _19461_/Q _16431_/B _16431_/C vssd1 vssd1 vccd1 vccd1 _16433_/B sky130_fd_sc_hd__and3_1
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13643_ _13643_/A vssd1 vssd1 vccd1 vccd1 _18394_/D sky130_fd_sc_hd__clkbuf_1
X_10855_ _10855_/A _10855_/B vssd1 vssd1 vccd1 vccd1 _10855_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10048__B1 _09989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12588__A2 _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19150_ _19688_/CLK _19150_/D vssd1 vssd1 vccd1 vccd1 _19150_/Q sky130_fd_sc_hd__dfxtp_1
X_13574_ _18371_/Q _13573_/X _13577_/S vssd1 vssd1 vccd1 vccd1 _13575_/A sky130_fd_sc_hd__mux2_1
X_16362_ _19435_/Q _16363_/C _19436_/Q vssd1 vssd1 vccd1 vccd1 _16364_/B sky130_fd_sc_hd__a21oi_1
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10786_ _11321_/A _10786_/B vssd1 vssd1 vccd1 vccd1 _10786_/Y sky130_fd_sc_hd__nand2_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18101_ _19815_/Q _18086_/X _18100_/Y _18097_/X vssd1 vssd1 vccd1 vccd1 _19815_/D
+ sky130_fd_sc_hd__o211a_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12525_ _12639_/A vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__clkbuf_2
X_15313_ _14617_/X _19070_/Q _15315_/S vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__mux2_1
X_16293_ _18079_/B vssd1 vssd1 vccd1 vccd1 _16293_/X sky130_fd_sc_hd__buf_4
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19081_ _19081_/CLK _19081_/D vssd1 vssd1 vccd1 vccd1 _19081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14606__S _14615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09496__A _09496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18032_ _19787_/Q _12066_/B _18038_/S vssd1 vssd1 vccd1 vccd1 _18033_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12456_ _12456_/A vssd1 vssd1 vccd1 vccd1 _12456_/X sky130_fd_sc_hd__clkbuf_1
X_15244_ _15244_/A vssd1 vssd1 vccd1 vccd1 _19039_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11407_ _09823_/X _11400_/Y _11402_/Y _11404_/Y _11406_/Y vssd1 vssd1 vccd1 vccd1
+ _11407_/X sky130_fd_sc_hd__o32a_1
XFILLER_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15175_ _15243_/S vssd1 vssd1 vccd1 vccd1 _15184_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12387_ _12387_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12389_/A sky130_fd_sc_hd__nand2_2
XFILLER_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output84_A _12200_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _14182_/A vssd1 vssd1 vccd1 vccd1 _14195_/S sky130_fd_sc_hd__buf_6
XFILLER_153_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11338_ _11331_/Y _11333_/Y _11335_/Y _11337_/Y _09572_/A vssd1 vssd1 vccd1 vccd1
+ _11338_/X sky130_fd_sc_hd__o221a_4
XFILLER_4_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10771__A1 _09434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18934_ _19382_/CLK _18934_/D vssd1 vssd1 vccd1 vccd1 _18934_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14057_ _13845_/X _18546_/Q _14063_/S vssd1 vssd1 vccd1 vccd1 _14058_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14341__S _14343_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11269_ _18577_/Q _18848_/Q _19072_/Q _18816_/Q _10969_/A _09511_/A vssd1 vssd1 vccd1
+ vccd1 _11269_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16239__A0 _13614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13008_ _13008_/A vssd1 vssd1 vccd1 vccd1 _13008_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18865_ _19089_/CLK _18865_/D vssd1 vssd1 vccd1 vccd1 _18865_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11720__A0 _18130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11266__A _11266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15961__A _15983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17816_ _17733_/A _17658_/X _17815_/X _17386_/A vssd1 vssd1 vccd1 vccd1 _17816_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_94_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18796_ _19054_/CLK _18796_/D vssd1 vssd1 vccd1 vccd1 _18796_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15462__A1 _13391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17747_ _17659_/X _17744_/X _17746_/X vssd1 vssd1 vccd1 vccd1 _17747_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14959_ _14959_/A vssd1 vssd1 vccd1 vccd1 _18925_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17678_ _17765_/A _17680_/B _17800_/A _17677_/X vssd1 vssd1 vccd1 vccd1 _17678_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12809__B _14197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19417_ _19699_/CLK _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12028__A1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16629_ _19520_/Q _16634_/B _16628_/Y vssd1 vssd1 vccd1 vccd1 _19520_/D sky130_fd_sc_hd__o21a_1
XFILLER_23_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16792__A _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16962__A1 _16932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19348_ _19357_/CLK _19348_/D vssd1 vssd1 vccd1 vccd1 _19348_/Q sky130_fd_sc_hd__dfxtp_2
X_09101_ _18077_/A _18075_/A _09236_/C _09236_/D vssd1 vssd1 vccd1 vccd1 _11528_/B
+ sky130_fd_sc_hd__and4bb_2
XFILLER_149_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19279_ _19311_/CLK _19279_/D vssd1 vssd1 vccd1 vccd1 _19279_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10685__S1 _10567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11539__A0 _11538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10211__B1 _09909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09934_ _10186_/S vssd1 vssd1 vccd1 vccd1 _10137_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_132_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13161__C1 _13160_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09865_ _10150_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _09865_/X sky130_fd_sc_hd__or2_1
XANTENNA_input8_A io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11176__A _18780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10080__A _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11607__C _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09796_ _11390_/A vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_85_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16178__S _16180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13391__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11904__A _11904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12019__A1 _19406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _10640_/A vssd1 vssd1 vccd1 vccd1 _10705_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_107_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17310__B _17319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ _10571_/A vssd1 vssd1 vccd1 vccd1 _10571_/Y sky130_fd_sc_hd__inv_2
XFILLER_139_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14426__S _14428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12310_ _12310_/A _17867_/B vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__xor2_1
XFILLER_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _19733_/Q _15606_/B _13345_/S vssd1 vssd1 vccd1 vccd1 _13290_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ _12241_/A vssd1 vssd1 vccd1 vccd1 _17305_/A sky130_fd_sc_hd__buf_2
XFILLER_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12742__A2 _12739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12172_ _12122_/A _12122_/B _12148_/A _12171_/Y vssd1 vssd1 vccd1 vccd1 _12173_/B
+ sky130_fd_sc_hd__a31o_2
X_11123_ _11123_/A vssd1 vssd1 vccd1 vccd1 _11173_/S sky130_fd_sc_hd__clkbuf_4
X_16980_ _19646_/Q _16984_/B vssd1 vssd1 vccd1 vccd1 _16980_/X sky130_fd_sc_hd__or2_1
XANTENNA__14161__S _14169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11054_ _18389_/Q _18650_/Q _18549_/Q _18884_/Q _11241_/S _11012_/A vssd1 vssd1 vccd1
+ vccd1 _11055_/B sky130_fd_sc_hd__mux4_1
X_15931_ _13519_/X _19299_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15932_/A sky130_fd_sc_hd__mux2_1
XFILLER_27_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10702__B _12457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10005_ _11335_/A vssd1 vssd1 vccd1 vccd1 _10289_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18650_ _19301_/CLK _18650_/D vssd1 vssd1 vccd1 vccd1 _18650_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15862_ _15862_/A vssd1 vssd1 vccd1 vccd1 _19268_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10600__S1 _09419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16641__B1 _14290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17601_ _17605_/A _17605_/B vssd1 vssd1 vccd1 vccd1 _17601_/Y sky130_fd_sc_hd__nand2_1
X_14813_ _18858_/Q _13981_/X _14821_/S vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__mux2_1
X_18581_ _19076_/CLK _18581_/D vssd1 vssd1 vccd1 vccd1 _18581_/Q sky130_fd_sc_hd__dfxtp_1
X_15793_ _13528_/X _19238_/Q _15793_/S vssd1 vssd1 vccd1 vccd1 _15794_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14397__A _14443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__C1 _09658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13505__S _13507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17532_ _17532_/A vssd1 vssd1 vccd1 vccd1 _17532_/X sky130_fd_sc_hd__buf_2
X_14744_ _14560_/X _18828_/Q _14748_/S vssd1 vssd1 vccd1 vccd1 _14745_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17197__A1 _12219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11956_ _11956_/A _11956_/B vssd1 vssd1 vccd1 vccd1 _11959_/A sky130_fd_sc_hd__and2_1
XFILLER_72_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17463_ _17534_/A _17463_/B vssd1 vssd1 vccd1 vccd1 _17463_/X sky130_fd_sc_hd__or2_1
X_10907_ _18919_/Q _18685_/Q _19367_/Q _19015_/Q _10904_/X _11072_/A vssd1 vssd1 vccd1
+ vccd1 _10907_/X sky130_fd_sc_hd__mux4_1
X_11887_ _11887_/A vssd1 vssd1 vccd1 vccd1 _11962_/A sky130_fd_sc_hd__clkbuf_2
X_14675_ _14675_/A vssd1 vssd1 vccd1 vccd1 _18797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19202_ _19202_/CLK _19202_/D vssd1 vssd1 vccd1 vccd1 _19202_/Q sky130_fd_sc_hd__dfxtp_1
X_16414_ _19454_/Q _16414_/B vssd1 vssd1 vccd1 vccd1 _16415_/B sky130_fd_sc_hd__and2_1
XFILLER_73_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10838_ _18457_/Q _19048_/Q _19210_/Q _18425_/Q _09626_/A _10837_/X vssd1 vssd1 vccd1
+ vccd1 _10839_/B sky130_fd_sc_hd__mux4_1
X_13626_ _13626_/A vssd1 vssd1 vccd1 vccd1 _18386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17394_ _17573_/S vssd1 vssd1 vccd1 vccd1 _17577_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_73_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19133_ _19389_/CLK _19133_/D vssd1 vssd1 vccd1 vccd1 _19133_/Q sky130_fd_sc_hd__dfxtp_1
X_16345_ _19431_/Q _16341_/C _16344_/Y vssd1 vssd1 vccd1 vccd1 _19431_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13557_ _15041_/A vssd1 vssd1 vccd1 vccd1 _13557_/X sky130_fd_sc_hd__clkbuf_2
X_10769_ _10769_/A _10769_/B vssd1 vssd1 vccd1 vccd1 _10769_/X sky130_fd_sc_hd__or2_1
XFILLER_121_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ _19829_/Q _12508_/B _12508_/C _19830_/Q vssd1 vssd1 vccd1 vccd1 _12536_/B
+ sky130_fd_sc_hd__or4b_4
X_19064_ _19471_/CLK _19064_/D vssd1 vssd1 vccd1 vccd1 _19064_/Q sky130_fd_sc_hd__dfxtp_1
X_13488_ _13228_/X _18343_/Q _13492_/S vssd1 vssd1 vccd1 vccd1 _13489_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16276_ _16282_/A _16276_/B vssd1 vssd1 vccd1 vccd1 _16277_/A sky130_fd_sc_hd__and2_1
XFILLER_173_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10992__A1 _18981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18015_ _18015_/A vssd1 vssd1 vccd1 vccd1 _19779_/D sky130_fd_sc_hd__clkbuf_1
X_12439_ _19662_/Q _17020_/A _12416_/B _12438_/Y _12230_/X vssd1 vssd1 vccd1 vccd1
+ _12440_/B sky130_fd_sc_hd__a311o_1
X_15227_ _15227_/A vssd1 vssd1 vccd1 vccd1 _19031_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17647__S _17716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14860__A _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09954__A _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15158_ _15158_/A vssd1 vssd1 vccd1 vccd1 _15167_/S sky130_fd_sc_hd__buf_4
XFILLER_126_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15167__S _15167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _14109_/A vssd1 vssd1 vccd1 vccd1 _14118_/S sky130_fd_sc_hd__buf_4
X_15089_ _15089_/A vssd1 vssd1 vccd1 vccd1 _15089_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18917_ _18917_/CLK _18917_/D vssd1 vssd1 vccd1 vccd1 _18917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18082__C1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _18639_/Q _18974_/Q _10785_/S vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__mux2_1
XFILLER_110_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18848_ _19712_/CLK _18848_/D vssd1 vssd1 vccd1 vccd1 _18848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_0_clock clock vssd1 vssd1 vccd1 vccd1 clkbuf_0_clock/X sky130_fd_sc_hd__clkbuf_16
XFILLER_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09581_ _09760_/A _09555_/X _09573_/X _09833_/A _09580_/Y vssd1 vssd1 vccd1 vccd1
+ _12479_/B sky130_fd_sc_hd__o32a_4
XFILLER_94_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18779_ _19740_/CLK _18779_/D vssd1 vssd1 vccd1 vccd1 _18779_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_leaf_175_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10107__S0 _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10658__S1 _11298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_0_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__11868__A2_N _12454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12185__B1 _15601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15077__S _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09917_ _10158_/A _09916_/X _09823_/A vssd1 vssd1 vccd1 vccd1 _09917_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _10670_/S vssd1 vssd1 vccd1 vccd1 _10546_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09779_ _10381_/S vssd1 vssd1 vccd1 vccd1 _10215_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _19637_/Q _11809_/Y _11810_/S vssd1 vssd1 vccd1 vccd1 _11810_/X sky130_fd_sc_hd__mux2_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12790_ _19588_/Q _12633_/X _12634_/X _19456_/Q _12789_/X vssd1 vssd1 vccd1 vccd1
+ _13399_/B sky130_fd_sc_hd__a221o_4
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10346__S0 _10215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12449__B _12449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11741_ _19635_/Q vssd1 vssd1 vccd1 vccd1 _16951_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16926__A1 _19626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14460_ _14460_/A vssd1 vssd1 vccd1 vccd1 _18715_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ _11618_/A _18114_/A _11672_/S vssd1 vssd1 vccd1 vccd1 _11672_/X sky130_fd_sc_hd__mux2_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13411_ _13411_/A vssd1 vssd1 vccd1 vccd1 _15482_/S sky130_fd_sc_hd__buf_4
X_10623_ _10623_/A vssd1 vssd1 vccd1 vccd1 _11321_/A sky130_fd_sc_hd__clkbuf_4
X_14391_ _13864_/X _18685_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14392_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14156__S _14158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13342_ _19453_/Q _12636_/X _13341_/X vssd1 vssd1 vccd1 vccd1 _13342_/X sky130_fd_sc_hd__o21a_1
X_16130_ _16129_/X _19352_/Q _16140_/S vssd1 vssd1 vccd1 vccd1 _16131_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10554_ _10559_/A _10550_/X _10553_/X _09450_/A vssd1 vssd1 vccd1 vccd1 _10554_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13995__S _13995_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16061_ _16059_/X _19340_/Q _16083_/S vssd1 vssd1 vccd1 vccd1 _16062_/A sky130_fd_sc_hd__mux2_1
X_13273_ _15079_/A vssd1 vssd1 vccd1 vccd1 _14601_/A sky130_fd_sc_hd__clkbuf_2
X_10485_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10485_/Y sky130_fd_sc_hd__nor2_1
X_15012_ _15012_/A vssd1 vssd1 vccd1 vccd1 _15012_/X sky130_fd_sc_hd__clkbuf_2
X_12224_ _12224_/A _12224_/B vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09774__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10726__B2 _10725_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19820_ _19834_/CLK _19820_/D vssd1 vssd1 vccd1 vccd1 _19820_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09592__A1 _09590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ _16989_/A _12156_/C _19650_/Q vssd1 vssd1 vccd1 vccd1 _12155_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_118_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_3_2_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_69_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_193_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19245_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11106_ _18579_/Q _18850_/Q _19074_/Q _18818_/Q _11074_/S _10971_/A vssd1 vssd1 vccd1
+ vccd1 _11106_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19751_ _19756_/CLK _19751_/D vssd1 vssd1 vccd1 vccd1 _19751_/Q sky130_fd_sc_hd__dfxtp_1
X_16963_ _16963_/A _16971_/B vssd1 vssd1 vccd1 vccd1 _16963_/X sky130_fd_sc_hd__or2_1
XFILLER_2_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12086_ _12087_/A _17215_/A vssd1 vssd1 vccd1 vccd1 _12088_/A sky130_fd_sc_hd__and2_1
XANTENNA__11528__B _11528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18702_ _19384_/CLK _18702_/D vssd1 vssd1 vccd1 vccd1 _18702_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15715__S _15721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11037_ _11032_/X _11035_/X _11036_/X _11111_/A _11022_/X vssd1 vssd1 vccd1 vccd1
+ _11044_/B sky130_fd_sc_hd__o221a_1
X_15914_ _19292_/Q _14605_/A _15920_/S vssd1 vssd1 vccd1 vccd1 _15915_/A sky130_fd_sc_hd__mux2_1
X_19682_ _19694_/CLK _19682_/D vssd1 vssd1 vccd1 vccd1 _19682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16894_ _16896_/B _16896_/C _16868_/X vssd1 vssd1 vccd1 vccd1 _16894_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18633_ _18902_/CLK _18633_/D vssd1 vssd1 vccd1 vccd1 _18633_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15845_ _15845_/A vssd1 vssd1 vccd1 vccd1 _19261_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15016__A _15099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18564_ _19285_/CLK _18564_/D vssd1 vssd1 vccd1 vccd1 _18564_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15776_ _13608_/X _19231_/Q _15776_/S vssd1 vssd1 vccd1 vccd1 _15777_/A sky130_fd_sc_hd__mux2_1
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _19561_/Q _12518_/A _12987_/X _13012_/A vssd1 vssd1 vccd1 vccd1 _12988_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _17716_/S _17510_/X _17514_/X vssd1 vssd1 vccd1 vccd1 _17515_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14727_ _14727_/A vssd1 vssd1 vccd1 vccd1 _18820_/D sky130_fd_sc_hd__clkbuf_1
X_11939_ _19642_/Q _19641_/Q _11939_/C vssd1 vssd1 vccd1 vccd1 _11994_/C sky130_fd_sc_hd__and3_1
X_18495_ _18987_/CLK _18495_/D vssd1 vssd1 vccd1 vccd1 _18495_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12651__B2 _18262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10888__S1 _11174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_131_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19759_/CLK sky130_fd_sc_hd__clkbuf_16
X_17446_ _17262_/X _17217_/X _17446_/S vssd1 vssd1 vccd1 vccd1 _17446_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10662__B1 _09602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14658_ _14658_/A vssd1 vssd1 vccd1 vccd1 _18789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13609_ _18382_/Q _13608_/X _13609_/S vssd1 vssd1 vccd1 vccd1 _13610_/A sky130_fd_sc_hd__mux2_1
X_17377_ _17374_/X _17375_/X _17511_/S vssd1 vssd1 vccd1 vccd1 _17377_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14066__S _14074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14589_ _14589_/A vssd1 vssd1 vccd1 vccd1 _14589_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19116_ _19280_/CLK _19116_/D vssd1 vssd1 vccd1 vccd1 _19116_/Q sky130_fd_sc_hd__dfxtp_1
X_16328_ _16331_/B _16331_/C _16293_/X vssd1 vssd1 vccd1 vccd1 _16328_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_158_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16145__A2 _15615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_146_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19712_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19047_ _19241_/CLK _19047_/D vssd1 vssd1 vccd1 vccd1 _19047_/Q sky130_fd_sc_hd__dfxtp_1
X_16259_ _16259_/A vssd1 vssd1 vccd1 vccd1 _19399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12706__A2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09684__A _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10623__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13116__C1 _13234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13667__A0 _13191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09702_ _09840_/S vssd1 vssd1 vccd1 vccd1 _10094_/S sky130_fd_sc_hd__buf_2
XFILLER_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09633_ _18479_/Q _19070_/Q _19232_/Q _18447_/Q _09538_/A _09547_/A vssd1 vssd1 vccd1
+ vccd1 _09634_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17125__B _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09564_ _09803_/A _09558_/X _09820_/A vssd1 vssd1 vccd1 vccd1 _09564_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_130_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09495_ _11151_/S vssd1 vssd1 vccd1 vccd1 _09496_/A sky130_fd_sc_hd__buf_4
XANTENNA__12642__B2 _19339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10879__S1 _10817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09859__A _09859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15592__A0 _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10270_ _10270_/A vssd1 vssd1 vccd1 vccd1 _10272_/A sky130_fd_sc_hd__buf_2
XFILLER_3_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10803__S1 _10802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13960_ _18516_/Q _13959_/X _13963_/S vssd1 vssd1 vccd1 vccd1 _13961_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12911_ _19745_/Q vssd1 vssd1 vccd1 vccd1 _16021_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_86_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13891_ _13889_/X _18496_/Q _13903_/S vssd1 vssd1 vccd1 vccd1 _13892_/A sky130_fd_sc_hd__mux2_1
X_15630_ hold7/A _13359_/X _15629_/Y _12544_/X vssd1 vssd1 vccd1 vccd1 _15630_/X sky130_fd_sc_hd__o211a_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ _19590_/Q _12697_/X _12503_/A _19458_/Q _12841_/X vssd1 vssd1 vccd1 vccd1
+ _13415_/B sky130_fd_sc_hd__a221o_4
XFILLER_46_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15561_/A vssd1 vssd1 vccd1 vccd1 _19155_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _12773_/A vssd1 vssd1 vccd1 vccd1 _12773_/X sky130_fd_sc_hd__buf_2
XFILLER_42_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15270__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17300_ _17550_/S vssd1 vssd1 vccd1 vccd1 _17653_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14512_ _14512_/A vssd1 vssd1 vccd1 vccd1 _18739_/D sky130_fd_sc_hd__clkbuf_1
X_11724_ _11782_/B vssd1 vssd1 vccd1 vccd1 _17391_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18280_ _19731_/CLK _18280_/D vssd1 vssd1 vccd1 vccd1 _18280_/Q sky130_fd_sc_hd__dfxtp_1
X_15492_ _15492_/A vssd1 vssd1 vccd1 vccd1 _19143_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17410_/B _12405_/A _17251_/S vssd1 vssd1 vccd1 vccd1 _17231_/X sky130_fd_sc_hd__mux2_1
X_11655_ _19330_/Q _11653_/X _15488_/A vssd1 vssd1 vccd1 vccd1 _11655_/Y sky130_fd_sc_hd__o21ai_1
X_14443_ _13940_/X _18709_/Q _14443_/S vssd1 vssd1 vccd1 vccd1 _14444_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_63_clock clkbuf_opt_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19540_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_156_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12195__A _12195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16890__A _16890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _18589_/Q _18860_/Q _19084_/Q _18828_/Q _10763_/S _09590_/X vssd1 vssd1 vccd1
+ vccd1 _10606_/X sky130_fd_sc_hd__mux4_1
X_17162_ _17175_/A _17149_/X _17140_/A _19706_/Q vssd1 vssd1 vccd1 vccd1 _17163_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11586_ _17165_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11586_/Y sky130_fd_sc_hd__nor2_1
X_14374_ _14430_/A vssd1 vssd1 vccd1 vccd1 _14443_/S sky130_fd_sc_hd__buf_6
XFILLER_167_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16113_ _16113_/A vssd1 vssd1 vccd1 vccd1 _19349_/D sky130_fd_sc_hd__clkbuf_1
X_13325_ _16912_/B _13260_/X _13261_/X _16501_/B _13324_/X vssd1 vssd1 vccd1 vccd1
+ _13325_/X sky130_fd_sc_hd__a221o_4
X_10537_ _10277_/A _10536_/X _10297_/A vssd1 vssd1 vccd1 vccd1 _10537_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_123_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17093_ _17093_/A vssd1 vssd1 vccd1 vccd1 _19692_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12923__A _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_78_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19725_/CLK sky130_fd_sc_hd__clkbuf_16
X_16044_ _16044_/A vssd1 vssd1 vccd1 vccd1 _19337_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10468_ _09727_/A _10461_/X _10463_/X _10467_/X _09753_/A vssd1 vssd1 vccd1 vccd1
+ _10468_/X sky130_fd_sc_hd__a311o_4
XANTENNA__11047__S1 _10990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13256_ _19763_/Q _19764_/Q _13256_/C vssd1 vssd1 vccd1 vccd1 _13281_/B sky130_fd_sc_hd__and3_1
XFILLER_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12207_ _19413_/Q _12093_/X _12203_/X _12206_/Y vssd1 vssd1 vccd1 vccd1 _16290_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_123_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13187_ _13154_/X _13186_/X _13164_/X vssd1 vssd1 vccd1 vccd1 _13187_/Y sky130_fd_sc_hd__a21oi_1
X_10399_ _09761_/A _10388_/X _10397_/X _09834_/A _10398_/Y vssd1 vssd1 vccd1 vccd1
+ _12466_/B sky130_fd_sc_hd__o32a_4
X_19803_ _19845_/CLK _19803_/D vssd1 vssd1 vccd1 vccd1 _19803_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12138_ _12020_/X _12467_/B _12137_/Y vssd1 vssd1 vccd1 vccd1 _17790_/A sky130_fd_sc_hd__a21oi_4
XFILLER_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17995_ _17995_/A vssd1 vssd1 vccd1 vccd1 _19770_/D sky130_fd_sc_hd__clkbuf_1
X_16946_ _16946_/A vssd1 vssd1 vccd1 vccd1 _16970_/A sky130_fd_sc_hd__clkbuf_2
X_12069_ _12274_/B vssd1 vssd1 vccd1 vccd1 _12069_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19734_ _19734_/CLK _19734_/D vssd1 vssd1 vccd1 vccd1 _19734_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__10558__S0 _10763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19665_ _19668_/CLK _19665_/D vssd1 vssd1 vccd1 vccd1 _19665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16877_ _16879_/B _16879_/C _16868_/X vssd1 vssd1 vccd1 vccd1 _16877_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11675__A2 _12445_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17260__A0 _17215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18616_ _19365_/CLK _18616_/D vssd1 vssd1 vccd1 vccd1 _18616_/Q sky130_fd_sc_hd__dfxtp_1
X_15828_ _15839_/A vssd1 vssd1 vccd1 vccd1 _15837_/S sky130_fd_sc_hd__buf_6
Xclkbuf_leaf_16_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19387_/CLK sky130_fd_sc_hd__clkbuf_16
X_19596_ _19598_/CLK _19596_/D vssd1 vssd1 vccd1 vccd1 _19596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_48_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18547_ _19300_/CLK _18547_/D vssd1 vssd1 vccd1 vccd1 _18547_/Q sky130_fd_sc_hd__dfxtp_1
X_15759_ _13583_/X _19223_/Q _15765_/S vssd1 vssd1 vccd1 vccd1 _15760_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15180__S _15184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09280_ _12817_/A _16937_/B _09280_/C _09280_/D vssd1 vssd1 vccd1 vccd1 _09280_/X
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__09679__A _09980_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18478_ _19261_/CLK _18478_/D vssd1 vssd1 vccd1 vccd1 _18478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17429_ _17994_/S vssd1 vssd1 vccd1 vccd1 _17831_/A sky130_fd_sc_hd__buf_2
XFILLER_147_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16118__A2 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__S1 _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11838__A1_N _11890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10353__A _19726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_125_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15355__S _15361_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10469__A3 _10468_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__S _10499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12863__B2 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11184__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09616_ _09369_/A _09604_/X _09615_/X _09472_/A _19737_/Q vssd1 vssd1 vccd1 vccd1
+ _11413_/A sky130_fd_sc_hd__a32o_4
XFILLER_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13812__A0 _13191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ _09547_/A vssd1 vssd1 vccd1 vccd1 _09547_/X sky130_fd_sc_hd__buf_2
XFILLER_169_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15090__S _15093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13603__S _13609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09617_/A vssd1 vssd1 vccd1 vccd1 _09760_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10641__A3 _18828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11440_ _11443_/A _11446_/A _11443_/C _10402_/A vssd1 vssd1 vccd1 vccd1 _11440_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11277__S1 _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11051__B1 _11254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13839__A _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10962__S _10962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _11364_/X _11366_/X _11368_/X _11370_/X _09754_/X vssd1 vssd1 vccd1 vccd1
+ _11371_/X sky130_fd_sc_hd__a221o_1
XFILLER_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ _19317_/Q _18729_/Q _18766_/Q _18340_/Q _09682_/A _10314_/A vssd1 vssd1 vccd1
+ vccd1 _10323_/B sky130_fd_sc_hd__mux4_1
X_13110_ _13110_/A vssd1 vssd1 vccd1 vccd1 _18298_/D sky130_fd_sc_hd__clkbuf_1
X_14090_ _13893_/X _18561_/Q _14096_/S vssd1 vssd1 vccd1 vccd1 _14091_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13041_ _19719_/Q _12667_/B _13143_/S vssd1 vssd1 vccd1 vccd1 _13041_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10253_ _19286_/Q _19124_/Q _18533_/Q _18303_/Q _10247_/X _10238_/X vssd1 vssd1 vccd1
+ vccd1 _10254_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10263__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10788__S0 _09519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input46_A io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _10184_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10184_/X sky130_fd_sc_hd__or2_1
XFILLER_105_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16800_ _19573_/Q _16800_/B _16800_/C vssd1 vssd1 vccd1 vccd1 _16809_/D sky130_fd_sc_hd__and3_1
XFILLER_121_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17780_ _17726_/A _17726_/B _17777_/B _17779_/X vssd1 vssd1 vccd1 vccd1 _17780_/X
+ sky130_fd_sc_hd__o31a_1
X_14992_ _18942_/Q vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16731_ _19553_/Q _16731_/B _16731_/C vssd1 vssd1 vccd1 vccd1 _16736_/C sky130_fd_sc_hd__and3_1
XFILLER_120_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13943_ _14519_/A vssd1 vssd1 vccd1 vccd1 _13943_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19450_ _19550_/CLK _19450_/D vssd1 vssd1 vccd1 vccd1 _19450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16662_ _19530_/Q _16669_/D vssd1 vssd1 vccd1 vccd1 _16664_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13874_ _13941_/S vssd1 vssd1 vccd1 vccd1 _13887_/S sky130_fd_sc_hd__buf_2
XFILLER_75_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18401_ _19314_/CLK _18401_/D vssd1 vssd1 vccd1 vccd1 _18401_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10960__S0 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15613_ _15613_/A vssd1 vssd1 vccd1 vccd1 _15613_/Y sky130_fd_sc_hd__inv_2
X_19381_ _19502_/CLK _19381_/D vssd1 vssd1 vccd1 vccd1 _19381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12825_ _19740_/Q _12824_/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12825_/X sky130_fd_sc_hd__mux2_1
X_16593_ _16890_/A vssd1 vssd1 vccd1 vccd1 _16806_/A sky130_fd_sc_hd__buf_2
XFILLER_62_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14609__S _14615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18332_ _19245_/CLK _18332_/D vssd1 vssd1 vccd1 vccd1 _18332_/Q sky130_fd_sc_hd__dfxtp_1
X_15544_ _15543_/X _19152_/Q _15544_/S vssd1 vssd1 vccd1 vccd1 _15545_/A sky130_fd_sc_hd__mux2_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09499__A _10633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ hold10/A _12752_/X _11347_/A _12755_/X vssd1 vssd1 vccd1 vccd1 _18266_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_43_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12082__A2 _12465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15556__A0 _19723_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _16947_/A _11706_/B _11706_/C vssd1 vssd1 vccd1 vccd1 _11707_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _19720_/CLK _18263_/D vssd1 vssd1 vccd1 vccd1 _18263_/Q sky130_fd_sc_hd__dfxtp_2
X_15475_ _19710_/Q _16024_/S _13423_/B vssd1 vssd1 vccd1 vccd1 _15475_/X sky130_fd_sc_hd__a21o_1
X_12687_ _18274_/Q _12687_/B vssd1 vssd1 vccd1 vccd1 _12687_/X sky130_fd_sc_hd__or2_1
XFILLER_147_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17214_ _17214_/A vssd1 vssd1 vccd1 vccd1 _17722_/B sky130_fd_sc_hd__clkbuf_2
X_14426_ _13915_/X _18701_/Q _14428_/S vssd1 vssd1 vccd1 vccd1 _14427_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18194_ input37/X _18178_/X _18188_/X _18193_/X _17114_/A vssd1 vssd1 vccd1 vccd1
+ _18195_/B sky130_fd_sc_hd__a32o_1
X_11638_ _11638_/A _11638_/B vssd1 vssd1 vccd1 vccd1 _11639_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11268__S1 _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17145_ _17145_/A _17145_/B _17145_/C _17145_/D vssd1 vssd1 vccd1 vccd1 _17145_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13749__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10872__S _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14357_ _13921_/X _18671_/Q _14365_/S vssd1 vssd1 vccd1 vccd1 _14358_/A sky130_fd_sc_hd__mux2_1
XFILLER_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ _11569_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _17175_/C sky130_fd_sc_hd__and2_1
XFILLER_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13308_ _12848_/A _13299_/Y _13307_/X _13051_/A vssd1 vssd1 vccd1 vccd1 _13308_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_144_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17076_ _17076_/A vssd1 vssd1 vccd1 vccd1 _19684_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14288_ _14288_/A vssd1 vssd1 vccd1 vccd1 _18643_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16027_ _19746_/Q _16028_/B vssd1 vssd1 vccd1 vccd1 _16039_/C sky130_fd_sc_hd__or2_2
X_13239_ _15073_/A vssd1 vssd1 vccd1 vccd1 _14595_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09633__S1 _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16284__A1 _12126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17978_ _17978_/A vssd1 vssd1 vccd1 vccd1 _19762_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13098__B2 _19343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16929_ input69/X _16929_/B vssd1 vssd1 vccd1 vccd1 _16929_/X sky130_fd_sc_hd__or2_1
XFILLER_37_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19717_ _19720_/CLK _19717_/D vssd1 vssd1 vccd1 vccd1 _19717_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_38_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15903__S _15909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10112__S _10112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19648_ _19649_/CLK _19648_/D vssd1 vssd1 vccd1 vccd1 _19648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09401_ _18781_/Q vssd1 vssd1 vccd1 vccd1 _11211_/A sky130_fd_sc_hd__inv_2
X_19579_ _19581_/CLK _19579_/D vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09332_ _19855_/Q vssd1 vssd1 vccd1 vccd1 _09351_/A sky130_fd_sc_hd__buf_4
XFILLER_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17536__A1 _11512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13270__A1 _15598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09263_ _19826_/Q _19825_/Q _19823_/Q _19824_/Q vssd1 vssd1 vccd1 vccd1 _09270_/A
+ sky130_fd_sc_hd__or4b_1
X_09194_ _19851_/Q vssd1 vssd1 vccd1 vccd1 _09194_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13022__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09872__S1 _09871_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkbuf_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__11907__A _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12836__B2 _19330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15813__S _15815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _18487_/Q _18982_/Q _10940_/S vssd1 vssd1 vccd1 vccd1 _10940_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17775__A1 _17779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__S0 _11172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10871_ _11184_/A _10871_/B vssd1 vssd1 vccd1 vccd1 _10871_/X sky130_fd_sc_hd__or2_1
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_1_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__12738__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12610_ _19331_/Q _12600_/Y _12604_/X _12609_/X vssd1 vssd1 vccd1 vccd1 _12610_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15114__A _15171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ _18376_/Q _13589_/X _13593_/S vssd1 vssd1 vccd1 vccd1 _13591_/A sky130_fd_sc_hd__mux2_1
XPHY_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12457__B _12457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10075__A1 _10684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12541_ _19536_/Q _12507_/X _12511_/X _19504_/Q _12540_/X vssd1 vssd1 vccd1 vccd1
+ _12542_/C sky130_fd_sc_hd__a221o_4
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13013__A1 _19562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15260_ _15260_/A vssd1 vssd1 vccd1 vccd1 _19045_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12472_ _12474_/A _12472_/B vssd1 vssd1 vccd1 vccd1 _12472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14211_ _14268_/S vssd1 vssd1 vccd1 vccd1 _14220_/S sky130_fd_sc_hd__buf_2
XANTENNA__10692__S _10692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ _11423_/A vssd1 vssd1 vccd1 vccd1 _11423_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15191_ _19015_/Q _15022_/X _15195_/S vssd1 vssd1 vccd1 vccd1 _15192_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12772__B1 _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14142_ _14142_/A vssd1 vssd1 vccd1 vccd1 _18583_/D sky130_fd_sc_hd__clkbuf_1
X_11354_ _11354_/A _12470_/B vssd1 vssd1 vccd1 vccd1 _11437_/B sky130_fd_sc_hd__nand2_1
XFILLER_153_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11089__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _10305_/A vssd1 vssd1 vccd1 vccd1 _11439_/A sky130_fd_sc_hd__inv_2
XFILLER_125_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15784__A _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14073_ _14073_/A vssd1 vssd1 vccd1 vccd1 _18553_/D sky130_fd_sc_hd__clkbuf_1
X_11285_ _11239_/Y _11465_/D _11284_/Y vssd1 vssd1 vccd1 vccd1 _11285_/X sky130_fd_sc_hd__a21o_1
X_18950_ _19329_/CLK _18950_/D vssd1 vssd1 vccd1 vccd1 _18950_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_153_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10236_ _10236_/A vssd1 vssd1 vccd1 vccd1 _10250_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13024_ _15031_/A vssd1 vssd1 vccd1 vccd1 _14553_/A sky130_fd_sc_hd__clkbuf_2
X_17901_ _17466_/X _17898_/X _17900_/Y _17532_/A vssd1 vssd1 vccd1 vccd1 _17901_/X
+ sky130_fd_sc_hd__o211a_1
X_18881_ _19298_/CLK _18881_/D vssd1 vssd1 vccd1 vccd1 _18881_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output152_A _16286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11817__A _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17832_ _17835_/A _17835_/B _17832_/S vssd1 vssd1 vccd1 vccd1 _17832_/X sky130_fd_sc_hd__mux2_1
X_10167_ _10167_/A vssd1 vssd1 vccd1 vccd1 _10167_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17763_ _10491_/Y _17652_/X _17762_/X vssd1 vssd1 vccd1 vccd1 _19723_/D sky130_fd_sc_hd__a21oi_1
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14975_ _14975_/A vssd1 vssd1 vccd1 vccd1 _18933_/D sky130_fd_sc_hd__clkbuf_1
X_10098_ _18408_/Q _18669_/Q _18568_/Q _18903_/Q _10137_/S _09714_/A vssd1 vssd1 vccd1
+ vccd1 _10099_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16714_ _16714_/A vssd1 vssd1 vccd1 vccd1 _16762_/A sky130_fd_sc_hd__clkbuf_4
X_19502_ _19502_/CLK _19502_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_2
X_13926_ _13925_/X _18507_/Q _13935_/S vssd1 vssd1 vccd1 vccd1 _13927_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17694_ _17696_/A _17696_/B vssd1 vssd1 vccd1 vccd1 _17694_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19433_ _19583_/CLK _19433_/D vssd1 vssd1 vccd1 vccd1 _19433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16645_ _19525_/Q _16642_/A _16644_/Y vssd1 vssd1 vccd1 vccd1 _19525_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13857_ _14537_/A vssd1 vssd1 vccd1 vccd1 _13857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14339__S _14343_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11552__A _16000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ _19814_/Q vssd1 vssd1 vccd1 vccd1 _14642_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19364_ _19364_/CLK _19364_/D vssd1 vssd1 vccd1 vccd1 _19364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16576_ _16585_/A _16576_/B _16578_/B vssd1 vssd1 vccd1 vccd1 _19506_/D sky130_fd_sc_hd__nor3_1
XFILLER_50_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13788_ _13788_/A vssd1 vssd1 vccd1 vccd1 _18458_/D sky130_fd_sc_hd__clkbuf_1
X_18315_ _19663_/CLK _18315_/D vssd1 vssd1 vccd1 vccd1 _18315_/Q sky130_fd_sc_hd__dfxtp_1
X_15527_ _15527_/A vssd1 vssd1 vccd1 vccd1 _19148_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12739_ _12744_/A vssd1 vssd1 vccd1 vccd1 _12739_/X sky130_fd_sc_hd__buf_6
X_19295_ _19389_/CLK _19295_/D vssd1 vssd1 vccd1 vccd1 _19295_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11702__D _11702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10161__S1 _09888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18246_ _18246_/A vssd1 vssd1 vccd1 vccd1 _19865_/D sky130_fd_sc_hd__clkbuf_1
X_15458_ _15458_/A vssd1 vssd1 vccd1 vccd1 _19134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09759__A1 _09667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ _13889_/X _18693_/Q _14417_/S vssd1 vssd1 vccd1 vccd1 _14410_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18177_ _18177_/A vssd1 vssd1 vccd1 vccd1 _19842_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14074__S _14074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09759__B2 _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15389_ _15854_/B _15389_/B vssd1 vssd1 vccd1 vccd1 _15446_/A sky130_fd_sc_hd__nor2_4
XANTENNA__12383__A _12383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11110__S0 _09624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12763__B1 _10303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17128_ _17114_/A _09210_/X _17115_/X _17127_/Y vssd1 vssd1 vccd1 vccd1 _17128_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_171_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09950_ _18936_/Q _18702_/Q _19384_/Q _19032_/Q _10112_/S _10218_/A vssd1 vssd1 vccd1
+ vccd1 _09951_/B sky130_fd_sc_hd__mux4_1
X_17059_ _19677_/Q _15536_/X _17061_/S vssd1 vssd1 vccd1 vccd1 _17060_/A sky130_fd_sc_hd__mux2_1
XFILLER_104_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09881_ _10341_/S vssd1 vssd1 vccd1 vccd1 _09952_/S sky130_fd_sc_hd__clkbuf_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__A2 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16302__B _16302_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16009__A1 _19331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17206__A0 _17662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15633__S _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17133__B _17133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13243__A1 input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09315_ _19696_/Q _09315_/B vssd1 vssd1 vccd1 vccd1 _11804_/B sky130_fd_sc_hd__nand2_1
XFILLER_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18182__B2 _19844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__S1 _09871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ _19834_/Q vssd1 vssd1 vccd1 vccd1 _16623_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13389__A _17028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15940__A0 _13531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _11589_/A _09208_/A _11556_/B _17108_/B vssd1 vssd1 vccd1 vccd1 _09213_/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12293__A _19417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12754__B1 _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17693__A0 _17696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10017__S _10017_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _09367_/A _11057_/X _11069_/X _09470_/A _19711_/Q vssd1 vssd1 vccd1 vccd1
+ _11070_/X sky130_fd_sc_hd__a32o_2
XFILLER_131_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput79 _12092_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[17] sky130_fd_sc_hd__buf_2
XFILLER_89_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10021_ _18411_/Q _18672_/Q _18571_/Q _18906_/Q _09776_/A _10056_/A vssd1 vssd1 vccd1
+ vccd1 _10021_/X sky130_fd_sc_hd__mux4_1
XFILLER_102_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10541__A _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14760_ _14760_/A vssd1 vssd1 vccd1 vccd1 _18835_/D sky130_fd_sc_hd__clkbuf_1
X_11972_ _19340_/Q _11653_/X _16114_/A vssd1 vssd1 vccd1 vccd1 _11972_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13711_ _13711_/A vssd1 vssd1 vccd1 vccd1 _18424_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10923_ _19305_/Q _18717_/Q _18754_/Q _18328_/Q _10852_/S _10837_/A vssd1 vssd1 vccd1
+ vccd1 _10923_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11493__B1 _18100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14691_ _14691_/A vssd1 vssd1 vccd1 vccd1 _18804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10391__S1 _10436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16430_ _16431_/B _16431_/C _16429_/Y vssd1 vssd1 vccd1 vccd1 _19460_/D sky130_fd_sc_hd__o21a_1
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13642_ _12999_/X _18394_/Q _13642_/S vssd1 vssd1 vccd1 vccd1 _13643_/A sky130_fd_sc_hd__mux2_1
X_10854_ _18617_/Q _18952_/Q _10854_/S vssd1 vssd1 vccd1 vccd1 _10855_/B sky130_fd_sc_hd__mux2_1
XFILLER_32_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16361_ _19435_/Q _16363_/C _16360_/Y vssd1 vssd1 vccd1 vccd1 _19435_/D sky130_fd_sc_hd__o21a_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _15057_/A vssd1 vssd1 vccd1 vccd1 _13573_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10785_ _18618_/Q _18953_/Q _10785_/S vssd1 vssd1 vccd1 vccd1 _10786_/B sky130_fd_sc_hd__mux2_1
X_18100_ _18100_/A _18128_/B vssd1 vssd1 vccd1 vccd1 _18100_/Y sky130_fd_sc_hd__nand2_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15312_ _15312_/A vssd1 vssd1 vccd1 vccd1 _19069_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ _13391_/A _12955_/B vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__and2_1
X_19080_ _19113_/CLK _19080_/D vssd1 vssd1 vccd1 vccd1 _19080_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16292_ _19414_/Q vssd1 vssd1 vccd1 vccd1 _16292_/Y sky130_fd_sc_hd__inv_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18031_ _18031_/A vssd1 vssd1 vccd1 vccd1 _19786_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15931__A0 _13519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15243_ _19039_/Q _15098_/X _15243_/S vssd1 vssd1 vccd1 vccd1 _15244_/A sky130_fd_sc_hd__mux2_1
X_12455_ _12462_/B _12455_/B vssd1 vssd1 vccd1 vccd1 _12456_/A sky130_fd_sc_hd__and2b_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12745__B1 _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11406_ _11402_/A _11405_/X _09823_/X vssd1 vssd1 vccd1 vccd1 _11406_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15174_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15243_/S sky130_fd_sc_hd__buf_4
X_12386_ _12386_/A vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__inv_2
XFILLER_126_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14125_ _15854_/A _15317_/B vssd1 vssd1 vccd1 vccd1 _14182_/A sky130_fd_sc_hd__nor2_2
XFILLER_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _10779_/A _11336_/X _09484_/A vssd1 vssd1 vccd1 vccd1 _11337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_114_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14498__A0 _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18933_ _19502_/CLK _18933_/D vssd1 vssd1 vccd1 vccd1 _18933_/Q sky130_fd_sc_hd__dfxtp_1
X_14056_ _14056_/A vssd1 vssd1 vccd1 vccd1 _18545_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output77_A _12035_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ _18385_/Q _18646_/Q _18545_/Q _18880_/Q _11112_/X _10910_/A vssd1 vssd1 vccd1
+ vccd1 _11268_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12650__B _18262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13007_ _13179_/A vssd1 vssd1 vccd1 vccd1 _13007_/X sky130_fd_sc_hd__clkbuf_2
X_10219_ _09773_/A _10216_/Y _10218_/Y _10214_/A vssd1 vssd1 vccd1 vccd1 _10219_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15019__A _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18864_ _19088_/CLK _18864_/D vssd1 vssd1 vccd1 vccd1 _18864_/Q sky130_fd_sc_hd__dfxtp_1
X_11199_ _10937_/A _11196_/X _11198_/X vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__a21o_1
XFILLER_121_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11181__C1 _10883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11720__A1 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17815_ _17419_/X _17656_/X _17814_/Y _17852_/A vssd1 vssd1 vccd1 vccd1 _17815_/X
+ sky130_fd_sc_hd__o211a_1
X_18795_ _19245_/CLK _18795_/D vssd1 vssd1 vccd1 vccd1 _18795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11159__S0 _10904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15453__S _15455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17746_ _17743_/A _17743_/B _17672_/A _17745_/Y vssd1 vssd1 vccd1 vccd1 _17746_/X
+ sky130_fd_sc_hd__o211a_1
X_14958_ _18925_/Q vssd1 vssd1 vccd1 vccd1 _14959_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_36_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _14589_/A vssd1 vssd1 vccd1 vccd1 _13909_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17677_ _17917_/A _17680_/A vssd1 vssd1 vccd1 vccd1 _17677_/X sky130_fd_sc_hd__or2_1
XFILLER_35_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14889_ _18892_/Q _13988_/X _14893_/S vssd1 vssd1 vccd1 vccd1 _14890_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16628_ _19520_/Q _16634_/B _16590_/X vssd1 vssd1 vccd1 vccd1 _16628_/Y sky130_fd_sc_hd__a21oi_1
X_19416_ _19416_/CLK _19416_/D vssd1 vssd1 vccd1 vccd1 _19416_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__14422__A0 _13909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13225__A1 input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12097__B _19406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10039__A1 _10046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16559_ _19500_/Q hold3/X _16559_/C vssd1 vssd1 vccd1 vccd1 _16561_/B sky130_fd_sc_hd__and3_1
X_19347_ _19349_/CLK _19347_/D vssd1 vssd1 vccd1 vccd1 _19347_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_149_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09100_ _19835_/Q vssd1 vssd1 vccd1 vccd1 _09236_/D sky130_fd_sc_hd__clkbuf_2
XANTENNA__13701__S _13703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19278_ _19278_/CLK _19278_/D vssd1 vssd1 vccd1 vccd1 _19278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17911__A1 _17907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18229_ _18229_/A vssd1 vssd1 vccd1 vccd1 _18229_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_164_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12736__A0 _18255_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__A1 _17166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_171_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14532__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09933_ _09733_/A _09930_/X _09932_/X vssd1 vssd1 vccd1 vccd1 _09933_/X sky130_fd_sc_hd__a21o_1
XFILLER_131_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ _19323_/Q _18735_/Q _18772_/Q _18346_/Q _09846_/X _09839_/A vssd1 vssd1 vccd1
+ vccd1 _09865_/B sky130_fd_sc_hd__mux4_1
XFILLER_113_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10070__S0 _09500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09964_/A vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10080__B _12477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17144__A _17163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13391__B _13391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16983__A _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_96_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16194__S _16202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14707__S _14709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10570_ _18495_/Q _18990_/Q _11320_/S vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16166__B1 _13430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09229_ _11573_/A vssd1 vssd1 vccd1 vccd1 _11508_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12240_ _12240_/A vssd1 vssd1 vccd1 vccd1 _17835_/A sky130_fd_sc_hd__clkinv_2
XFILLER_108_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10202__A1 _09844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _12118_/A _12146_/A _12170_/Y vssd1 vssd1 vccd1 vccd1 _12171_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_135_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12751__A _12751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _18779_/Q vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__buf_2
XANTENNA__12470__B _12470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11053_ _18581_/Q _18852_/Q _19076_/Q _18820_/Q _10940_/S _11005_/X vssd1 vssd1 vccd1
+ vccd1 _11053_/X sky130_fd_sc_hd__mux4_1
X_15930_ _15930_/A vssd1 vssd1 vccd1 vccd1 _19298_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10004_ _10014_/A _10004_/B vssd1 vssd1 vccd1 vccd1 _10004_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10061__S0 _09500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ _19268_/Q _14528_/A _15865_/S vssd1 vssd1 vccd1 vccd1 _15862_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14678__A _14700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17600_ _17605_/A _17605_/B _17775_/S vssd1 vssd1 vccd1 vccd1 _17600_/X sky130_fd_sc_hd__mux2_1
X_14812_ _14858_/S vssd1 vssd1 vccd1 vccd1 _14821_/S sky130_fd_sc_hd__buf_2
X_18580_ _19074_/CLK _18580_/D vssd1 vssd1 vccd1 vccd1 _18580_/Q sky130_fd_sc_hd__dfxtp_1
X_15792_ _15792_/A vssd1 vssd1 vccd1 vccd1 _19237_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17531_ _17672_/A vssd1 vssd1 vccd1 vccd1 _17532_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14743_ _14743_/A vssd1 vssd1 vccd1 vccd1 _18827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11955_ _11955_/A _17221_/A vssd1 vssd1 vccd1 vccd1 _11956_/B sky130_fd_sc_hd__or2_1
XFILLER_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ _11220_/A vssd1 vssd1 vccd1 vccd1 _11072_/A sky130_fd_sc_hd__clkbuf_4
X_17462_ _17462_/A vssd1 vssd1 vccd1 vccd1 _17462_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_44_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14674_ _14563_/X _18797_/Q _14676_/S vssd1 vssd1 vccd1 vccd1 _14675_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11886_ _19640_/Q _19639_/Q _11886_/C vssd1 vssd1 vccd1 vccd1 _11939_/C sky130_fd_sc_hd__and3_1
XFILLER_33_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16413_ _19453_/Q _16409_/B _16412_/Y vssd1 vssd1 vccd1 vccd1 _19453_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19201_ _19201_/CLK _19201_/D vssd1 vssd1 vccd1 vccd1 _19201_/Q sky130_fd_sc_hd__dfxtp_1
X_13625_ _12828_/X _18386_/Q _13631_/S vssd1 vssd1 vccd1 vccd1 _13626_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10837_ _10837_/A vssd1 vssd1 vccd1 vccd1 _10837_/X sky130_fd_sc_hd__buf_2
X_17393_ _17393_/A vssd1 vssd1 vccd1 vccd1 _17573_/S sky130_fd_sc_hd__clkbuf_2
X_19132_ _19326_/CLK _19132_/D vssd1 vssd1 vccd1 vccd1 _19132_/Q sky130_fd_sc_hd__dfxtp_1
X_16344_ _16344_/A _16351_/C vssd1 vssd1 vccd1 vccd1 _16344_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15302__A _15302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ _13556_/A vssd1 vssd1 vccd1 vccd1 _18365_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10768_ _18394_/Q _18655_/Q _18554_/Q _18889_/Q _11297_/S _09600_/A vssd1 vssd1 vccd1
+ vccd1 _10769_/B sky130_fd_sc_hd__mux4_1
XFILLER_146_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12507_ _13004_/A vssd1 vssd1 vccd1 vccd1 _12507_/X sky130_fd_sc_hd__buf_2
X_19063_ _19382_/CLK _19063_/D vssd1 vssd1 vccd1 vccd1 _19063_/Q sky130_fd_sc_hd__dfxtp_1
X_16275_ _16275_/A vssd1 vssd1 vccd1 vccd1 _19406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13487_ _13487_/A vssd1 vssd1 vccd1 vccd1 _18342_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10699_ _10074_/X _10689_/Y _10694_/X _10698_/Y _09658_/X vssd1 vssd1 vccd1 vccd1
+ _10699_/X sky130_fd_sc_hd__o311a_1
X_18014_ _19779_/Q _11879_/A _18016_/S vssd1 vssd1 vccd1 vccd1 _18015_/A sky130_fd_sc_hd__mux2_1
X_15226_ _19031_/Q _15073_/X _15228_/S vssd1 vssd1 vccd1 vccd1 _15227_/A sky130_fd_sc_hd__mux2_1
X_12438_ _17020_/A _12416_/B _19662_/Q vssd1 vssd1 vccd1 vccd1 _12438_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14860__B _14860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15157_ _15157_/A vssd1 vssd1 vccd1 vccd1 _19000_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14352__S _14354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12369_ _12369_/A _12369_/B vssd1 vssd1 vccd1 vccd1 _12369_/Y sky130_fd_sc_hd__nand2_1
XFILLER_99_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11941__A1 _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14108_ _14108_/A vssd1 vssd1 vccd1 vccd1 _18569_/D sky130_fd_sc_hd__clkbuf_1
X_15088_ _15088_/A vssd1 vssd1 vccd1 vccd1 _18971_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13143__A0 _19725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15972__A _15983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18916_ _19012_/CLK _18916_/D vssd1 vssd1 vccd1 vccd1 _18916_/Q sky130_fd_sc_hd__dfxtp_1
X_14039_ _14611_/A vssd1 vssd1 vccd1 vccd1 _14039_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10181__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18847_ _19297_/CLK _18847_/D vssd1 vssd1 vccd1 vccd1 _18847_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09580_ _19736_/Q vssd1 vssd1 vccd1 vccd1 _09580_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18778_ _19071_/CLK _18778_/D vssd1 vssd1 vccd1 vccd1 _18778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_118_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17729_ _17597_/A _17721_/Y _17728_/X _17422_/A vssd1 vssd1 vccd1 vccd1 _17729_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_24_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10107__S1 _09714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__S0 _10660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12421__A2 _12482_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14262__S _14264_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10291__S0 _10260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09916_ _19323_/Q _18735_/Q _18772_/Q _18346_/Q _10114_/S _09888_/X vssd1 vssd1 vccd1
+ vccd1 _09916_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11145__C1 _09465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09880__A _10274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__S0 _09981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09847_ _18602_/Q _18873_/Q _19097_/Q _18841_/Q _09846_/X _09839_/A vssd1 vssd1 vccd1
+ vccd1 _09847_/X sky130_fd_sc_hd__mux4_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15093__S _15093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11915__A _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13606__S _13609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _10260_/A vssd1 vssd1 vccd1 vccd1 _10381_/S sky130_fd_sc_hd__buf_2
XFILLER_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__A1 _17696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _19332_/Q _11733_/X _11734_/X _11739_/X _11691_/X vssd1 vssd1 vccd1 vccd1
+ _11740_/X sky130_fd_sc_hd__o221a_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10030__S _10030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16926__A2 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _19853_/Q vssd1 vssd1 vccd1 vccd1 _18114_/A sky130_fd_sc_hd__buf_4
XFILLER_42_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14437__S _14439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13410_ _13398_/X _13408_/X _13409_/Y _13403_/X _18252_/Q vssd1 vssd1 vccd1 vccd1
+ _13410_/X sky130_fd_sc_hd__a32o_4
XFILLER_139_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10622_ _10689_/A _10622_/B vssd1 vssd1 vccd1 vccd1 _10622_/Y sky130_fd_sc_hd__nor2_1
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14390_ _14390_/A vssd1 vssd1 vccd1 vccd1 _18684_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12412__A2 _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12465__B _12465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ _19581_/Q _12638_/X _13340_/X _13265_/X vssd1 vssd1 vccd1 vccd1 _13341_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_155_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10423__B2 _19724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _10617_/A _10553_/B vssd1 vssd1 vccd1 vccd1 _10553_/X sky130_fd_sc_hd__or2_1
XANTENNA__10266__A _10518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16060_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16083_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_143_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13272_ _13051_/X _13255_/X _13258_/Y _13271_/X vssd1 vssd1 vccd1 vccd1 _15079_/A
+ sky130_fd_sc_hd__a22o_2
X_10484_ _18928_/Q _18694_/Q _19376_/Q _19024_/Q _10274_/A _10348_/A vssd1 vssd1 vccd1
+ vccd1 _10485_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17639__A0 _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15011_ _15011_/A vssd1 vssd1 vccd1 vccd1 _18947_/D sky130_fd_sc_hd__clkbuf_1
X_12223_ _12223_/A _12223_/B vssd1 vssd1 vccd1 vccd1 _12224_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14172__S _14180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10187__B1 _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12154_ _19347_/Q _11859_/X _12037_/X _12153_/Y _12102_/X vssd1 vssd1 vccd1 vccd1
+ _12154_/X sky130_fd_sc_hd__o221a_1
XFILLER_123_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11105_ _18387_/Q _18648_/Q _18547_/Q _18882_/Q _09624_/A _11020_/X vssd1 vssd1 vccd1
+ vccd1 _11105_/X sky130_fd_sc_hd__mux4_1
XFILLER_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19750_ _19779_/CLK _19750_/D vssd1 vssd1 vccd1 vccd1 _19750_/Q sky130_fd_sc_hd__dfxtp_1
X_16962_ _16932_/A _16956_/X _16961_/X _16954_/X vssd1 vssd1 vccd1 vccd1 _19638_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14900__S _14904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12085_ _19788_/Q _11445_/A _12143_/S vssd1 vssd1 vccd1 vccd1 _17215_/A sky130_fd_sc_hd__mux2_2
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18701_ _19256_/CLK _18701_/D vssd1 vssd1 vccd1 vccd1 _18701_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10034__S0 _09415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11036_ _18917_/Q _18683_/Q _19365_/Q _19013_/Q _11149_/A _09512_/A vssd1 vssd1 vccd1
+ vccd1 _11036_/X sky130_fd_sc_hd__mux4_1
X_15913_ _15913_/A vssd1 vssd1 vccd1 vccd1 _19291_/D sky130_fd_sc_hd__clkbuf_1
X_19681_ _19694_/CLK _19681_/D vssd1 vssd1 vccd1 vccd1 _19681_/Q sky130_fd_sc_hd__dfxtp_1
X_16893_ _19609_/Q _16889_/B _16892_/Y vssd1 vssd1 vccd1 vccd1 _19609_/D sky130_fd_sc_hd__o21a_1
XFILLER_103_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18632_ _19127_/CLK _18632_/D vssd1 vssd1 vccd1 vccd1 _18632_/Q sky130_fd_sc_hd__dfxtp_1
X_15844_ _13602_/X _19261_/Q _15848_/S vssd1 vssd1 vccd1 vccd1 _15845_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11544__B _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18563_ _19284_/CLK _18563_/D vssd1 vssd1 vccd1 vccd1 _18563_/Q sky130_fd_sc_hd__dfxtp_1
X_15775_ _15775_/A vssd1 vssd1 vccd1 vccd1 _19230_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _19147_/Q _12895_/X _12958_/A _19337_/Q _12986_/X vssd1 vssd1 vccd1 vccd1
+ _12987_/X sky130_fd_sc_hd__a221o_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _14534_/X _18820_/Q _14726_/S vssd1 vssd1 vccd1 vccd1 _14727_/A sky130_fd_sc_hd__mux2_1
X_17514_ _17653_/A _17514_/B vssd1 vssd1 vccd1 vccd1 _17514_/X sky130_fd_sc_hd__or2_1
X_11938_ _16967_/A _11939_/C _19642_/Q vssd1 vssd1 vccd1 vccd1 _11938_/Y sky130_fd_sc_hd__a21oi_1
X_18494_ _19085_/CLK _18494_/D vssd1 vssd1 vccd1 vccd1 _18494_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _17267_/X _17277_/X _17448_/S vssd1 vssd1 vccd1 vccd1 _17445_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10662__A1 _09597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14657_ _14537_/X _18789_/Q _14665_/S vssd1 vssd1 vccd1 vccd1 _14658_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18119__A1 _09351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11869_ _17630_/A _11950_/A _11949_/A vssd1 vssd1 vccd1 vccd1 _11870_/B sky130_fd_sc_hd__o21a_1
XFILLER_159_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15032__A _15099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ _15092_/A vssd1 vssd1 vccd1 vccd1 _13608_/X sky130_fd_sc_hd__clkbuf_2
X_17376_ _17396_/A vssd1 vssd1 vccd1 vccd1 _17511_/S sky130_fd_sc_hd__clkbuf_2
X_14588_ _14588_/A vssd1 vssd1 vccd1 vccd1 _18767_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13061__C1 _13060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16327_ _19425_/Q _16322_/C _16326_/Y vssd1 vssd1 vccd1 vccd1 _19425_/D sky130_fd_sc_hd__o21a_1
X_19115_ _19373_/CLK _19115_/D vssd1 vssd1 vccd1 vccd1 _19115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13539_ _18360_/Q _13538_/X _13545_/S vssd1 vssd1 vccd1 vccd1 _13540_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_158_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19046_ _19306_/CLK _19046_/D vssd1 vssd1 vccd1 vccd1 _19046_/Q sky130_fd_sc_hd__dfxtp_1
X_16258_ _16266_/A _16258_/B vssd1 vssd1 vccd1 vccd1 _16259_/A sky130_fd_sc_hd__or2_1
XFILLER_174_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15209_ _19023_/Q _15047_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15210_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15178__S _15184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12391__A _12391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16189_ _13541_/X _19368_/Q _16191_/S vssd1 vssd1 vccd1 vccd1 _16190_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09701_ _09868_/A vssd1 vssd1 vccd1 vccd1 _09840_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_101_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09632_ _09632_/A vssd1 vssd1 vccd1 vccd1 _10682_/A sky130_fd_sc_hd__buf_2
XFILLER_95_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10350__B1 _10297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _09563_/A vssd1 vssd1 vccd1 vccd1 _09820_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15641__S _15649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13950__A _14049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ _11219_/S vssd1 vssd1 vccd1 vccd1 _11151_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_130_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10785__S _10785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15592__A1 _12689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12285__B _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12158__A1 _19411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13397__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10814__A _10878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10264__S0 _10260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14720__S _14726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12910_ _12910_/A vssd1 vssd1 vccd1 vccd1 _18288_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13890_ _13922_/A vssd1 vssd1 vccd1 vccd1 _13903_/S sky130_fd_sc_hd__buf_4
XFILLER_101_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12841_ _19522_/Q _12939_/S _12953_/A _16529_/B _12840_/X vssd1 vssd1 vccd1 vccd1
+ _12841_/X sky130_fd_sc_hd__a221o_1
XFILLER_62_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _15559_/X _19155_/Q _15570_/S vssd1 vssd1 vccd1 vccd1 _15561_/A sky130_fd_sc_hd__mux2_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12772_ _18278_/Q _12766_/X _10080_/A _12769_/X vssd1 vssd1 vccd1 vccd1 _18278_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _13934_/X _18739_/Q _14511_/S vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__mux2_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _12447_/B _11722_/Y _11723_/S vssd1 vssd1 vccd1 vccd1 _11782_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10644__A1 _10074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14167__S _14169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15491_ _15489_/X _19143_/Q _15517_/S vssd1 vssd1 vccd1 vccd1 _15492_/A sky130_fd_sc_hd__mux2_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13071__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17230_/A vssd1 vssd1 vccd1 vccd1 _17410_/B sky130_fd_sc_hd__clkbuf_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ _14442_/A vssd1 vssd1 vccd1 vccd1 _18708_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15583__A1 _15582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11654_ _12184_/A vssd1 vssd1 vccd1 vccd1 _15488_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12397__A1 _12391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _09390_/A _10602_/X _10604_/X vssd1 vssd1 vccd1 vccd1 _10605_/X sky130_fd_sc_hd__a21o_1
X_17161_ _17161_/A vssd1 vssd1 vccd1 vccd1 _19705_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14373_ _15245_/B _16169_/B vssd1 vssd1 vccd1 vccd1 _14430_/A sky130_fd_sc_hd__nand2_2
XFILLER_11_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11585_ _18135_/A _18132_/A _11585_/C _11585_/D vssd1 vssd1 vccd1 vccd1 _11586_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18163__A _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16112_ _16111_/X _19349_/Q _16112_/S vssd1 vssd1 vccd1 vccd1 _16113_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13324_ _19548_/Q _12583_/X _13054_/X _19516_/Q _13323_/X vssd1 vssd1 vccd1 vccd1
+ _13324_/X sky130_fd_sc_hd__a221o_1
XFILLER_156_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17092_ _19692_/Q _15620_/X _17094_/S vssd1 vssd1 vccd1 vccd1 _17093_/A sky130_fd_sc_hd__mux2_1
X_10536_ _19281_/Q _19119_/Q _18528_/Q _18298_/Q _10481_/S _10262_/A vssd1 vssd1 vccd1
+ vccd1 _10536_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13346__B1 _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16043_ _16042_/X _19337_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16044_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13255_ input18/X _13134_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _13255_/X sky130_fd_sc_hd__a21o_1
X_10467_ _10250_/A _10464_/X _10466_/X _10243_/A vssd1 vssd1 vccd1 vccd1 _10467_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_109_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12206_ _11884_/X _12204_/Y _12256_/C _11835_/X vssd1 vssd1 vccd1 vccd1 _12206_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_124_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10255__S0 _10247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13186_ _19727_/Q _15572_/B _13360_/S vssd1 vssd1 vccd1 vccd1 _13186_/X sky130_fd_sc_hd__mux2_1
X_10398_ _19725_/Q vssd1 vssd1 vccd1 vccd1 _10398_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19802_ _19802_/CLK _19802_/D vssd1 vssd1 vccd1 vccd1 _19802_/Q sky130_fd_sc_hd__dfxtp_1
X_12137_ _18116_/A _12021_/X _12022_/X vssd1 vssd1 vccd1 vccd1 _12137_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11109__C1 _09553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17994_ _19770_/Q _19802_/Q _17994_/S vssd1 vssd1 vccd1 vccd1 _17995_/A sky130_fd_sc_hd__mux2_1
XFILLER_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19733_ _19736_/CLK _19733_/D vssd1 vssd1 vccd1 vccd1 _19733_/Q sky130_fd_sc_hd__dfxtp_4
X_16945_ _13410_/X _16943_/X _16944_/X _16933_/X vssd1 vssd1 vccd1 vccd1 _19632_/D
+ sky130_fd_sc_hd__o211a_1
X_12068_ _12068_/A vssd1 vssd1 vccd1 vccd1 _12274_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10558__S1 _09590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _11085_/A _11019_/B vssd1 vssd1 vccd1 vccd1 _11019_/Y sky130_fd_sc_hd__nor2_1
XFILLER_37_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19664_ _19667_/CLK _19664_/D vssd1 vssd1 vccd1 vccd1 _19664_/Q sky130_fd_sc_hd__dfxtp_1
X_16876_ _19603_/Q _16873_/B _16875_/Y vssd1 vssd1 vccd1 vccd1 _19603_/D sky130_fd_sc_hd__o21a_1
XFILLER_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17260__A1 _17722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18615_ _19367_/CLK _18615_/D vssd1 vssd1 vccd1 vccd1 _18615_/Q sky130_fd_sc_hd__dfxtp_1
X_15827_ _15827_/A vssd1 vssd1 vccd1 vccd1 _19253_/D sky130_fd_sc_hd__clkbuf_1
X_19595_ _19598_/CLK _19595_/D vssd1 vssd1 vccd1 vccd1 _19595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15461__S _15482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12085__A0 _19788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15758_ _15758_/A vssd1 vssd1 vccd1 vccd1 _19222_/D sky130_fd_sc_hd__clkbuf_1
X_18546_ _19298_/CLK _18546_/D vssd1 vssd1 vccd1 vccd1 _18546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10635__A1 _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14709_ _14614_/X _18813_/Q _14709_/S vssd1 vssd1 vccd1 vccd1 _14710_/A sky130_fd_sc_hd__mux2_1
X_15689_ _14592_/X _19192_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15690_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14077__S _14085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18477_ _19264_/CLK _18477_/D vssd1 vssd1 vccd1 vccd1 _18477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17428_ _11612_/X _17427_/X _12727_/X vssd1 vssd1 vccd1 vccd1 _17428_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_159_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17359_ _17359_/A vssd1 vssd1 vccd1 vccd1 _17359_/Y sky130_fd_sc_hd__inv_2
XFILLER_147_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09695__A _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19029_ _19502_/CLK _19029_/D vssd1 vssd1 vccd1 vccd1 _19029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10634__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17079__A1 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15636__S _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10020__C1 _10684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13945__A _18089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17251__A1 _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ _09606_/X _09609_/X _09611_/X _09613_/X _09614_/X vssd1 vssd1 vccd1 vccd1
+ _09615_/X sky130_fd_sc_hd__a221o_2
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09546_ _10680_/A vssd1 vssd1 vccd1 vccd1 _10014_/A sky130_fd_sc_hd__buf_2
XFILLER_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_0_0_clock_A clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ _09477_/A vssd1 vssd1 vccd1 vccd1 _09617_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_169_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_192_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19247_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11051__A1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13839__B _14197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ _11373_/A _11369_/X _09740_/X vssd1 vssd1 vccd1 vccd1 _11370_/X sky130_fd_sc_hd__o21a_1
XFILLER_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10321_ _10361_/A _10321_/B vssd1 vssd1 vccd1 vccd1 _10321_/X sky130_fd_sc_hd__or2_1
XFILLER_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ _13040_/A vssd1 vssd1 vccd1 vccd1 _18294_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10252_ _10323_/A _10251_/X _09728_/A vssd1 vssd1 vccd1 vccd1 _10252_/X sky130_fd_sc_hd__o21a_1
XFILLER_140_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10788__S1 _09506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ _18933_/Q _18699_/Q _19381_/Q _19029_/Q _09854_/X _09676_/A vssd1 vssd1 vccd1
+ vccd1 _10184_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14450__S _14456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_130_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19793_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18019__A0 _19781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input39_A io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14991_ _14991_/A vssd1 vssd1 vccd1 vccd1 _18941_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12303__A1 _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16730_ _16731_/B _16731_/C _19553_/Q vssd1 vssd1 vccd1 vccd1 _16732_/B sky130_fd_sc_hd__a21oi_1
XFILLER_115_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13942_ _13942_/A vssd1 vssd1 vccd1 vccd1 _18512_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16661_ _16806_/A vssd1 vssd1 vccd1 vccd1 _16696_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_145_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19299_/CLK sky130_fd_sc_hd__clkbuf_16
X_13873_ _14553_/A vssd1 vssd1 vccd1 vccd1 _13873_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15281__S _15289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18400_ _19314_/CLK _18400_/D vssd1 vssd1 vccd1 vccd1 _18400_/Q sky130_fd_sc_hd__dfxtp_1
X_15612_ _15629_/A vssd1 vssd1 vccd1 vccd1 _15612_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_90_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10960__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _09315_/B _13408_/B _13143_/S vssd1 vssd1 vccd1 vccd1 _12824_/X sky130_fd_sc_hd__mux2_1
X_16592_ _19511_/Q _16596_/C _16591_/Y vssd1 vssd1 vccd1 vccd1 _19511_/D sky130_fd_sc_hd__o21a_1
X_19380_ _19380_/CLK _19380_/D vssd1 vssd1 vccd1 vccd1 _19380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_131_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15543_ _19721_/Q _15542_/X _15543_/S vssd1 vssd1 vccd1 vccd1 _15543_/X sky130_fd_sc_hd__mux2_1
X_18331_ _19307_/CLK _18331_/D vssd1 vssd1 vccd1 vccd1 _18331_/Q sky130_fd_sc_hd__dfxtp_1
X_12755_ _12769_/A vssd1 vssd1 vccd1 vccd1 _12755_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11706_ _16947_/A _11706_/B _11706_/C vssd1 vssd1 vccd1 vccd1 _11706_/X sky130_fd_sc_hd__or3_1
XFILLER_15_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _19201_/CLK _18262_/D vssd1 vssd1 vccd1 vccd1 _18262_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13016__C1 _13015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15556__A1 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15474_ _15474_/A vssd1 vssd1 vccd1 vccd1 _16024_/S sky130_fd_sc_hd__buf_2
X_12686_ _19611_/Q _12501_/X _12503_/X _19479_/Q _12685_/X vssd1 vssd1 vccd1 vccd1
+ _12687_/B sky130_fd_sc_hd__a221o_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14425_ _14425_/A vssd1 vssd1 vccd1 vccd1 _18700_/D sky130_fd_sc_hd__clkbuf_1
X_17213_ _17743_/B _12089_/A _17261_/S vssd1 vssd1 vccd1 vccd1 _17213_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18193_ _18234_/A vssd1 vssd1 vccd1 vccd1 _18193_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11637_ _11608_/B _17317_/A _11606_/X vssd1 vssd1 vccd1 vccd1 _11638_/B sky130_fd_sc_hd__a21oi_4
XFILLER_129_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17144_ _17163_/A vssd1 vssd1 vccd1 vccd1 _17160_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__10476__S0 _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14356_ _14356_/A vssd1 vssd1 vccd1 vccd1 _14365_/S sky130_fd_sc_hd__buf_4
X_11568_ _11565_/A _11513_/A _09327_/A _11559_/A vssd1 vssd1 vccd1 vccd1 _11672_/S
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13307_ _13360_/S _10077_/Y _12942_/S _13306_/Y vssd1 vssd1 vccd1 vccd1 _13307_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_157_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17075_ _19684_/Q _15574_/X _17083_/S vssd1 vssd1 vccd1 vccd1 _17076_/A sky130_fd_sc_hd__mux2_1
X_10519_ _10519_/A vssd1 vssd1 vccd1 vccd1 _10519_/Y sky130_fd_sc_hd__inv_2
XFILLER_155_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14287_ _14290_/A _18220_/B vssd1 vssd1 vccd1 vccd1 _14288_/A sky130_fd_sc_hd__and2_2
X_11499_ _12861_/A vssd1 vssd1 vccd1 vccd1 _11499_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_170_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16026_ _16026_/A vssd1 vssd1 vccd1 vccd1 _19334_/D sky130_fd_sc_hd__clkbuf_1
X_13238_ _13234_/X _13236_/Y _13237_/Y vssd1 vssd1 vccd1 vccd1 _15073_/A sky130_fd_sc_hd__a21oi_4
XFILLER_170_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17237__A _17237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _13153_/X _13165_/Y _13168_/Y vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__a21oi_4
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17977_ _16126_/A _19794_/Q _17979_/S vssd1 vssd1 vccd1 vccd1 _17978_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19716_ _19720_/CLK _19716_/D vssd1 vssd1 vccd1 vccd1 _19716_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_66_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16928_ _19627_/Q _12674_/X _16927_/X _16269_/X vssd1 vssd1 vccd1 vccd1 _19627_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_38_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17233__A1 _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19647_ _19695_/CLK _19647_/D vssd1 vssd1 vccd1 vccd1 _19647_/Q sky130_fd_sc_hd__dfxtp_1
X_16859_ _19597_/Q _16856_/B _16858_/Y vssd1 vssd1 vccd1 vccd1 _19597_/D sky130_fd_sc_hd__o21a_1
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09400_ _18510_/Q _19005_/Q _10602_/S vssd1 vssd1 vccd1 vccd1 _09400_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19578_ _19581_/CLK _19578_/D vssd1 vssd1 vccd1 vccd1 _19578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09331_ _09331_/A vssd1 vssd1 vccd1 vccd1 _18122_/A sky130_fd_sc_hd__buf_2
X_18529_ _19120_/CLK _18529_/D vssd1 vssd1 vccd1 vccd1 _18529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _19832_/Q _19831_/Q _19834_/Q _19833_/Q vssd1 vssd1 vccd1 vccd1 _12508_/C
+ sky130_fd_sc_hd__or4bb_4
XFILLER_139_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16744__B1 _16718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14535__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ _14297_/B _11522_/A vssd1 vssd1 vccd1 vccd1 _09193_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15366__S _15372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12533__B2 _19344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14286__A1 input48/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_62_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19502_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__14286__B2 _18125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11195__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10942__S1 _11174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_166_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ _18919_/Q _18685_/Q _19367_/Q _19015_/Q _10873_/S _11174_/A vssd1 vssd1 vccd1
+ vccd1 _10871_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_77_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19731_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_72_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09529_ _18643_/Q vssd1 vssd1 vccd1 vccd1 _10920_/A sky130_fd_sc_hd__inv_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10539__A _19722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12540_ _19440_/Q _12515_/X _12539_/X vssd1 vssd1 vccd1 vccd1 _12540_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11272__A1 _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12471_ _12474_/A _12471_/B vssd1 vssd1 vccd1 vccd1 _12471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14210_ _14210_/A vssd1 vssd1 vccd1 vccd1 _18613_/D sky130_fd_sc_hd__clkbuf_1
X_11422_ _11422_/A vssd1 vssd1 vccd1 vccd1 _11433_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_15190_ _15190_/A vssd1 vssd1 vccd1 vccd1 _19014_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_165_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12473__B _12473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14141_ _18583_/Q _13969_/X _14147_/S vssd1 vssd1 vccd1 vccd1 _14142_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11353_ _11443_/A _11446_/A _11443_/C _10402_/A _11352_/Y vssd1 vssd1 vccd1 vccd1
+ _11439_/C sky130_fd_sc_hd__a311o_1
XANTENNA__10274__A _10274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19324_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_152_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10304_ _10304_/A _10304_/B vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__or2_1
XFILLER_141_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14072_ _13867_/X _18553_/Q _14074_/S vssd1 vssd1 vccd1 vccd1 _14073_/A sky130_fd_sc_hd__mux2_1
X_11284_ _11284_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _11284_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15276__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17900_ _17490_/X _17897_/Y _17899_/Y vssd1 vssd1 vccd1 vccd1 _17900_/Y sky130_fd_sc_hd__a21oi_1
X_13023_ _11538_/X _13021_/X _13022_/X vssd1 vssd1 vccd1 vccd1 _15031_/A sky130_fd_sc_hd__o21a_4
XANTENNA__14180__S _14180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10235_ _09713_/A _10232_/X _10234_/X vssd1 vssd1 vccd1 vccd1 _10235_/X sky130_fd_sc_hd__a21o_1
X_18880_ _19268_/CLK _18880_/D vssd1 vssd1 vccd1 vccd1 _18880_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_105_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17831_ _17831_/A vssd1 vssd1 vccd1 vccd1 _17831_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10166_ _18503_/Q _18998_/Q _10166_/S vssd1 vssd1 vccd1 vccd1 _10167_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output145_A _11975_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10550__A3 _18830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17762_ _12060_/A _17737_/X _17760_/X _17761_/X vssd1 vssd1 vccd1 vccd1 _17762_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14974_ _18933_/Q vssd1 vssd1 vccd1 vccd1 _14975_/A sky130_fd_sc_hd__clkbuf_1
X_10097_ _18600_/Q _18871_/Q _19095_/Q _18839_/Q _10093_/S _09715_/A vssd1 vssd1 vccd1
+ vccd1 _10097_/X sky130_fd_sc_hd__mux4_1
XFILLER_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19501_ _19502_/CLK _19501_/D vssd1 vssd1 vccd1 vccd1 _19501_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10299__C1 _09831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16713_ _16737_/A _16713_/B _16722_/D vssd1 vssd1 vccd1 vccd1 _19547_/D sky130_fd_sc_hd__nor3_1
XFILLER_48_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13925_ _14605_/A vssd1 vssd1 vccd1 vccd1 _13925_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17693_ _17696_/A _17696_/B _17896_/S vssd1 vssd1 vccd1 vccd1 _17693_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17766__A2 _17215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19432_ _19436_/CLK _19432_/D vssd1 vssd1 vccd1 vccd1 _19432_/Q sky130_fd_sc_hd__dfxtp_1
X_16644_ _16666_/A _16644_/B vssd1 vssd1 vccd1 vccd1 _16644_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13856_ _13856_/A vssd1 vssd1 vccd1 vccd1 _18485_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12807_ _14642_/C _14998_/A vssd1 vssd1 vccd1 vccd1 _15173_/A sky130_fd_sc_hd__nand2_1
X_19363_ _19364_/CLK _19363_/D vssd1 vssd1 vccd1 vccd1 _19363_/Q sky130_fd_sc_hd__dfxtp_1
X_16575_ _19506_/Q _19505_/Q _16575_/C vssd1 vssd1 vccd1 vccd1 _16578_/B sky130_fd_sc_hd__and3_1
X_13787_ _12999_/X _18458_/Q _13787_/S vssd1 vssd1 vccd1 vccd1 _13788_/A sky130_fd_sc_hd__mux2_1
XFILLER_163_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10999_ _11195_/A _10999_/B vssd1 vssd1 vccd1 vccd1 _10999_/X sky130_fd_sc_hd__or2_1
XFILLER_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18314_ _19071_/CLK _18314_/D vssd1 vssd1 vccd1 vccd1 _18314_/Q sky130_fd_sc_hd__dfxtp_1
X_15526_ _15524_/X _19148_/Q _15544_/S vssd1 vssd1 vccd1 vccd1 _15527_/A sky130_fd_sc_hd__mux2_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _17795_/A vssd1 vssd1 vccd1 vccd1 _12744_/A sky130_fd_sc_hd__buf_2
XFILLER_124_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19294_ _19326_/CLK _19294_/D vssd1 vssd1 vccd1 vccd1 _19294_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18245_ _18248_/A _18245_/B vssd1 vssd1 vccd1 vccd1 _18246_/A sky130_fd_sc_hd__and2_1
X_15457_ _19134_/Q _15095_/X _15459_/S vssd1 vssd1 vccd1 vccd1 _15458_/A sky130_fd_sc_hd__mux2_1
X_12669_ _12557_/X _12667_/X _12668_/Y _12549_/X _18263_/Q vssd1 vssd1 vccd1 vccd1
+ _12669_/X sky130_fd_sc_hd__a32o_4
XFILLER_31_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14408_ _14430_/A vssd1 vssd1 vccd1 vccd1 _14417_/S sky130_fd_sc_hd__buf_4
X_18176_ _18190_/A _18176_/B vssd1 vssd1 vccd1 vccd1 _18177_/A sky130_fd_sc_hd__and2_1
X_15388_ _15388_/A vssd1 vssd1 vccd1 vccd1 _19103_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11110__S1 _11020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14339_ _13896_/X _18663_/Q _14343_/S vssd1 vssd1 vccd1 vccd1 _14340_/A sky130_fd_sc_hd__mux2_1
X_17127_ _17127_/A _17127_/B vssd1 vssd1 vccd1 vccd1 _17127_/Y sky130_fd_sc_hd__nor2_1
XFILLER_171_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10184__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ _17058_/A vssd1 vssd1 vccd1 vccd1 _19676_/D sky130_fd_sc_hd__clkbuf_1
X_16009_ _16008_/X _19331_/Q _16025_/S vssd1 vssd1 vccd1 vccd1 _16010_/A sky130_fd_sc_hd__mux2_1
X_09880_ _10274_/A vssd1 vssd1 vccd1 vccd1 _10341_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__14090__S _14096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10621__S0 _10566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11727__B _17252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11219__S _11219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15914__S _15920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12818__A2 _12817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17206__A1 _12195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09314_ _11699_/A _11700_/B _11702_/D vssd1 vssd1 vccd1 vccd1 _11743_/C sky130_fd_sc_hd__a21o_2
XFILLER_40_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17430__A _17831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10688__S0 _10566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12451__B1 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09245_ _09274_/C vssd1 vssd1 vccd1 vccd1 _16622_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09176_ _09176_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _17108_/B sky130_fd_sc_hd__nand2_2
XFILLER_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12754__A1 hold13/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09883__A _09955_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17693__A1 _17696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_92_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15096__S _15099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11918__A _18146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13609__S _13609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10020_ _09768_/A _10016_/Y _10018_/Y _10684_/A vssd1 vssd1 vccd1 vccd1 _10020_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_88_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11190__B1 _10883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__B _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15824__S _15826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17605__A _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11971_ _12011_/C _12372_/A _11970_/X vssd1 vssd1 vccd1 vccd1 _11971_/X sky130_fd_sc_hd__or3b_1
XANTENNA__17748__A2 _17741_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13710_ _12945_/X _18424_/Q _13714_/S vssd1 vssd1 vccd1 vccd1 _13711_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12690__A0 _12689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ _11116_/A vssd1 vssd1 vccd1 vccd1 _10981_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15125__A _15171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14690_ _14585_/X _18804_/Q _14698_/S vssd1 vssd1 vccd1 vccd1 _14691_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12468__B _12468_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _13641_/A vssd1 vssd1 vccd1 vccd1 _18393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ _10853_/A vssd1 vssd1 vccd1 vccd1 _10853_/Y sky130_fd_sc_hd__inv_2
XFILLER_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16360_ _19435_/Q _16363_/C _16359_/X vssd1 vssd1 vccd1 vccd1 _16360_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11245__A1 _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13572_ _13572_/A vssd1 vssd1 vccd1 vccd1 _18370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10679__S0 _10055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ _10784_/A vssd1 vssd1 vccd1 vccd1 _10784_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11193__A1_N _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _14614_/X _19069_/Q _15311_/S vssd1 vssd1 vccd1 vccd1 _15312_/A sky130_fd_sc_hd__mux2_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _13391_/B vssd1 vssd1 vccd1 vccd1 _12955_/B sky130_fd_sc_hd__inv_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16291_ _16291_/A vssd1 vssd1 vccd1 vccd1 _19413_/D sky130_fd_sc_hd__clkbuf_1
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15242_ _15242_/A vssd1 vssd1 vccd1 vccd1 _19038_/D sky130_fd_sc_hd__clkbuf_1
X_18030_ _19786_/Q _12066_/A _18038_/S vssd1 vssd1 vccd1 vccd1 _18031_/A sky130_fd_sc_hd__mux2_1
X_12454_ _12454_/A _12461_/B vssd1 vssd1 vccd1 vccd1 _12454_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12745__A1 hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11405_ _19329_/Q _18741_/Q _18778_/Q _18352_/Q _09815_/X _09788_/A vssd1 vssd1 vccd1
+ vccd1 _11405_/X sky130_fd_sc_hd__mux4_1
X_15173_ _15173_/A _15173_/B vssd1 vssd1 vccd1 vccd1 _15230_/A sky130_fd_sc_hd__nor2_2
XANTENNA__15795__A _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12385_ _12385_/A _17899_/B vssd1 vssd1 vccd1 vccd1 _12386_/A sky130_fd_sc_hd__nor2_1
XFILLER_165_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14124_ _18096_/A _14860_/B _14715_/C _14642_/C vssd1 vssd1 vccd1 vccd1 _15317_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11336_ _19279_/Q _19117_/Q _18526_/Q _18296_/Q _10633_/S _10060_/A vssd1 vssd1 vccd1
+ vccd1 _11336_/X sky130_fd_sc_hd__mux4_1
XFILLER_125_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18932_ _19380_/CLK _18932_/D vssd1 vssd1 vccd1 vccd1 _18932_/Q sky130_fd_sc_hd__dfxtp_1
X_14055_ _13837_/X _18545_/Q _14063_/S vssd1 vssd1 vccd1 vccd1 _14056_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11267_ _11033_/X _11264_/Y _11266_/Y _11232_/A vssd1 vssd1 vccd1 vccd1 _11267_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13006_ _13055_/A vssd1 vssd1 vccd1 vccd1 _13006_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10218_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10218_/Y sky130_fd_sc_hd__nand2_1
X_18863_ _19119_/CLK _18863_/D vssd1 vssd1 vccd1 vccd1 _18863_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11198_ _11242_/A _11197_/X _11257_/A vssd1 vssd1 vccd1 vccd1 _11198_/X sky130_fd_sc_hd__a21o_1
X_17814_ _17659_/X _17811_/X _17813_/X vssd1 vssd1 vccd1 vccd1 _17814_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_121_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10149_ _19320_/Q _18732_/Q _18769_/Q _18343_/Q _09846_/X _09871_/X vssd1 vssd1 vccd1
+ vccd1 _10150_/B sky130_fd_sc_hd__mux4_1
XFILLER_95_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18794_ _19180_/CLK _18794_/D vssd1 vssd1 vccd1 vccd1 _18794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11159__S1 _11033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17745_ _17812_/A _17745_/B vssd1 vssd1 vccd1 vccd1 _17745_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14957_ _14957_/A vssd1 vssd1 vccd1 vccd1 _18924_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12659__A _13008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15035__A _15035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ _13908_/A vssd1 vssd1 vccd1 vccd1 _18501_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17676_ _17680_/A _17680_/B vssd1 vssd1 vccd1 vccd1 _17676_/Y sky130_fd_sc_hd__nand2_1
X_14888_ _14888_/A vssd1 vssd1 vccd1 vccd1 _18891_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19415_ _19699_/CLK _19415_/D vssd1 vssd1 vccd1 vccd1 _19415_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_74_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ _16659_/A vssd1 vssd1 vccd1 vccd1 _16634_/B sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13839_ _19814_/Q _14197_/B _15854_/A vssd1 vssd1 vccd1 vccd1 _16622_/B sky130_fd_sc_hd__or3_4
XANTENNA__17250__A _17250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09968__A _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19346_ _19349_/CLK _19346_/D vssd1 vssd1 vccd1 vccd1 _19346_/Q sky130_fd_sc_hd__dfxtp_2
X_16558_ hold3/X _16559_/C _19500_/Q vssd1 vssd1 vccd1 vccd1 _16560_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10444__C1 _09812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__A1 input32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15509_ _15478_/X _15505_/X _15507_/Y _15508_/X hold12/X vssd1 vssd1 vccd1 vccd1
+ _15509_/X sky130_fd_sc_hd__a32o_4
XANTENNA__14085__S _14085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19277_ _19310_/CLK _19277_/D vssd1 vssd1 vccd1 vccd1 _19277_/Q sky130_fd_sc_hd__dfxtp_1
X_16489_ _16546_/A vssd1 vssd1 vccd1 vccd1 _16489_/X sky130_fd_sc_hd__buf_2
X_18228_ _18228_/A vssd1 vssd1 vccd1 vccd1 _19860_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15909__S _15909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18159_ input59/X _18155_/X _18066_/S _12657_/X _18077_/A vssd1 vssd1 vccd1 vccd1
+ _18160_/B sky130_fd_sc_hd__a32o_1
XFILLER_11_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18081__A _18081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14813__S _14821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _09690_/A _09931_/X _10195_/A vssd1 vssd1 vccd1 vccd1 _09932_/X sky130_fd_sc_hd__a21o_1
XFILLER_104_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09863_ _10148_/A _09863_/B vssd1 vssd1 vccd1 vccd1 _09863_/X sky130_fd_sc_hd__or2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09460__S0 _09441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11711__A2 _11710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _10214_/A vssd1 vssd1 vccd1 vccd1 _09964_/A sky130_fd_sc_hd__buf_2
XFILLER_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10070__S1 _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_39_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10817__A _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ _19859_/Q _13619_/A _09225_/Y _09226_/X _09227_/Y vssd1 vssd1 vccd1 vccd1
+ _09230_/B sky130_fd_sc_hd__o221a_2
XFILLER_167_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11086__S0 _10969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09159_ _09186_/A _09186_/B _09176_/B vssd1 vssd1 vccd1 vccd1 _17165_/A sky130_fd_sc_hd__or3b_2
XFILLER_107_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12170_ _12170_/A _17222_/A vssd1 vssd1 vccd1 vccd1 _12170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17319__B _17319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11648__A _19394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ _09476_/A _11109_/X _11119_/X _09576_/A _11120_/Y vssd1 vssd1 vccd1 vccd1
+ _12444_/B sky130_fd_sc_hd__o32a_4
XFILLER_150_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11052_ _09416_/A _11049_/X _11051_/X vssd1 vssd1 vccd1 vccd1 _11052_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09118__A _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _19196_/Q _18810_/Q _19260_/Q _18379_/Q _09776_/A _09547_/X vssd1 vssd1 vccd1
+ vccd1 _10004_/B sky130_fd_sc_hd__mux4_1
XFILLER_88_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15860_ _15860_/A vssd1 vssd1 vccd1 vccd1 _19267_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10061__S1 _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14101__A0 _13909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input21_A io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ _14811_/A vssd1 vssd1 vccd1 vccd1 _18857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_92_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15791_ _13525_/X _19237_/Q _15793_/S vssd1 vssd1 vccd1 vccd1 _15792_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09659__A1 _09640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17530_ _17530_/A vssd1 vssd1 vccd1 vccd1 _17672_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14742_ _14557_/X _18827_/Q _14748_/S vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11954_ _11955_/A _17221_/A vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11466__B2 _12442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905_ _11020_/A vssd1 vssd1 vccd1 vccd1 _11220_/A sky130_fd_sc_hd__buf_2
XANTENNA__10674__C1 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17461_ _17461_/A _17463_/B vssd1 vssd1 vccd1 vccd1 _17468_/B sky130_fd_sc_hd__nand2_1
X_14673_ _14673_/A vssd1 vssd1 vccd1 vccd1 _18796_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17325__C_N _17190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11885_ _16963_/A _11886_/C _19640_/Q vssd1 vssd1 vccd1 vccd1 _11885_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_output108_A _17175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19200_ _19264_/CLK _19200_/D vssd1 vssd1 vccd1 vccd1 _19200_/Q sky130_fd_sc_hd__dfxtp_1
X_16412_ _16427_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _16412_/Y sky130_fd_sc_hd__nor2_1
X_13624_ _13624_/A vssd1 vssd1 vccd1 vccd1 _18385_/D sky130_fd_sc_hd__clkbuf_1
X_10836_ _11075_/A vssd1 vssd1 vccd1 vccd1 _10837_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17392_ _17739_/S vssd1 vssd1 vccd1 vccd1 _17392_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19131_ _19325_/CLK _19131_/D vssd1 vssd1 vccd1 vccd1 _19131_/Q sky130_fd_sc_hd__dfxtp_1
X_16343_ _16355_/D vssd1 vssd1 vccd1 vccd1 _16351_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13555_ _18365_/Q _13554_/X _13561_/S vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10767_ _18586_/Q _18857_/Q _19081_/Q _18825_/Q _10030_/S _09707_/A vssd1 vssd1 vccd1
+ vccd1 _10767_/X sky130_fd_sc_hd__mux4_1
XFILLER_160_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ _12782_/A vssd1 vssd1 vccd1 vccd1 _13004_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_146_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16274_ _18150_/A _16274_/B vssd1 vssd1 vccd1 vccd1 _16275_/A sky130_fd_sc_hd__or2_1
X_19062_ _19471_/CLK _19062_/D vssd1 vssd1 vccd1 vccd1 _19062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ _13209_/X _18342_/Q _13492_/S vssd1 vssd1 vccd1 vccd1 _13487_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _10585_/A _10695_/X _10697_/X vssd1 vssd1 vccd1 vccd1 _10698_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12718__A1 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12718__B2 _12694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15225_ _15225_/A vssd1 vssd1 vccd1 vccd1 _19030_/D sky130_fd_sc_hd__clkbuf_1
X_18013_ _18013_/A vssd1 vssd1 vccd1 vccd1 _19778_/D sky130_fd_sc_hd__clkbuf_1
X_12437_ _11686_/X _12433_/Y _12435_/Y _12436_/X vssd1 vssd1 vccd1 vccd1 _12437_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_154_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14860__C _18091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15156_ _19000_/Q _15076_/X _15156_/S vssd1 vssd1 vccd1 vccd1 _15157_/A sky130_fd_sc_hd__mux2_1
X_12368_ _19659_/Q _12394_/C vssd1 vssd1 vccd1 vccd1 _12368_/X sky130_fd_sc_hd__and2_1
X_14107_ _13918_/X _18569_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _14108_/A sky130_fd_sc_hd__mux2_1
X_11319_ _11319_/A vssd1 vssd1 vccd1 vccd1 _11319_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11558__A _17174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15087_ _18971_/Q _15086_/X _15093_/S vssd1 vssd1 vccd1 vccd1 _15088_/A sky130_fd_sc_hd__mux2_1
X_12299_ _11884_/X _12297_/Y _12343_/C _11962_/A vssd1 vssd1 vccd1 vccd1 _12299_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_113_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13143__A1 _12590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18915_ _19074_/CLK _18915_/D vssd1 vssd1 vccd1 vccd1 _18915_/Q sky130_fd_sc_hd__dfxtp_1
X_14038_ _14038_/A vssd1 vssd1 vccd1 vccd1 _18540_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10181__B _12471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17245__A _17245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18846_ _19328_/CLK _18846_/D vssd1 vssd1 vccd1 vccd1 _18846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16093__B1 _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18777_ _19328_/CLK _18777_/D vssd1 vssd1 vccd1 vccd1 _18777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15989_ _15989_/A vssd1 vssd1 vccd1 vccd1 _19325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17728_ _17537_/X _17725_/Y _17727_/X vssd1 vssd1 vccd1 vccd1 _17728_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17659_ _17659_/A vssd1 vssd1 vccd1 vccd1 _17659_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12957__A1 _19146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19329_ _19329_/CLK _19329_/D vssd1 vssd1 vccd1 vccd1 _19329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10637__A _10689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13382__B2 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10291__S1 _10263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09915_ _10209_/A vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__buf_2
XFILLER_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09846_ _10186_/S vssd1 vssd1 vccd1 vccd1 _09846_/X sky130_fd_sc_hd__clkbuf_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11240__S0 _11173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__S1 _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _10520_/S vssd1 vssd1 vccd1 vccd1 _10260_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14634__A1 input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16994__A _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14634__B2 _18114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14718__S _14726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11670_ _11670_/A vssd1 vssd1 vccd1 vccd1 _11890_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10621_ _19182_/Q _18796_/Q _19246_/Q _18365_/Q _10566_/X _10586_/X vssd1 vssd1 vccd1
+ vccd1 _10622_/B sky130_fd_sc_hd__mux4_1
XFILLER_23_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13340_ _19167_/Q _12784_/X _12532_/X _19357_/Q _13339_/X vssd1 vssd1 vccd1 vccd1
+ _13340_/X sky130_fd_sc_hd__a221o_2
XANTENNA__10423__A2 _10411_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17887__A1 _11512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10552_ _18399_/Q _18660_/Q _18559_/Q _18894_/Q _10542_/A _09443_/A vssd1 vssd1 vccd1
+ vccd1 _10553_/B sky130_fd_sc_hd__mux4_1
XFILLER_127_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13858__A _13941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13271_ _12848_/A _13270_/X _12831_/X vssd1 vssd1 vccd1 vccd1 _13271_/X sky130_fd_sc_hd__o21a_1
X_10483_ _10482_/A _10480_/Y _10482_/Y _10531_/A vssd1 vssd1 vccd1 vccd1 _10483_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12762__A _12769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15010_ _18947_/Q _15009_/X _15013_/S vssd1 vssd1 vccd1 vccd1 _15011_/A sky130_fd_sc_hd__mux2_1
XFILLER_136_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12222_ _12173_/A _12173_/B _12196_/A _12195_/A _12168_/A vssd1 vssd1 vccd1 vccd1
+ _12223_/B sky130_fd_sc_hd__a221o_1
XANTENNA_input69_A io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10187__A1 _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _11858_/S _12150_/Y _12226_/C _12152_/X vssd1 vssd1 vccd1 vccd1 _12153_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11104_ _11278_/A _11104_/B vssd1 vssd1 vccd1 vccd1 _11104_/Y sky130_fd_sc_hd__nor2_1
X_16961_ _19638_/Q _16971_/B vssd1 vssd1 vccd1 vccd1 _16961_/X sky130_fd_sc_hd__or2_1
X_12084_ _17768_/B _12084_/B vssd1 vssd1 vccd1 vccd1 _12087_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14689__A _14700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18700_ _19320_/CLK _18700_/D vssd1 vssd1 vccd1 vccd1 _18700_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11035_ _11033_/X _11034_/X _09531_/A vssd1 vssd1 vccd1 vccd1 _11035_/X sky130_fd_sc_hd__a21o_1
X_15912_ _19291_/Q _14601_/A _15920_/S vssd1 vssd1 vccd1 vccd1 _15913_/A sky130_fd_sc_hd__mux2_1
X_19680_ _19688_/CLK _19680_/D vssd1 vssd1 vccd1 vccd1 _19680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11231__S0 _11265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10034__S1 _09443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16892_ _16915_/A _16896_/C vssd1 vssd1 vccd1 vccd1 _16892_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12884__B1 _12883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18631_ _18902_/CLK _18631_/D vssd1 vssd1 vccd1 vccd1 _18631_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15843_ _15843_/A vssd1 vssd1 vccd1 vccd1 _19260_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18562_ _19377_/CLK _18562_/D vssd1 vssd1 vccd1 vccd1 _18562_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12986_ _19673_/Q _12817_/X _12680_/A _19640_/Q vssd1 vssd1 vccd1 vccd1 _12986_/X
+ sky130_fd_sc_hd__a22o_1
X_15774_ _13605_/X _19230_/Q _15776_/S vssd1 vssd1 vccd1 vccd1 _15775_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17513_ _17615_/B _17512_/X _17524_/S vssd1 vssd1 vccd1 vccd1 _17514_/B sky130_fd_sc_hd__mux2_1
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _14725_/A vssd1 vssd1 vccd1 vccd1 _18819_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11937_ _12654_/B vssd1 vssd1 vccd1 vccd1 _12230_/A sky130_fd_sc_hd__buf_2
XANTENNA__10111__A1 _09667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18493_ _19374_/CLK _18493_/D vssd1 vssd1 vccd1 vccd1 _18493_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10111__B2 _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11841__A _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17444_/A vssd1 vssd1 vccd1 vccd1 _17444_/Y sky130_fd_sc_hd__clkinv_2
X_14656_ _14713_/S vssd1 vssd1 vccd1 vccd1 _14665_/S sky130_fd_sc_hd__buf_2
X_11868_ _12208_/A _12454_/A _11890_/C _19864_/Q vssd1 vssd1 vccd1 vccd1 _17642_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18119__A2 _18091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10819_ _11184_/A _10819_/B vssd1 vssd1 vccd1 vccd1 _10819_/X sky130_fd_sc_hd__or2_1
XFILLER_32_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13607_ _13607_/A vssd1 vssd1 vccd1 vccd1 _18381_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11560__B _11560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17375_ _17293_/X _17289_/X _17375_/S vssd1 vssd1 vccd1 vccd1 _17375_/X sky130_fd_sc_hd__mux2_1
X_14587_ _14585_/X _18767_/Q _14599_/S vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__mux2_1
X_11799_ _11794_/X _11797_/X _11798_/Y vssd1 vssd1 vccd1 vccd1 _11799_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19114_ _19370_/CLK _19114_/D vssd1 vssd1 vccd1 vccd1 _19114_/Q sky130_fd_sc_hd__dfxtp_1
X_16326_ _16344_/A _16331_/C vssd1 vssd1 vccd1 vccd1 _16326_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ _15022_/A vssd1 vssd1 vccd1 vccd1 _13538_/X sky130_fd_sc_hd__buf_2
XFILLER_158_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19045_ _19239_/CLK _19045_/D vssd1 vssd1 vccd1 vccd1 _19045_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15459__S _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16257_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16266_/A sky130_fd_sc_hd__clkbuf_1
X_13469_ _13469_/A vssd1 vssd1 vccd1 vccd1 _18334_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14363__S _14365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15217_/S sky130_fd_sc_hd__buf_4
X_16188_ _16188_/A vssd1 vssd1 vccd1 vccd1 _19367_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11288__A _11288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15983__A _15983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ _18992_/Q _15051_/X _15145_/S vssd1 vssd1 vccd1 vccd1 _15140_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13116__A1 _13132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09700_ _09700_/A vssd1 vssd1 vccd1 vccd1 _09868_/A sky130_fd_sc_hd__buf_2
XFILLER_101_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18055__A1 _12321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11222__S0 _11074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__B1 _12521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16066__A0 _15536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09631_ _11335_/A _09629_/X _09630_/X vssd1 vssd1 vccd1 vccd1 _09631_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18829_ _19245_/CLK _18829_/D vssd1 vssd1 vccd1 vccd1 _18829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10350__A1 _10394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15922__S _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13008__A _13008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _09630_/A vssd1 vssd1 vccd1 vccd1 _09563_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ _18641_/Q vssd1 vssd1 vccd1 vccd1 _11219_/S sky130_fd_sc_hd__buf_2
XFILLER_64_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_0_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13442__S _13448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09221__A _11618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13355__B2 _19358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09654__S0 _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10264__S1 _10263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14304__A0 _13845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11118__B1 _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18046__A1 _19414_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12330__A2 _12477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09829_ _09829_/A vssd1 vssd1 vccd1 vccd1 _09830_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15804__A0 _13544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _16331_/B _13005_/A _12839_/X vssd1 vssd1 vccd1 vccd1 _12840_/X sky130_fd_sc_hd__o21a_1
XFILLER_74_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _18277_/Q _12766_/X _10082_/A _12769_/X vssd1 vssd1 vccd1 vccd1 _18277_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14448__S _14456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _12159_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _11722_/Y sky130_fd_sc_hd__nand2_2
X_14510_ _14510_/A vssd1 vssd1 vccd1 vccd1 _18738_/D sky130_fd_sc_hd__clkbuf_1
X_15490_ _15636_/S vssd1 vssd1 vccd1 vccd1 _15517_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__B _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11653_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11653_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14441_ _13937_/X _18708_/Q _14443_/S vssd1 vssd1 vccd1 vccd1 _14442_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10604_ _09688_/A _10603_/X _09982_/A vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__a21o_1
XFILLER_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14372_ _14372_/A _15173_/B vssd1 vssd1 vccd1 vccd1 _16169_/B sky130_fd_sc_hd__nor2_1
X_17160_ _17160_/A _17160_/B vssd1 vssd1 vccd1 vccd1 _17161_/A sky130_fd_sc_hd__and2_1
XFILLER_128_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11584_ _18138_/A _11584_/B _19865_/Q vssd1 vssd1 vccd1 vccd1 _11585_/D sky130_fd_sc_hd__or3b_1
XFILLER_167_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13323_ _19452_/Q _12962_/X _13322_/X vssd1 vssd1 vccd1 vccd1 _13323_/X sky130_fd_sc_hd__o21a_1
X_16111_ _12233_/X _15582_/X _16110_/Y vssd1 vssd1 vccd1 vccd1 _16111_/X sky130_fd_sc_hd__a21o_1
X_10535_ _10535_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10535_/Y sky130_fd_sc_hd__nor2_1
X_17091_ _17091_/A vssd1 vssd1 vccd1 vccd1 _19691_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14183__S _14191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16042_ _15515_/X _16041_/Y _16052_/S vssd1 vssd1 vccd1 vccd1 _16042_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13254_ _13254_/A vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_124_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10466_ _10509_/A _10466_/B vssd1 vssd1 vccd1 vccd1 _10466_/X sky130_fd_sc_hd__or2_1
XFILLER_89_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ _19652_/Q _16993_/A _12205_/C vssd1 vssd1 vccd1 vccd1 _12256_/C sky130_fd_sc_hd__and3_1
XFILLER_89_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10255__S1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ _19608_/Q _12501_/X _12503_/X _19476_/Q _13184_/X vssd1 vssd1 vccd1 vccd1
+ _15572_/B sky130_fd_sc_hd__a221o_2
XFILLER_124_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10397_ _10390_/Y _10392_/Y _10394_/Y _10396_/Y _09830_/A vssd1 vssd1 vccd1 vccd1
+ _10397_/X sky130_fd_sc_hd__o221a_4
XFILLER_97_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19801_ _19802_/CLK _19801_/D vssd1 vssd1 vccd1 vccd1 _19801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12136_ _12126_/A _11963_/X _12129_/X _12135_/X vssd1 vssd1 vccd1 vccd1 _12136_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_2_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17993_ _17993_/A vssd1 vssd1 vccd1 vccd1 _19769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_151_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19732_ _19734_/CLK _19732_/D vssd1 vssd1 vccd1 vccd1 _19732_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_78_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16944_ _19632_/Q _16957_/B vssd1 vssd1 vccd1 vccd1 _16944_/X sky130_fd_sc_hd__or2_1
X_12067_ _12369_/A _12067_/B _12176_/B vssd1 vssd1 vccd1 vccd1 _12067_/X sky130_fd_sc_hd__or3_1
XFILLER_78_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16048__A0 _15522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11018_ _19175_/Q _18789_/Q _19239_/Q _18358_/Q _11149_/A _09512_/A vssd1 vssd1 vccd1
+ vccd1 _11019_/B sky130_fd_sc_hd__mux4_1
X_19663_ _19663_/CLK _19663_/D vssd1 vssd1 vccd1 vccd1 _19663_/Q sky130_fd_sc_hd__dfxtp_1
X_16875_ _16883_/A _16879_/C vssd1 vssd1 vccd1 vccd1 _16875_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18614_ _18917_/CLK _18614_/D vssd1 vssd1 vccd1 vccd1 _18614_/Q sky130_fd_sc_hd__dfxtp_1
X_15826_ _13576_/X _19253_/Q _15826_/S vssd1 vssd1 vccd1 vccd1 _15827_/A sky130_fd_sc_hd__mux2_1
X_19594_ _19594_/CLK _19594_/D vssd1 vssd1 vccd1 vccd1 _19594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18545_ _19268_/CLK _18545_/D vssd1 vssd1 vccd1 vccd1 _18545_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12085__A1 _11445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _13579_/X _19222_/Q _15765_/S vssd1 vssd1 vccd1 vccd1 _15758_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__A _18263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12969_ _19747_/Q vssd1 vssd1 vccd1 vccd1 _16039_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_61_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _14708_/A vssd1 vssd1 vccd1 vccd1 _18812_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18476_ _19197_/CLK _18476_/D vssd1 vssd1 vccd1 vccd1 _18476_/Q sky130_fd_sc_hd__dfxtp_1
X_15688_ _15688_/A vssd1 vssd1 vccd1 vccd1 _19191_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ _17596_/A vssd1 vssd1 vccd1 vccd1 _17427_/X sky130_fd_sc_hd__clkbuf_2
X_14639_ input44/X _18148_/A _18029_/A _14623_/X _18116_/A vssd1 vssd1 vccd1 vccd1
+ _18213_/B sky130_fd_sc_hd__a32o_1
XFILLER_158_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17358_ _17548_/B _17357_/X _17456_/S vssd1 vssd1 vccd1 vccd1 _17359_/A sky130_fd_sc_hd__mux2_1
XFILLER_119_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16309_ _19456_/Q _19457_/Q _19459_/Q _19458_/Q vssd1 vssd1 vccd1 vccd1 _16426_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_119_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17289_ _12383_/A _17463_/B _17293_/S vssd1 vssd1 vccd1 vccd1 _17289_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17720__B1 _17719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19028_ _19124_/CLK _19028_/D vssd1 vssd1 vccd1 vccd1 _19028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14821__S _14821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13945__B _14787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10650__A _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17787__A0 _17790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15652__S _15660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09614_ _09614_/A vssd1 vssd1 vccd1 vccd1 _09614_/X sky130_fd_sc_hd__buf_4
XFILLER_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09650__S _10785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09545_ _10721_/A vssd1 vssd1 vccd1 vccd1 _10680_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12577__A _17026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14268__S _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13172__S _13172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ _09476_/A vssd1 vssd1 vccd1 vccd1 _09477_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13900__S _13903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13132__D_N _12571_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_4_0_clock_A clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15099__S _15099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10320_ _19189_/Q _18803_/Q _19253_/Q _18372_/Q _09682_/A _10314_/A vssd1 vssd1 vccd1
+ vccd1 _10321_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_162_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10251_ _19318_/Q _18730_/Q _18767_/Q _18341_/Q _10247_/X _09712_/A vssd1 vssd1 vccd1
+ vccd1 _10251_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14731__S _14737_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10011__B1 _09485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10182_ _10182_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__nor2_1
XFILLER_132_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18019__A1 _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14990_ _18941_/Q vssd1 vssd1 vccd1 vccd1 _14991_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_93_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13941_ _13940_/X _18512_/Q _13941_/S vssd1 vssd1 vccd1 vccd1 _13942_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16660_ _16660_/A _16660_/B _16669_/D vssd1 vssd1 vccd1 vccd1 _19529_/D sky130_fd_sc_hd__nor3_1
XFILLER_35_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13872_ _13872_/A vssd1 vssd1 vccd1 vccd1 _18490_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _15611_/A vssd1 vssd1 vccd1 vccd1 _19164_/D sky130_fd_sc_hd__clkbuf_1
X_12823_ _16836_/B _12633_/X _12634_/X _16423_/B _12822_/X vssd1 vssd1 vccd1 vccd1
+ _13408_/B sky130_fd_sc_hd__a221o_4
X_16591_ _19511_/Q _16596_/C _16590_/X vssd1 vssd1 vccd1 vccd1 _16591_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14178__S _14180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12487__A _17294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13082__S _13143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18330_ _19306_/CLK _18330_/D vssd1 vssd1 vccd1 vccd1 _18330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10078__B1 _09833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15542_ _15519_/X _15540_/X _15541_/Y _15508_/X hold13/X vssd1 vssd1 vccd1 vccd1
+ _15542_/X sky130_fd_sc_hd__a32o_4
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11814__B2 _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12754_ hold13/A _12752_/X _10597_/A _12747_/X vssd1 vssd1 vccd1 vccd1 _18265_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10173__S0 _09904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16202__A0 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _19634_/Q _11705_/B vssd1 vssd1 vccd1 vccd1 _11706_/C sky130_fd_sc_hd__xnor2_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18261_ _19201_/CLK _18261_/D vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfxtp_2
X_12685_ _16706_/C _12507_/X _12511_/X _19511_/Q _12684_/X vssd1 vssd1 vccd1 vccd1
+ _12685_/X sky130_fd_sc_hd__a221o_1
X_15473_ _15473_/A vssd1 vssd1 vccd1 vccd1 _19140_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18174__A _18234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _17240_/S vssd1 vssd1 vccd1 vccd1 _17261_/S sky130_fd_sc_hd__clkbuf_2
X_14424_ _13912_/X _18700_/Q _14428_/S vssd1 vssd1 vccd1 vccd1 _14425_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _11681_/A _17239_/A vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__xnor2_4
X_18192_ _18233_/A vssd1 vssd1 vccd1 vccd1 _18231_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_129_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11578__B1 _19855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17143_ _17143_/A vssd1 vssd1 vccd1 vccd1 _19700_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14355_ _14355_/A vssd1 vssd1 vccd1 vccd1 _18670_/D sky130_fd_sc_hd__clkbuf_1
X_11567_ _11567_/A _11713_/B _17177_/A _11566_/X vssd1 vssd1 vccd1 vccd1 _11840_/A
+ sky130_fd_sc_hd__nor4b_4
XFILLER_156_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10476__S1 _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__A _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10518_ _18496_/Q _18991_/Q _10518_/S vssd1 vssd1 vccd1 vccd1 _10519_/A sky130_fd_sc_hd__mux2_1
X_13306_ _13306_/A _13306_/B vssd1 vssd1 vccd1 vccd1 _13306_/Y sky130_fd_sc_hd__nand2_1
XFILLER_143_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17074_ _17085_/A vssd1 vssd1 vccd1 vccd1 _17083_/S sky130_fd_sc_hd__clkbuf_2
X_14286_ input48/X _14282_/X _14277_/X _14278_/X _18125_/A vssd1 vssd1 vccd1 vccd1
+ _18220_/B sky130_fd_sc_hd__a32o_2
XFILLER_171_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11498_ _12832_/A vssd1 vssd1 vccd1 vccd1 _12861_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09618__S0 _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16025_ _16024_/X _19334_/Q _16025_/S vssd1 vssd1 vccd1 vccd1 _16026_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15737__S _15743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13237_ input16/X _13117_/X _13120_/X vssd1 vssd1 vccd1 vccd1 _13237_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_170_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10449_ _10461_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10449_/X sky130_fd_sc_hd__or2_1
XFILLER_171_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10002__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13168_ input11/X _13166_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _13168_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_152_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12119_ _12056_/A _12089_/A _12088_/A vssd1 vssd1 vccd1 vccd1 _12120_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11566__A _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15038__A _15038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ _19567_/Q _12518_/A _13098_/X _12707_/X vssd1 vssd1 vccd1 vccd1 _13099_/X
+ sky130_fd_sc_hd__a211o_1
X_17976_ _17976_/A vssd1 vssd1 vccd1 vccd1 _19761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19715_ _19724_/CLK _19715_/D vssd1 vssd1 vccd1 vccd1 _19715_/Q sky130_fd_sc_hd__dfxtp_4
X_16927_ input68/X _16929_/B vssd1 vssd1 vccd1 vccd1 _16927_/X sky130_fd_sc_hd__or2_1
XFILLER_66_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19646_ _19695_/CLK _19646_/D vssd1 vssd1 vccd1 vccd1 _19646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16858_ _16883_/A _16862_/C vssd1 vssd1 vccd1 vccd1 _16858_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15809_ _13551_/X _19245_/Q _15815_/S vssd1 vssd1 vccd1 vccd1 _15810_/A sky130_fd_sc_hd__mux2_1
X_19577_ _19583_/CLK _19577_/D vssd1 vssd1 vccd1 vccd1 _19577_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14088__S _14096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16789_ _16799_/A _16789_/B _16798_/D vssd1 vssd1 vccd1 vccd1 _19570_/D sky130_fd_sc_hd__nor3_1
XANTENNA__16992__A1 _15568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09330_ _11918_/B vssd1 vssd1 vccd1 vccd1 _12735_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__10069__B1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18528_ _19282_/CLK _18528_/D vssd1 vssd1 vccd1 vccd1 _18528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09261_ _12660_/B _12490_/A vssd1 vssd1 vccd1 vccd1 _09261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18459_ _19247_/CLK _18459_/D vssd1 vssd1 vccd1 vccd1 _18459_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16744__A1 _16752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18084__A _18097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09192_ _19854_/Q _19853_/Q _19852_/Q _19851_/Q vssd1 vssd1 vccd1 vccd1 _11522_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_14_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__A _19719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15647__S _15649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16332__A _16341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09645__S _09645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_152_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14787__A _18089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17163__A _17163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_109_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09528_ _10347_/A _09521_/Y _09527_/Y _09557_/A vssd1 vssd1 vccd1 vccd1 _09528_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _18478_/Q _19069_/Q _19231_/Q _18446_/Q _09980_/S _09390_/A vssd1 vssd1 vccd1
+ vccd1 _09459_/X sky130_fd_sc_hd__mux4_1
XPHY_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16735__A1 _16736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14726__S _14726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ _12474_/A _12470_/B vssd1 vssd1 vccd1 vccd1 _12470_/Y sky130_fd_sc_hd__nor2_1
XFILLER_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ _11419_/X _09664_/A _11420_/Y vssd1 vssd1 vccd1 vccd1 _11492_/D sky130_fd_sc_hd__a21o_2
XFILLER_138_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14140_ _14140_/A vssd1 vssd1 vccd1 vccd1 _18582_/D sky130_fd_sc_hd__clkbuf_1
X_11352_ _11441_/B vssd1 vssd1 vccd1 vccd1 _11352_/Y sky130_fd_sc_hd__inv_2
XFILLER_125_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _10303_/A _12468_/B vssd1 vssd1 vccd1 vccd1 _10304_/B sky130_fd_sc_hd__nor2_1
XFILLER_152_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14071_ _14071_/A vssd1 vssd1 vccd1 vccd1 _18552_/D sky130_fd_sc_hd__clkbuf_1
X_11283_ _11239_/A _11238_/A _11260_/X _12442_/B vssd1 vssd1 vccd1 vccd1 _11465_/D
+ sky130_fd_sc_hd__o22ai_2
XFILLER_152_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13022_ input2/X _12974_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _13022_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input51_A io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _09690_/A _10233_/X _10404_/A vssd1 vssd1 vccd1 vccd1 _10234_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11327__A3 _18829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17830_ _17830_/A vssd1 vssd1 vccd1 vccd1 _19729_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10290__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ _10158_/Y _10160_/Y _10162_/Y _10164_/Y _09831_/X vssd1 vssd1 vccd1 vccd1
+ _10165_/X sky130_fd_sc_hd__o221a_1
XFILLER_121_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17761_ _17937_/A vssd1 vssd1 vccd1 vccd1 _17761_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14973_ _14973_/A vssd1 vssd1 vccd1 vccd1 _18932_/D sky130_fd_sc_hd__clkbuf_1
X_10096_ _09715_/X _10093_/X _10095_/X vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19500_ _19619_/CLK _19500_/D vssd1 vssd1 vccd1 vccd1 _19500_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15292__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16712_ _19547_/Q _19546_/Q _19545_/Q _16712_/D vssd1 vssd1 vccd1 vccd1 _16722_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__13805__S _13809_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13924_ _13924_/A vssd1 vssd1 vccd1 vccd1 _18506_/D sky130_fd_sc_hd__clkbuf_1
X_17692_ _17648_/S _17505_/Y _17402_/A vssd1 vssd1 vccd1 vccd1 _17692_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19431_ _19524_/CLK _19431_/D vssd1 vssd1 vccd1 vccd1 _19431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_142_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16643_ _19525_/Q _16650_/B _16650_/C vssd1 vssd1 vccd1 vccd1 _16644_/B sky130_fd_sc_hd__and3_1
XANTENNA__17620__C1 _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13855_ _13854_/X _18485_/Q _13855_/S vssd1 vssd1 vccd1 vccd1 _13856_/A sky130_fd_sc_hd__mux2_1
XFILLER_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13106__A _15047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12806_ _19811_/Q _14297_/B vssd1 vssd1 vccd1 vccd1 _14998_/A sky130_fd_sc_hd__and2_1
X_19362_ _19736_/CLK _19362_/D vssd1 vssd1 vccd1 vccd1 _19362_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16574_ _19505_/Q _16575_/C _19506_/Q vssd1 vssd1 vccd1 vccd1 _16576_/B sky130_fd_sc_hd__a21oi_1
X_13786_ _13786_/A vssd1 vssd1 vccd1 vccd1 _18457_/D sky130_fd_sc_hd__clkbuf_1
X_10998_ _18390_/Q _18651_/Q _18550_/Q _18885_/Q _11011_/A _11012_/A vssd1 vssd1 vccd1
+ vccd1 _10999_/B sky130_fd_sc_hd__mux4_1
X_18313_ _19328_/CLK _18313_/D vssd1 vssd1 vccd1 vccd1 _18313_/Q sky130_fd_sc_hd__dfxtp_1
X_15525_ _15636_/S vssd1 vssd1 vccd1 vccd1 _15544_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12737_ _12737_/A vssd1 vssd1 vccd1 vccd1 _18255_/D sky130_fd_sc_hd__clkbuf_1
X_19293_ _19390_/CLK _19293_/D vssd1 vssd1 vccd1 vccd1 _19293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ input57/X _14274_/X _18229_/X _18234_/X _18144_/A vssd1 vssd1 vccd1 vccd1
+ _18245_/B sky130_fd_sc_hd__a32o_1
XFILLER_31_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15456_ _15456_/A vssd1 vssd1 vccd1 vccd1 _19133_/D sky130_fd_sc_hd__clkbuf_1
X_12668_ _12713_/A _18263_/Q vssd1 vssd1 vccd1 vccd1 _12668_/Y sky130_fd_sc_hd__nand2_1
XFILLER_169_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14407_ _14407_/A vssd1 vssd1 vccd1 vccd1 _18692_/D sky130_fd_sc_hd__clkbuf_1
X_18175_ input63/X _18155_/X _18168_/X _18174_/X _18087_/A vssd1 vssd1 vccd1 vccd1
+ _18176_/B sky130_fd_sc_hd__a32o_1
X_11619_ _11619_/A vssd1 vssd1 vccd1 vccd1 _18125_/A sky130_fd_sc_hd__buf_2
X_15387_ _19103_/Q _15098_/X _15387_/S vssd1 vssd1 vccd1 vccd1 _15388_/A sky130_fd_sc_hd__mux2_1
X_12599_ _19427_/Q _12600_/B _12606_/B vssd1 vssd1 vccd1 vccd1 _12599_/X sky130_fd_sc_hd__or3_1
XFILLER_128_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17126_ _18122_/A _17126_/B _17126_/C _17126_/D vssd1 vssd1 vccd1 vccd1 _17127_/B
+ sky130_fd_sc_hd__or4_1
X_14338_ _14338_/A vssd1 vssd1 vccd1 vccd1 _18662_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17057_ _19676_/Q _12669_/X _17061_/S vssd1 vssd1 vccd1 vccd1 _17058_/A sky130_fd_sc_hd__mux2_1
X_14269_ _14269_/A vssd1 vssd1 vccd1 vccd1 _18640_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16008_ _12130_/X _16007_/Y _13423_/B vssd1 vssd1 vccd1 vccd1 _16008_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11723__A0 _12447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_191_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19309_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12279__A1 _19416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17968_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_39_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_110_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__S0 _10339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19629_ _19663_/CLK _19629_/D vssd1 vssd1 vccd1 vccd1 _19629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17711__A _17910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09313_ _19708_/Q _09309_/X _09130_/X _09312_/Y vssd1 vssd1 vccd1 vccd1 _11702_/D
+ sky130_fd_sc_hd__o211a_4
XFILLER_90_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12451__A1 _18100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _19826_/Q _19825_/Q _19824_/Q _19823_/Q vssd1 vssd1 vccd1 vccd1 _09274_/C
+ sky130_fd_sc_hd__or4_2
XFILLER_22_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12203__A1 _19349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ _17117_/A _09338_/C _09175_/C vssd1 vssd1 vccd1 vccd1 _11556_/B sky130_fd_sc_hd__or3_2
XANTENNA__09604__C1 _09374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12754__A2 _12752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_144_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19235_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15377__S _15383_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11918__B _11918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16997__A _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__B2 _19722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__B1 _11632_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_159_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19364_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11190__A1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13625__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11934__A _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _11915_/A _11969_/B _11969_/D _11969_/C vssd1 vssd1 vccd1 vccd1 _11970_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10921_ _11024_/A vssd1 vssd1 vccd1 vccd1 _11116_/A sky130_fd_sc_hd__buf_2
XANTENNA__13219__B1 _13218_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11493__A2 _11492_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15840__S _15848_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13640_ _12981_/X _18393_/Q _13642_/S vssd1 vssd1 vccd1 vccd1 _13641_/A sky130_fd_sc_hd__mux2_1
X_10852_ _18489_/Q _18984_/Q _10852_/S vssd1 vssd1 vccd1 vccd1 _10853_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10128__S0 _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _18370_/Q _13570_/X _13577_/S vssd1 vssd1 vccd1 vccd1 _13572_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14456__S _14456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10783_ _18490_/Q _18985_/Q _11318_/S vssd1 vssd1 vccd1 vccd1 _10784_/A sky130_fd_sc_hd__mux2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15310_ _15310_/A vssd1 vssd1 vccd1 vccd1 _19068_/D sky130_fd_sc_hd__clkbuf_1
X_12522_ _12522_/A vssd1 vssd1 vccd1 vccd1 _13391_/A sky130_fd_sc_hd__buf_2
XFILLER_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16290_ _16298_/A _16290_/B vssd1 vssd1 vccd1 vccd1 _16291_/A sky130_fd_sc_hd__and2_1
XFILLER_13_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15241_ _19038_/Q _15095_/X _15243_/S vssd1 vssd1 vccd1 vccd1 _15242_/A sky130_fd_sc_hd__mux2_1
X_12453_ _12453_/A _12461_/B vssd1 vssd1 vccd1 vccd1 _12453_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11404_ _11404_/A _11404_/B vssd1 vssd1 vccd1 vccd1 _11404_/Y sky130_fd_sc_hd__nor2_1
X_12384_ _12385_/A _17899_/B vssd1 vssd1 vccd1 vccd1 _12387_/A sky130_fd_sc_hd__nand2_1
X_15172_ _15172_/A vssd1 vssd1 vccd1 vccd1 _19007_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11953__A0 _19783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15287__S _15289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11335_ _11335_/A _11335_/B vssd1 vssd1 vccd1 vccd1 _11335_/Y sky130_fd_sc_hd__nor2_1
X_14123_ _14123_/A vssd1 vssd1 vccd1 vccd1 _18576_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14191__S _14191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _19124_/CLK _18931_/D vssd1 vssd1 vccd1 vccd1 _18931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14054_ _14122_/S vssd1 vssd1 vccd1 vccd1 _14063_/S sky130_fd_sc_hd__clkbuf_4
X_11266_ _11266_/A _11266_/B vssd1 vssd1 vccd1 vccd1 _11266_/Y sky130_fd_sc_hd__nand2_1
X_13005_ _13005_/A vssd1 vssd1 vccd1 vccd1 _13005_/X sky130_fd_sc_hd__clkbuf_2
X_10217_ _18630_/Q _18965_/Q _10217_/S vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18862_ _19374_/CLK _18862_/D vssd1 vssd1 vccd1 vccd1 _18862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11197_ _18482_/Q _18977_/Q _11241_/S vssd1 vssd1 vccd1 vccd1 _11197_/X sky130_fd_sc_hd__mux2_1
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17813_ _17810_/A _17810_/B _17672_/A _17812_/Y vssd1 vssd1 vccd1 vccd1 _17813_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10148_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10148_/X sky130_fd_sc_hd__or2_1
X_18793_ _19180_/CLK _18793_/D vssd1 vssd1 vccd1 vccd1 _18793_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17744_ _17742_/X _17745_/B _17744_/S vssd1 vssd1 vccd1 vccd1 _17744_/X sky130_fd_sc_hd__mux2_1
X_14956_ _18924_/Q vssd1 vssd1 vccd1 vccd1 _14957_/A sky130_fd_sc_hd__clkbuf_1
X_10079_ _10080_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _11427_/A sky130_fd_sc_hd__or2_1
XFILLER_130_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13907_ _13905_/X _18501_/Q _13919_/S vssd1 vssd1 vccd1 vccd1 _13908_/A sky130_fd_sc_hd__mux2_1
X_17675_ _17479_/X _17674_/Y _17483_/X vssd1 vssd1 vccd1 vccd1 _17675_/X sky130_fd_sc_hd__a21o_1
XFILLER_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14887_ _18891_/Q _13985_/X _14893_/S vssd1 vssd1 vccd1 vccd1 _14888_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15750__S _15754_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19414_ _19423_/CLK _19414_/D vssd1 vssd1 vccd1 vccd1 _19414_/Q sky130_fd_sc_hd__dfxtp_2
X_16626_ _09241_/A _17133_/A _16626_/C _16626_/D vssd1 vssd1 vccd1 vccd1 _16659_/A
+ sky130_fd_sc_hd__and4bb_4
X_13838_ _19811_/Q _14297_/B vssd1 vssd1 vccd1 vccd1 _15854_/A sky130_fd_sc_hd__or2_2
XFILLER_51_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10119__S0 _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19345_ _19349_/CLK _19345_/D vssd1 vssd1 vccd1 vccd1 _19345_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_44_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16557_ hold3/A _16559_/C _16556_/Y vssd1 vssd1 vccd1 vccd1 _19499_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12433__A1 _12432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__A _19584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ _13769_/A vssd1 vssd1 vccd1 vccd1 _18449_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15051__A _15051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15508_ _15549_/A vssd1 vssd1 vccd1 vccd1 _15508_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19276_ _19370_/CLK _19276_/D vssd1 vssd1 vccd1 vccd1 _19276_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12984__A2 _12974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16488_ _19480_/Q _16485_/B _16487_/Y vssd1 vssd1 vccd1 vccd1 _19480_/D sky130_fd_sc_hd__o21a_1
XFILLER_148_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10995__B2 _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18227_ _18231_/A _18227_/B vssd1 vssd1 vccd1 vccd1 _18228_/A sky130_fd_sc_hd__and2_1
XFILLER_30_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19380_/CLK sky130_fd_sc_hd__clkbuf_16
X_15439_ _15439_/A vssd1 vssd1 vccd1 vccd1 _19125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10195__A _10195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18158_ _18158_/A vssd1 vssd1 vccd1 vccd1 _19837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17109_ _17109_/A _17109_/B _12462_/B vssd1 vssd1 vccd1 vccd1 _17169_/B sky130_fd_sc_hd__or3b_2
XFILLER_172_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18089_ _18089_/A _18091_/B vssd1 vssd1 vccd1 vccd1 _18089_/Y sky130_fd_sc_hd__nand2_1
XFILLER_132_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_171_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09931_ _18505_/Q _19000_/Q _09931_/S vssd1 vssd1 vccd1 vccd1 _09931_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_clock clkbuf_opt_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19383_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13161__A2 _12507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _19195_/Q _18809_/Q _19259_/Q _18378_/Q _09846_/X _09839_/A vssd1 vssd1 vccd1
+ vccd1 _09863_/B sky130_fd_sc_hd__mux4_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09460__S1 _10031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _10345_/A vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__clkbuf_2
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10358__S0 _09700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10132__C1 _09831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15660__S _15660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_14_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19292_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12585__A _16622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10530__S0 _10433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19385_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_167_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09227_ _19855_/Q _19810_/Q vssd1 vssd1 vccd1 vccd1 _09227_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09158_ _09158_/A _09158_/B _09211_/B vssd1 vssd1 vccd1 vccd1 _17168_/A sky130_fd_sc_hd__and3_1
XANTENNA__11086__S1 _11266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16626__B_N _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ _09207_/A vssd1 vssd1 vccd1 vccd1 _17175_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_163_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11120_ _19709_/Q vssd1 vssd1 vccd1 vccd1 _11120_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18076__C1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11051_ _09393_/A _11050_/X _11254_/A vssd1 vssd1 vccd1 vccd1 _11051_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15835__S _15837_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10002_ _09665_/A _09991_/X _10001_/X _09756_/A _19733_/Q vssd1 vssd1 vccd1 vccd1
+ _10082_/A sky130_fd_sc_hd__a32o_4
XFILLER_131_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14810_ _18857_/Q _13978_/X _14810_/S vssd1 vssd1 vccd1 vccd1 _14811_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15790_ _15790_/A vssd1 vssd1 vccd1 vccd1 _19236_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10349__S0 _10341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12479__B _12479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14741_ _14741_/A vssd1 vssd1 vccd1 vccd1 _18826_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input14_A io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12663__A1 _16778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10123__C1 _09813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__A2 _12443_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11953_ _19783_/Q _10648_/A _12028_/S vssd1 vssd1 vccd1 vccd1 _17221_/A sky130_fd_sc_hd__mux2_2
XFILLER_17_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17460_ _17844_/S vssd1 vssd1 vccd1 vccd1 _17710_/S sky130_fd_sc_hd__clkbuf_2
X_10904_ _11151_/S vssd1 vssd1 vccd1 vccd1 _10904_/X sky130_fd_sc_hd__clkbuf_4
X_14672_ _14560_/X _18796_/Q _14676_/S vssd1 vssd1 vccd1 vccd1 _14673_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11884_ _12074_/A vssd1 vssd1 vccd1 vccd1 _11884_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16411_ _19453_/Q _19452_/Q _16411_/C vssd1 vssd1 vccd1 vccd1 _16414_/B sky130_fd_sc_hd__and3_1
XFILLER_60_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13623_ _12801_/X _18385_/Q _13631_/S vssd1 vssd1 vccd1 vccd1 _13624_/A sky130_fd_sc_hd__mux2_1
X_17391_ _17391_/A vssd1 vssd1 vccd1 vccd1 _17739_/S sky130_fd_sc_hd__clkbuf_2
X_10835_ _11020_/A vssd1 vssd1 vccd1 vccd1 _11075_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19130_ _19386_/CLK _19130_/D vssd1 vssd1 vccd1 vccd1 _19130_/Q sky130_fd_sc_hd__dfxtp_1
X_16342_ _19431_/Q _19430_/Q _19429_/Q _16342_/D vssd1 vssd1 vccd1 vccd1 _16355_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_158_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13554_ _15038_/A vssd1 vssd1 vccd1 vccd1 _13554_/X sky130_fd_sc_hd__buf_2
X_10766_ _09671_/A _10763_/X _10765_/X vssd1 vssd1 vccd1 vccd1 _10766_/X sky130_fd_sc_hd__a21o_1
XFILLER_41_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19061_ _19619_/CLK _19061_/D vssd1 vssd1 vccd1 vccd1 _19061_/Q sky130_fd_sc_hd__dfxtp_1
X_12505_ _16879_/B _12501_/X _12503_/X _16466_/B vssd1 vssd1 vccd1 vccd1 _12542_/B
+ sky130_fd_sc_hd__a22o_2
X_16273_ _16273_/A vssd1 vssd1 vccd1 vccd1 _19405_/D sky130_fd_sc_hd__clkbuf_1
X_13485_ _13485_/A vssd1 vssd1 vccd1 vccd1 _18341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10697_ _10639_/X _10696_/X _10074_/A vssd1 vssd1 vccd1 vccd1 _10697_/X sky130_fd_sc_hd__o21a_1
XFILLER_157_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18012_ _19778_/Q _19399_/Q _18016_/S vssd1 vssd1 vccd1 vccd1 _18013_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15224_ _19030_/Q _15070_/X _15228_/S vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__mux2_1
X_12436_ _19359_/Q _12274_/B _12230_/X vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__o21a_1
XFILLER_138_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15155_ _15155_/A vssd1 vssd1 vccd1 vccd1 _18999_/D sky130_fd_sc_hd__clkbuf_1
X_12367_ _19659_/Q _12394_/C vssd1 vssd1 vccd1 vccd1 _12367_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14106_ _14106_/A vssd1 vssd1 vccd1 vccd1 _18568_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output82_A _11612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11318_ _18494_/Q _18989_/Q _11318_/S vssd1 vssd1 vccd1 vccd1 _11319_/A sky130_fd_sc_hd__mux2_1
X_12298_ _19656_/Q _17005_/A _12298_/C vssd1 vssd1 vccd1 vccd1 _12343_/C sky130_fd_sc_hd__and3_1
X_15086_ _15086_/A vssd1 vssd1 vccd1 vccd1 _15086_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11249_ _11254_/A _11246_/X _11248_/X _11134_/X vssd1 vssd1 vccd1 vccd1 _11249_/X
+ sky130_fd_sc_hd__o211a_1
X_18914_ _19736_/CLK _18914_/D vssd1 vssd1 vccd1 vccd1 _18914_/Q sky130_fd_sc_hd__dfxtp_1
X_14037_ _18540_/Q _14036_/X _14043_/S vssd1 vssd1 vccd1 vccd1 _14038_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10750__A_N _10749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18845_ _19389_/CLK _18845_/D vssd1 vssd1 vccd1 vccd1 _18845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17290__A0 _12358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18776_ _19375_/CLK _18776_/D vssd1 vssd1 vccd1 vccd1 _18776_/Q sky130_fd_sc_hd__dfxtp_1
X_15988_ _13602_/X _19325_/Q _15992_/S vssd1 vssd1 vccd1 vccd1 _15989_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17727_ _17722_/A _17722_/B _17530_/A _17726_/X vssd1 vssd1 vccd1 vccd1 _17727_/X
+ sky130_fd_sc_hd__o211a_1
X_14939_ _14939_/A vssd1 vssd1 vccd1 vccd1 _18915_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_82_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_0_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17658_ _17717_/S _17657_/Y _17402_/A vssd1 vssd1 vccd1 vccd1 _17658_/X sky130_fd_sc_hd__a21o_1
XFILLER_35_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16609_ _19517_/Q _19516_/Q _16609_/C vssd1 vssd1 vccd1 vccd1 _16613_/B sky130_fd_sc_hd__and3_1
XFILLER_90_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14096__S _14096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17589_ _17672_/A vssd1 vssd1 vccd1 vccd1 _17589_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19328_ _19328_/CLK _19328_/D vssd1 vssd1 vccd1 vccd1 _19328_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09283__B1 _19584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19259_ _19391_/CLK _19259_/D vssd1 vssd1 vccd1 vccd1 _19259_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14824__S _14832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16305__C1 _16914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10653__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09219__A _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09914_ _10174_/A _09914_/B vssd1 vssd1 vccd1 vccd1 _09914_/Y sky130_fd_sc_hd__nor2_1
XFILLER_120_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11145__A1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09845_ _09839_/X _09842_/X _09843_/X _10108_/A _09844_/X vssd1 vssd1 vccd1 vccd1
+ _09859_/B sky130_fd_sc_hd__o221a_1
XFILLER_98_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input6_A io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11240__S1 _11124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09776_/A vssd1 vssd1 vccd1 vccd1 _10520_/S sky130_fd_sc_hd__buf_2
XFILLER_27_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12645__A1 _16772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13903__S _13903_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15595__A0 _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10620_ _09369_/A _10610_/X _10619_/X _09472_/A _19719_/Q vssd1 vssd1 vccd1 vccd1
+ _10648_/A sky130_fd_sc_hd__a32o_2
XFILLER_169_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10959__B2 _19713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10551_ _10823_/A vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10423__A3 _10422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10482_/Y sky130_fd_sc_hd__nand2_1
X_13270_ _19732_/Q _15598_/B _13381_/S vssd1 vssd1 vccd1 vccd1 _13270_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12221_ _12221_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12224_/A sky130_fd_sc_hd__nor2_2
XFILLER_136_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12152_ _12322_/A _12322_/B _12149_/A vssd1 vssd1 vccd1 vccd1 _12152_/X sky130_fd_sc_hd__a21o_1
X_11103_ _18914_/Q _18680_/Q _19362_/Q _19010_/Q _09624_/A _11020_/X vssd1 vssd1 vccd1
+ vccd1 _11104_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13874__A _13941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ _17013_/A vssd1 vssd1 vccd1 vccd1 _16971_/B sky130_fd_sc_hd__clkbuf_1
X_12083_ _17756_/B _12053_/B _12241_/A vssd1 vssd1 vccd1 vccd1 _12084_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11136__A1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11034_ _18614_/Q _18949_/Q _11071_/S vssd1 vssd1 vccd1 vccd1 _11034_/X sky130_fd_sc_hd__mux2_1
X_15911_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15920_/S sky130_fd_sc_hd__clkbuf_4
X_16891_ _16891_/A vssd1 vssd1 vccd1 vccd1 _16896_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12884__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__S1 _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12884__B2 _12798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18630_ _19096_/CLK _18630_/D vssd1 vssd1 vccd1 vccd1 _18630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15842_ _13599_/X _19260_/Q _15848_/S vssd1 vssd1 vccd1 vccd1 _15843_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18561_ _19282_/CLK _18561_/D vssd1 vssd1 vccd1 vccd1 _18561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ _15773_/A vssd1 vssd1 vccd1 vccd1 _19229_/D sky130_fd_sc_hd__clkbuf_1
X_12985_ _13033_/A vssd1 vssd1 vccd1 vccd1 _13154_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ _17361_/X _17355_/X _17512_/S vssd1 vssd1 vccd1 vccd1 _17512_/X sky130_fd_sc_hd__mux2_1
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_157_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14724_ _14531_/X _18819_/Q _14726_/S vssd1 vssd1 vccd1 vccd1 _14725_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09799__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ _19339_/Q _11766_/X _12037_/A _11935_/X _16109_/A vssd1 vssd1 vccd1 vccd1
+ _11936_/X sky130_fd_sc_hd__o221a_1
XFILLER_27_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18492_ _18987_/CLK _18492_/D vssd1 vssd1 vccd1 vccd1 _18492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10742__S0 _11297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _17437_/X _17653_/B _17573_/S vssd1 vssd1 vccd1 vccd1 _17444_/A sky130_fd_sc_hd__mux2_1
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14655_ _14655_/A vssd1 vssd1 vccd1 vccd1 _18788_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11890_/B vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__buf_2
XFILLER_159_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13606_ _18381_/Q _13605_/X _13609_/S vssd1 vssd1 vccd1 vccd1 _13607_/A sky130_fd_sc_hd__mux2_1
X_10818_ _19274_/Q _19112_/Q _18521_/Q _18291_/Q _11049_/S _10817_/X vssd1 vssd1 vccd1
+ vccd1 _10819_/B sky130_fd_sc_hd__mux4_1
X_17374_ _17290_/X _17285_/X _17375_/S vssd1 vssd1 vccd1 vccd1 _17374_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14586_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14599_/S sky130_fd_sc_hd__buf_4
X_11798_ _19334_/Q _11653_/X _15488_/A vssd1 vssd1 vccd1 vccd1 _11798_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_159_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19113_ _19113_/CLK _19113_/D vssd1 vssd1 vccd1 vccd1 _19113_/Q sky130_fd_sc_hd__dfxtp_2
X_16325_ _16333_/D vssd1 vssd1 vccd1 vccd1 _16331_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13537_ _13537_/A vssd1 vssd1 vccd1 vccd1 _18359_/D sky130_fd_sc_hd__clkbuf_1
X_10749_ _12455_/B _10749_/B vssd1 vssd1 vccd1 vccd1 _10751_/A sky130_fd_sc_hd__and2b_1
XFILLER_174_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16425__A _16442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19044_ _19237_/CLK _19044_/D vssd1 vssd1 vccd1 vccd1 _19044_/Q sky130_fd_sc_hd__dfxtp_1
X_16256_ _16256_/A vssd1 vssd1 vccd1 vccd1 _19398_/D sky130_fd_sc_hd__clkbuf_1
X_13468_ _13070_/X _18334_/Q _13470_/S vssd1 vssd1 vccd1 vccd1 _13469_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15207_ _15207_/A vssd1 vssd1 vccd1 vccd1 _19022_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09568__A1 _09557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12419_/A _17906_/B vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__nand2_1
XFILLER_127_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16187_ _13538_/X _19367_/Q _16191_/S vssd1 vssd1 vccd1 vccd1 _16188_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ hold21/A _13399_/B vssd1 vssd1 vccd1 vccd1 _13399_/X sky130_fd_sc_hd__or2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15138_ _15138_/A vssd1 vssd1 vccd1 vccd1 _18991_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11288__B _12449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10583__C1 _09811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15510__A0 _19715_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__A2 _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15069_ _15069_/A vssd1 vssd1 vccd1 vccd1 _18965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11222__S1 _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09630_ _09630_/A vssd1 vssd1 vccd1 vccd1 _09630_/X sky130_fd_sc_hd__buf_2
XFILLER_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18828_ _19054_/CLK _18828_/D vssd1 vssd1 vccd1 vccd1 _18828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09561_ _09561_/A vssd1 vssd1 vccd1 vccd1 _09630_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18759_ _19054_/CLK _18759_/D vssd1 vssd1 vccd1 vccd1 _18759_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18087__A _18087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14819__S _14821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13723__S _13725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09492_ _09644_/A vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__buf_2
XANTENNA__09502__A _11033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10648__A _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11243__S _11243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13024__A _15031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_4_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16335__A _16344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13355__A2 _12606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09654__S1 _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10574__C1 _09644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15385__S _15387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13694__A _13762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17166__A _17166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11926__B _17201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09828_ _09817_/A _09827_/X _09767_/X vssd1 vssd1 vccd1 vccd1 _09828_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_111_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10972__S0 _10969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09759_ _09667_/X _09742_/X _09755_/X _09758_/X _19735_/Q vssd1 vssd1 vccd1 vccd1
+ _11416_/A sky130_fd_sc_hd__a32o_4
XANTENNA__14729__S _14737_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10629__B1 _09640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _18276_/Q _12766_/X _09975_/A _12769_/X vssd1 vssd1 vccd1 vccd1 _18276_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09412__A _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _19846_/Q _11720_/X _11721_/S vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__mux2_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14440_ _14440_/A vssd1 vssd1 vccd1 vccd1 _18707_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_120_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11652_ _11652_/A vssd1 vssd1 vccd1 vccd1 _11859_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10603_ _18493_/Q _18988_/Q _10603_/S vssd1 vssd1 vccd1 vccd1 _10603_/X sky130_fd_sc_hd__mux2_1
XFILLER_80_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14371_ _14642_/D _14371_/B _14715_/C vssd1 vssd1 vccd1 vccd1 _15173_/B sky130_fd_sc_hd__or3_1
XANTENNA__10992__S _11243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11583_ _19862_/Q vssd1 vssd1 vccd1 vccd1 _18138_/A sky130_fd_sc_hd__buf_4
XFILLER_7_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12773__A _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16245__A _16245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ _16116_/B _16108_/Y _16109_/X vssd1 vssd1 vccd1 vccd1 _16110_/Y sky130_fd_sc_hd__a21oi_1
X_13322_ _19580_/Q _13055_/X _13321_/X _13265_/X vssd1 vssd1 vccd1 vccd1 _13322_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_156_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17090_ _19691_/Q _15615_/X _17094_/S vssd1 vssd1 vccd1 vccd1 _17091_/A sky130_fd_sc_hd__mux2_1
X_10534_ _18464_/Q _19055_/Q _19217_/Q _18432_/Q _10433_/S _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10535_/B sky130_fd_sc_hd__mux4_1
XFILLER_7_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16041_ _16046_/B _16041_/B vssd1 vssd1 vccd1 vccd1 _16041_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13253_ _13253_/A vssd1 vssd1 vccd1 vccd1 _18307_/D sky130_fd_sc_hd__clkbuf_1
X_10465_ _19282_/Q _19120_/Q _18529_/Q _18299_/Q _10500_/S _09672_/A vssd1 vssd1 vccd1
+ vccd1 _10466_/B sky130_fd_sc_hd__mux4_1
X_12204_ _16993_/A _12205_/C _19652_/Q vssd1 vssd1 vccd1 vccd1 _12204_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_136_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13184_ _16697_/C _12952_/X _12511_/X _19508_/Q _13183_/X vssd1 vssd1 vccd1 vccd1
+ _13184_/X sky130_fd_sc_hd__a221o_1
X_10396_ _10378_/A _10395_/X _10297_/X vssd1 vssd1 vccd1 vccd1 _10396_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_83_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19800_ _19800_/CLK _19800_/D vssd1 vssd1 vccd1 vccd1 _19800_/Q sky130_fd_sc_hd__dfxtp_1
X_12135_ _12130_/X _12132_/X _12133_/Y _12134_/X vssd1 vssd1 vccd1 vccd1 _12135_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17992_ _19769_/Q _19801_/Q _17994_/S vssd1 vssd1 vccd1 vccd1 _17993_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16943_ _17010_/A vssd1 vssd1 vccd1 vccd1 _16943_/X sky130_fd_sc_hd__clkbuf_2
X_19731_ _19731_/CLK _19731_/D vssd1 vssd1 vccd1 vccd1 _19731_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_111_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12066_ _12066_/A _12066_/B _12066_/C vssd1 vssd1 vccd1 vccd1 _12176_/B sky130_fd_sc_hd__and3_1
XFILLER_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14059__A0 _13848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _11263_/S vssd1 vssd1 vccd1 vccd1 _11149_/A sky130_fd_sc_hd__buf_4
XFILLER_65_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19662_ _19695_/CLK _19662_/D vssd1 vssd1 vccd1 vccd1 _19662_/Q sky130_fd_sc_hd__dfxtp_1
X_16874_ _16874_/A vssd1 vssd1 vccd1 vccd1 _16879_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10232__S _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17796__A1 _12149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15825_ _15825_/A vssd1 vssd1 vccd1 vccd1 _19252_/D sky130_fd_sc_hd__clkbuf_1
X_18613_ _19076_/CLK _18613_/D vssd1 vssd1 vccd1 vccd1 _18613_/Q sky130_fd_sc_hd__dfxtp_1
X_19593_ _19688_/CLK _19593_/D vssd1 vssd1 vccd1 vccd1 _19593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15767_/A vssd1 vssd1 vccd1 vccd1 _15765_/S sky130_fd_sc_hd__buf_4
X_18544_ _19297_/CLK _18544_/D vssd1 vssd1 vccd1 vccd1 _18544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12968_ _19715_/Q _15505_/B _13381_/S vssd1 vssd1 vccd1 vccd1 _12968_/X sky130_fd_sc_hd__mux2_1
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10096__A1 _09715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15559__A0 _19724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14707_ _14611_/X _18812_/Q _14709_/S vssd1 vssd1 vccd1 vccd1 _14708_/A sky130_fd_sc_hd__mux2_1
X_11919_ _12159_/B vssd1 vssd1 vccd1 vccd1 _11919_/Y sky130_fd_sc_hd__inv_2
X_18475_ _19387_/CLK _18475_/D vssd1 vssd1 vccd1 vccd1 _18475_/Q sky130_fd_sc_hd__dfxtp_1
X_15687_ _14589_/X _19191_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15688_/A sky130_fd_sc_hd__mux2_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12899_ _16340_/B _12700_/X _12898_/X vssd1 vssd1 vccd1 vccd1 _12899_/X sky130_fd_sc_hd__o21a_1
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17426_ _17432_/A _17726_/A vssd1 vssd1 vccd1 vccd1 _17596_/A sky130_fd_sc_hd__nor2_1
X_14638_ _18229_/A vssd1 vssd1 vccd1 vccd1 _18029_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__13034__B2 _13234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17357_ _17355_/X _17356_/X _17512_/S vssd1 vssd1 vccd1 vccd1 _17357_/X sky130_fd_sc_hd__mux2_1
X_14569_ _14569_/A vssd1 vssd1 vccd1 vccd1 _14569_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10399__A2 _10388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16308_ _19423_/Q _12440_/A _12437_/X _12440_/Y _12556_/X vssd1 vssd1 vccd1 vccd1
+ _19423_/D sky130_fd_sc_hd__o221a_1
XFILLER_158_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17288_ _17284_/X _17287_/X _17448_/S vssd1 vssd1 vccd1 vccd1 _17288_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19027_ _19027_/CLK _19027_/D vssd1 vssd1 vccd1 vccd1 _19027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16239_ _13614_/X _19391_/Q _16239_/S vssd1 vssd1 vccd1 vccd1 _16240_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10020__A1 _09768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09961__A1 _09964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10931__A _19714_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clock_A clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15933__S _15937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17787__A1 _17790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09931__S _09931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15798__A0 _13535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09613_ _10614_/A _09612_/X _09450_/A vssd1 vssd1 vccd1 vccd1 _09613_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09544_ _18606_/Q _18877_/Q _19101_/Q _18845_/Q _10479_/S _09768_/A vssd1 vssd1 vccd1
+ vccd1 _09544_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12577__B _12577_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09475_ _18742_/Q _09474_/Y _09230_/B _09223_/B vssd1 vssd1 vccd1 vccd1 _09476_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__10378__A _10378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12593__A _17026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11131__S0 _10878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_105_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_8_0_clock_A clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11002__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ _10250_/A vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10011__A1 _10289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17475__B1 _09322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10181_ _10181_/A _12471_/B vssd1 vssd1 vccd1 vccd1 _10182_/B sky130_fd_sc_hd__nor2_1
XFILLER_160_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12839__A1 _16736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13940_ _14620_/A vssd1 vssd1 vccd1 vccd1 _13940_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10945__S0 _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15789__A0 _13522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13871_ _13870_/X _18490_/Q _13871_/S vssd1 vssd1 vccd1 vccd1 _13872_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15610_ _15609_/X _19164_/Q _15627_/S vssd1 vssd1 vccd1 vccd1 _15611_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12822_ _19521_/Q _12782_/X _12699_/X _19489_/Q _12821_/X vssd1 vssd1 vccd1 vccd1
+ _12822_/X sky130_fd_sc_hd__a221o_1
X_16590_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16590_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13264__B2 _19353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__B _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10078__A1 _09760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15541_ _15541_/A hold13/A vssd1 vssd1 vccd1 vccd1 _15541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_opt_3_0_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_12753_ hold11/A _12752_/X _11342_/A _12747_/X vssd1 vssd1 vccd1 vccd1 _18264_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10288__A _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10173__S1 _09905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11704_ _09296_/X _11801_/B _11703_/X _11698_/B vssd1 vssd1 vccd1 vccd1 _11705_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _19720_/CLK _18260_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_2
X_15472_ _15471_/Y _19140_/Q _15483_/S vssd1 vssd1 vccd1 vccd1 _15473_/A sky130_fd_sc_hd__mux2_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _19447_/Q _12515_/X _12683_/X vssd1 vssd1 vccd1 vccd1 _12684_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17211_ _17211_/A vssd1 vssd1 vccd1 vccd1 _17743_/B sky130_fd_sc_hd__clkbuf_2
X_14423_ _14423_/A vssd1 vssd1 vccd1 vccd1 _18699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13599__A _15083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18191_ _18191_/A vssd1 vssd1 vccd1 vccd1 _19846_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11635_ _19773_/Q _11284_/A _11678_/A vssd1 vssd1 vccd1 vccd1 _17239_/A sky130_fd_sc_hd__mux2_8
XFILLER_168_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17142_ _17142_/A _17142_/B vssd1 vssd1 vccd1 vccd1 _17143_/A sky130_fd_sc_hd__and2_1
XANTENNA__12775__B1 _11418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14354_ _13918_/X _18670_/Q _14354_/S vssd1 vssd1 vccd1 vccd1 _14355_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11566_ _11566_/A _17105_/A _11566_/C _11589_/B vssd1 vssd1 vccd1 vccd1 _11566_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_11_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13305_ _19615_/Q _12950_/X _12951_/X _19483_/Q _13304_/X vssd1 vssd1 vccd1 vccd1
+ _13306_/B sky130_fd_sc_hd__a221o_2
XFILLER_116_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15713__A0 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17073_ _17073_/A vssd1 vssd1 vccd1 vccd1 _19683_/D sky130_fd_sc_hd__clkbuf_1
X_10517_ _09666_/A _10507_/X _10516_/X _09757_/A _19722_/Q vssd1 vssd1 vccd1 vccd1
+ _11347_/A sky130_fd_sc_hd__a32o_4
XFILLER_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14285_ _14285_/A vssd1 vssd1 vccd1 vccd1 _18642_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14922__S _14926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11497_ _18743_/Q vssd1 vssd1 vccd1 vccd1 _12832_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_109_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09618__S1 _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16024_ _15495_/X _16023_/Y _16024_/S vssd1 vssd1 vccd1 vccd1 _16024_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13236_ _13153_/A _13235_/X _13164_/X vssd1 vssd1 vccd1 vccd1 _13236_/Y sky130_fd_sc_hd__a21oi_1
X_10448_ _18928_/Q _18694_/Q _19376_/Q _19024_/Q _10451_/S _10311_/A vssd1 vssd1 vccd1
+ vccd1 _10449_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10538__C1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10002__A1 _09665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15319__A _15387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10002__B2 _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ _13167_/A vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__clkbuf_2
X_10379_ _18499_/Q _18994_/Q _10435_/S vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12118_ _12118_/A _12118_/B vssd1 vssd1 vccd1 vccd1 _12122_/A sky130_fd_sc_hd__and2_1
XFILLER_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13098_ _19153_/Q _12895_/X _12677_/X _19343_/Q _13097_/X vssd1 vssd1 vccd1 vccd1
+ _13098_/X sky130_fd_sc_hd__a221o_1
XFILLER_97_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17975_ _19761_/Q _19793_/Q _17979_/S vssd1 vssd1 vccd1 vccd1 _17976_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11189__S0 _10873_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19714_ _19724_/CLK _19714_/D vssd1 vssd1 vccd1 vccd1 _19714_/Q sky130_fd_sc_hd__dfxtp_4
X_16926_ _19626_/Q _12674_/X _16925_/X _16269_/X vssd1 vssd1 vccd1 vccd1 _19626_/D
+ sky130_fd_sc_hd__o211a_1
X_12049_ _12110_/A vssd1 vssd1 vccd1 vccd1 _17756_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_120_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19645_ _19645_/CLK _19645_/D vssd1 vssd1 vccd1 vccd1 _19645_/Q sky130_fd_sc_hd__dfxtp_1
X_16857_ _16857_/A vssd1 vssd1 vccd1 vccd1 _16862_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14369__S _14369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15054__A _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15808_ _15808_/A vssd1 vssd1 vccd1 vccd1 _19244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19576_ _19581_/CLK _19576_/D vssd1 vssd1 vccd1 vccd1 _19576_/Q sky130_fd_sc_hd__dfxtp_1
X_16788_ _19570_/Q _19569_/Q _19568_/Q _16788_/D vssd1 vssd1 vccd1 vccd1 _16798_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__14452__A0 _13848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13255__A1 input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10069__A1 _10590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15739_ _13554_/X _19214_/Q _15743_/S vssd1 vssd1 vccd1 vccd1 _15740_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18527_ _19280_/CLK _18527_/D vssd1 vssd1 vccd1 vccd1 _18527_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18194__B2 _17114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09260_ _12602_/B _12605_/B vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__nor2_2
X_18458_ _19180_/CLK _18458_/D vssd1 vssd1 vccd1 vccd1 _18458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ _19810_/Q vssd1 vssd1 vccd1 vccd1 _14297_/B sky130_fd_sc_hd__buf_4
X_17409_ _17800_/A vssd1 vssd1 vccd1 vccd1 _17724_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18389_ _19237_/CLK _18389_/D vssd1 vssd1 vccd1 vccd1 _18389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10137__S _10137_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14832__S _14832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10529__C1 _09812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13448__S _13448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18250__D input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09227__A _19855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__clkbuf_2
XFILLER_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15663__S _15671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14787__B _14787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_31_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09527_ _10347_/A _09527_/B vssd1 vssd1 vccd1 vccd1 _09527_/Y sky130_fd_sc_hd__nand2_1
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18185__B2 _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09897__A _09905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09458_ _09981_/S vssd1 vssd1 vccd1 vccd1 _09980_/S sky130_fd_sc_hd__clkbuf_4
XPHY_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14746__A1 _18829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10836__A _11075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09389_ _18638_/Q _18973_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12757__B1 _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ _11420_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11420_/Y sky130_fd_sc_hd__nand2_1
XFILLER_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11351_ _11351_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _11441_/B sky130_fd_sc_hd__nand2_1
XFILLER_125_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14742__S _14748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10302_ _10303_/A _12468_/B vssd1 vssd1 vccd1 vccd1 _10304_/A sky130_fd_sc_hd__and2_1
X_14070_ _13864_/X _18552_/Q _14074_/S vssd1 vssd1 vccd1 vccd1 _14071_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11282_ _09476_/A _11272_/X _11281_/X _09576_/A _09311_/Y vssd1 vssd1 vccd1 vccd1
+ _12442_/B sky130_fd_sc_hd__o32a_4
XFILLER_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13182__B1 _13181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13021_ _13153_/A _13017_/X _13020_/X vssd1 vssd1 vccd1 vccd1 _13021_/X sky130_fd_sc_hd__a21bo_1
XFILLER_152_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10233_ _18501_/Q _18996_/Q _10368_/S vssd1 vssd1 vccd1 vccd1 _10233_/X sky130_fd_sc_hd__mux2_1
XFILLER_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17999__A1 _19393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input44_A io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10164_ _10158_/A _10163_/X _09823_/A vssd1 vssd1 vccd1 vccd1 _10164_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10091__S0 _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09137__A _19864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14972_ _18932_/Q vssd1 vssd1 vccd1 vccd1 _14973_/A sky130_fd_sc_hd__clkbuf_1
X_10095_ _10138_/A _10094_/X _10150_/A vssd1 vssd1 vccd1 vccd1 _10095_/X sky130_fd_sc_hd__a21o_1
X_17760_ _17646_/X _17741_/X _17759_/X _17386_/X vssd1 vssd1 vccd1 vccd1 _17760_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_48_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__S0 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16711_ _16715_/C _16715_/D _19547_/Q vssd1 vssd1 vccd1 vccd1 _16713_/B sky130_fd_sc_hd__a21oi_1
X_13923_ _13921_/X _18506_/Q _13935_/S vssd1 vssd1 vccd1 vccd1 _13924_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17691_ _17691_/A vssd1 vssd1 vccd1 vccd1 _19718_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12498__A _17026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14189__S _14191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19430_ _19436_/CLK _19430_/D vssd1 vssd1 vccd1 vccd1 _19430_/Q sky130_fd_sc_hd__dfxtp_1
X_16642_ _16642_/A _16642_/B vssd1 vssd1 vccd1 vccd1 _19524_/D sky130_fd_sc_hd__nor2_1
X_13854_ _14534_/A vssd1 vssd1 vccd1 vccd1 _13854_/X sky130_fd_sc_hd__buf_2
XANTENNA__13237__A1 input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _13435_/B vssd1 vssd1 vccd1 vccd1 _14642_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16573_ _19505_/Q _16575_/C _16572_/Y vssd1 vssd1 vccd1 vccd1 _19505_/D sky130_fd_sc_hd__o21a_1
X_19361_ _19361_/CLK _19361_/D vssd1 vssd1 vccd1 vccd1 _19361_/Q sky130_fd_sc_hd__dfxtp_1
X_13785_ _12981_/X _18457_/Q _13787_/S vssd1 vssd1 vccd1 vccd1 _13786_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10997_ _18781_/Q vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__buf_2
XFILLER_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15524_ _19717_/Q _15522_/X _15543_/S vssd1 vssd1 vccd1 vccd1 _15524_/X sky130_fd_sc_hd__mux2_1
X_18312_ _19375_/CLK _18312_/D vssd1 vssd1 vccd1 vccd1 _18312_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16187__A0 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ _18255_/Q _12735_/X _17520_/S vssd1 vssd1 vccd1 vccd1 _12737_/A sky130_fd_sc_hd__mux2_1
X_19292_ _19292_/CLK _19292_/D vssd1 vssd1 vccd1 vccd1 _19292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18243_ _18243_/A vssd1 vssd1 vccd1 vccd1 _19864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09600__A _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15455_ _19133_/Q _15092_/X _15455_/S vssd1 vssd1 vccd1 vccd1 _15456_/A sky130_fd_sc_hd__mux2_1
X_12667_ _18263_/Q _12667_/B vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__or2_1
XANTENNA__12748__B1 _10749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14406_ _13886_/X _18692_/Q _14406_/S vssd1 vssd1 vccd1 vccd1 _14407_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18174_ _18234_/A vssd1 vssd1 vccd1 vccd1 _18174_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11618_ _11618_/A vssd1 vssd1 vccd1 vccd1 _18127_/A sky130_fd_sc_hd__buf_2
X_15386_ _15386_/A vssd1 vssd1 vccd1 vccd1 _19102_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09613__B1 _09450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ _19620_/Q _16245_/A vssd1 vssd1 vccd1 vccd1 _12598_/X sky130_fd_sc_hd__or2_1
XFILLER_128_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10759__C1 _09602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15748__S _15754_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17125_ _17125_/A _18127_/A _18125_/A _18140_/A vssd1 vssd1 vccd1 vccd1 _17126_/D
+ sky130_fd_sc_hd__or4bb_1
X_14337_ _13893_/X _18662_/Q _14343_/S vssd1 vssd1 vccd1 vccd1 _14338_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14652__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11549_ _11738_/A vssd1 vssd1 vccd1 vccd1 _12179_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_144_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16433__A _16442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ _17056_/A vssd1 vssd1 vccd1 vccd1 _19675_/D sky130_fd_sc_hd__clkbuf_1
X_14268_ _18640_/Q _14048_/X _14268_/S vssd1 vssd1 vccd1 vccd1 _14269_/A sky130_fd_sc_hd__mux2_1
X_16007_ _16011_/A _16011_/C vssd1 vssd1 vccd1 vccd1 _16007_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_83_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13219_ _19574_/Q _13006_/X _13218_/X _13012_/X vssd1 vssd1 vccd1 vccd1 _13219_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_171_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14199_ _14255_/A vssd1 vssd1 vccd1 vccd1 _14268_/S sky130_fd_sc_hd__buf_6
XFILLER_140_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12920__A0 _19713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A1 _11722_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17958_/A vssd1 vssd1 vccd1 vccd1 _19753_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18079__B _18079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16909_ _19615_/Q _16906_/B _16908_/Y vssd1 vssd1 vccd1 vccd1 _19615_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14099__S _14107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17889_ _17920_/B _17889_/B vssd1 vssd1 vccd1 vccd1 _17889_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10385__S1 _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19628_ _19828_/CLK _19628_/D vssd1 vssd1 vccd1 vccd1 _19628_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11743__C _11743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12201__A _19413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19559_ _19564_/CLK _19559_/D vssd1 vssd1 vccd1 vccd1 _19559_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11334__S0 _10572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09312_ _19705_/Q _09311_/Y _19706_/Q vssd1 vssd1 vccd1 vccd1 _09312_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16178__A0 _13525_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09510__A _18642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _19699_/Q vssd1 vssd1 vccd1 vccd1 _12543_/B sky130_fd_sc_hd__buf_2
XFILLER_166_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09174_ _09174_/A _09174_/B vssd1 vssd1 vccd1 vccd1 _17117_/A sky130_fd_sc_hd__nand2_2
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15658__S _15660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12590__B _12590_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10517__A2 _10507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17174__A _17174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10920_ _10920_/A vssd1 vssd1 vccd1 vccd1 _11024_/A sky130_fd_sc_hd__buf_2
XFILLER_147_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _10962_/S vssd1 vssd1 vccd1 vccd1 _10852_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__14737__S _14737_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10128__S1 _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__S0 _10692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11950__A _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _15054_/A vssd1 vssd1 vccd1 vccd1 _13570_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10775_/Y _10777_/Y _10779_/Y _10781_/Y _09571_/A vssd1 vssd1 vccd1 vccd1
+ _10782_/X sky130_fd_sc_hd__o221a_2
XANTENNA__17905__A1 _19736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A vssd1 vssd1 vccd1 vccd1 _12565_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10453__A1 _09674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15240_ _15240_/A vssd1 vssd1 vccd1 vccd1 _19037_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15392__A1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12452_ _12462_/B vssd1 vssd1 vccd1 vccd1 _12461_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11403_ _19201_/Q _18815_/Q _19265_/Q _18384_/Q _11388_/S _09788_/A vssd1 vssd1 vccd1
+ vccd1 _11404_/B sky130_fd_sc_hd__mux4_1
X_15171_ _19007_/Q _15098_/X _15171_/S vssd1 vssd1 vccd1 vccd1 _15172_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14472__S _14478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _12383_/A vssd1 vssd1 vccd1 vccd1 _17899_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12781__A _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11953__A1 _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14122_ _13940_/X _18576_/Q _14122_/S vssd1 vssd1 vccd1 vccd1 _14123_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11334_ _18462_/Q _19053_/Q _19215_/Q _18430_/Q _10572_/S _09542_/A vssd1 vssd1 vccd1
+ vccd1 _11335_/B sky130_fd_sc_hd__mux4_1
XFILLER_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18930_ _19379_/CLK _18930_/D vssd1 vssd1 vccd1 vccd1 _18930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14053_ _14109_/A vssd1 vssd1 vccd1 vccd1 _14122_/S sky130_fd_sc_hd__buf_6
XFILLER_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11265_ _18609_/Q _18944_/Q _11265_/S vssd1 vssd1 vccd1 vccd1 _11266_/B sky130_fd_sc_hd__mux2_1
XFILLER_107_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12902__A0 _19712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13004_ _13004_/A vssd1 vssd1 vccd1 vccd1 _13004_/X sky130_fd_sc_hd__clkbuf_2
X_10216_ _10216_/A vssd1 vssd1 vccd1 vccd1 _10216_/Y sky130_fd_sc_hd__inv_2
XFILLER_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18861_ _19085_/CLK _18861_/D vssd1 vssd1 vccd1 vccd1 _18861_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output150_A _16282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ _18610_/Q _18945_/Q _11196_/S vssd1 vssd1 vccd1 vccd1 _11196_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13816__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17812_ _17812_/A _17812_/B vssd1 vssd1 vccd1 vccd1 _17812_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17841__B1 _17840_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10147_ _19192_/Q _18806_/Q _19256_/Q _18375_/Q _09930_/S _09871_/X vssd1 vssd1 vccd1
+ vccd1 _10148_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18792_ _19306_/CLK _18792_/D vssd1 vssd1 vccd1 vccd1 _18792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14955_ _14955_/A vssd1 vssd1 vccd1 vccd1 _18923_/D sky130_fd_sc_hd__clkbuf_1
X_17743_ _17743_/A _17743_/B vssd1 vssd1 vccd1 vccd1 _17745_/B sky130_fd_sc_hd__nand2_1
XFILLER_130_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12666__C1 _12665_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10078_ _09760_/A _10065_/X _10076_/X _09833_/A _10077_/Y vssd1 vssd1 vccd1 vccd1
+ _12477_/B sky130_fd_sc_hd__o32a_4
XFILLER_35_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13117__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_1_0_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ _13922_/A vssd1 vssd1 vccd1 vccd1 _13919_/S sky130_fd_sc_hd__buf_2
XFILLER_63_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17674_ _17674_/A vssd1 vssd1 vccd1 vccd1 _17674_/Y sky130_fd_sc_hd__inv_2
X_14886_ _14886_/A vssd1 vssd1 vccd1 vccd1 _18890_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19413_ _19699_/CLK _19413_/D vssd1 vssd1 vccd1 vccd1 _19413_/Q sky130_fd_sc_hd__dfxtp_2
X_16625_ _16625_/A _16625_/B _16625_/C _16625_/D vssd1 vssd1 vccd1 vccd1 _16626_/D
+ sky130_fd_sc_hd__or4_1
X_13837_ _14519_/A vssd1 vssd1 vccd1 vccd1 _13837_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12956__A _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__S1 _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16556_ hold3/A _16559_/C _16546_/X vssd1 vssd1 vccd1 vccd1 _16556_/Y sky130_fd_sc_hd__a21oi_1
X_19344_ _19357_/CLK _19344_/D vssd1 vssd1 vccd1 vccd1 _19344_/Q sky130_fd_sc_hd__dfxtp_2
X_13768_ _12801_/X _18449_/Q _13776_/S vssd1 vssd1 vccd1 vccd1 _13769_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12433__A2 _12432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__B input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10444__A1 _10297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09330__A _11918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15507_ _15541_/A hold12/A vssd1 vssd1 vccd1 vccd1 _15507_/Y sky130_fd_sc_hd__nand2_1
X_12719_ _18107_/A _11260_/X _12735_/S vssd1 vssd1 vccd1 vccd1 _12719_/X sky130_fd_sc_hd__mux2_1
X_16487_ _16524_/A _16493_/C vssd1 vssd1 vccd1 vccd1 _16487_/Y sky130_fd_sc_hd__nor2_1
X_19275_ _19308_/CLK _19275_/D vssd1 vssd1 vccd1 vccd1 _19275_/Q sky130_fd_sc_hd__dfxtp_1
X_13699_ _12851_/X _18419_/Q _13703_/S vssd1 vssd1 vccd1 vccd1 _13700_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11071__S _11071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15438_ _19125_/Q _15067_/X _15444_/S vssd1 vssd1 vccd1 vccd1 _15439_/A sky130_fd_sc_hd__mux2_1
X_18226_ input51/X _18197_/X _18188_/X _18193_/X _18132_/A vssd1 vssd1 vccd1 vccd1
+ _18227_/B sky130_fd_sc_hd__a32o_1
XFILLER_50_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18157_ _18170_/A _18157_/B vssd1 vssd1 vccd1 vccd1 _18158_/A sky130_fd_sc_hd__and2_1
X_15369_ _15369_/A vssd1 vssd1 vccd1 vccd1 _19094_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14382__S _14384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17108_ _17108_/A _17108_/B vssd1 vssd1 vccd1 vccd1 _17109_/B sky130_fd_sc_hd__nor2_1
X_18088_ _14787_/B _18086_/X _18087_/X _18084_/X vssd1 vssd1 vccd1 vccd1 _19810_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17039_ _19668_/Q _15481_/X _17039_/S vssd1 vssd1 vccd1 vccd1 _17040_/A sky130_fd_sc_hd__mux2_1
X_09930_ _18633_/Q _18968_/Q _09930_/S vssd1 vssd1 vccd1 vccd1 _09930_/X sky130_fd_sc_hd__mux2_1
XFILLER_104_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10415__S _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11100__A _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09861_ _10197_/A vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__clkbuf_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09792_ _10439_/A vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__clkbuf_2
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10358__S1 _10238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17722__A _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12585__B _12606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09226_ _19857_/Q _19812_/Q vssd1 vssd1 vccd1 vccd1 _09226_/X sky130_fd_sc_hd__and2_1
XFILLER_21_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12188__A1 _09331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09157_ _09328_/A _18102_/A vssd1 vssd1 vccd1 vccd1 _09158_/A sky130_fd_sc_hd__nor2_1
XFILLER_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11935__A1 _11932_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09088_ _09146_/C _09180_/C _11585_/C vssd1 vssd1 vccd1 vccd1 _09207_/A sky130_fd_sc_hd__nor3_1
XFILLER_162_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11010__A _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ _18485_/Q _18980_/Q _11050_/S vssd1 vssd1 vccd1 vccd1 _11050_/X sky130_fd_sc_hd__mux2_1
XFILLER_115_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09987__S0 _09599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10001_ _09993_/X _09996_/X _09998_/X _10000_/X _09752_/A vssd1 vssd1 vccd1 vccd1
+ _10001_/X sky130_fd_sc_hd__a221o_4
XFILLER_77_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09415__A _09415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12648__C1 _12647_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10349__S1 _10436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14740_ _14553_/X _18826_/Q _14748_/S vssd1 vssd1 vccd1 vccd1 _14741_/A sky130_fd_sc_hd__mux2_1
XFILLER_57_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11952_ _17696_/A _11952_/B vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__xnor2_1
XFILLER_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ _10965_/A _10897_/Y _10900_/Y _11160_/A vssd1 vssd1 vccd1 vccd1 _10903_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14671_ _14671_/A vssd1 vssd1 vccd1 vccd1 _18795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10674__B2 _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11883_ _19337_/Q _11766_/X _12037_/A _11881_/X _16109_/A vssd1 vssd1 vccd1 vccd1
+ _11883_/X sky130_fd_sc_hd__o221a_1
XFILLER_44_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16410_ _19452_/Q _16411_/C _16409_/Y vssd1 vssd1 vccd1 vccd1 _19452_/D sky130_fd_sc_hd__o21a_1
XFILLER_83_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13622_ _13690_/S vssd1 vssd1 vccd1 vccd1 _13631_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_72_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17390_ _17390_/A vssd1 vssd1 vccd1 vccd1 _17390_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10834_ _18642_/Q vssd1 vssd1 vccd1 vccd1 _11020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16341_ _16341_/A _16341_/B _16341_/C vssd1 vssd1 vccd1 vccd1 _19430_/D sky130_fd_sc_hd__nor3_1
X_13553_ _13553_/A vssd1 vssd1 vccd1 vccd1 _18364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10765_ _09589_/A _10764_/X _10743_/A vssd1 vssd1 vccd1 vccd1 _10765_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19060_ _19319_/CLK _19060_/D vssd1 vssd1 vccd1 vccd1 _19060_/Q sky130_fd_sc_hd__dfxtp_1
X_12504_ _19472_/Q vssd1 vssd1 vccd1 vccd1 _16466_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16272_ _18150_/A _16272_/B vssd1 vssd1 vccd1 vccd1 _16273_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_190_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19311_/CLK sky130_fd_sc_hd__clkbuf_16
X_13484_ _13191_/X _18341_/Q _13492_/S vssd1 vssd1 vccd1 vccd1 _13485_/A sky130_fd_sc_hd__mux2_1
X_10696_ _18588_/Q _18859_/Q _19083_/Q _18827_/Q _10579_/X _10705_/A vssd1 vssd1 vccd1
+ vccd1 _10696_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15223_ _15223_/A vssd1 vssd1 vccd1 vccd1 _19029_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15298__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18011_ _18011_/A vssd1 vssd1 vccd1 vccd1 _19777_/D sky130_fd_sc_hd__clkbuf_1
X_12435_ _12435_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12435_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13400__A _13400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15154_ _18999_/Q _15073_/X _15156_/S vssd1 vssd1 vccd1 vccd1 _15155_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_0_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12366_ _19420_/Q vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_153_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14105_ _13915_/X _18568_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _14106_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11317_ _09368_/A _11307_/X _11316_/X _09471_/A _19720_/Q vssd1 vssd1 vccd1 vccd1
+ _11342_/A sky130_fd_sc_hd__a32o_2
XFILLER_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15085_ _15085_/A vssd1 vssd1 vccd1 vccd1 _18970_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14930__S _14930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ _17005_/A _12298_/C _19656_/Q vssd1 vssd1 vccd1 vccd1 _12297_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18913_ _19711_/CLK _18913_/D vssd1 vssd1 vccd1 vccd1 _18913_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output75_A _11988_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__S0 _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14036_ _14608_/A vssd1 vssd1 vccd1 vccd1 _14036_/X sky130_fd_sc_hd__clkbuf_2
X_11248_ _11248_/A _11248_/B vssd1 vssd1 vccd1 vccd1 _11248_/X sky130_fd_sc_hd__or2_1
XFILLER_79_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11855__A _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18844_ _19388_/CLK _18844_/D vssd1 vssd1 vccd1 vccd1 _18844_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11179_ _18388_/Q _18649_/Q _18548_/Q _18883_/Q _11243_/S _11177_/A vssd1 vssd1 vccd1
+ vccd1 _11180_/B sky130_fd_sc_hd__mux4_1
XFILLER_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18775_ _19326_/CLK _18775_/D vssd1 vssd1 vccd1 vccd1 _18775_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12103__A1 _19345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15987_ _15987_/A vssd1 vssd1 vccd1 vccd1 _19324_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15761__S _15765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17726_ _17726_/A _17726_/B _17726_/C vssd1 vssd1 vccd1 vccd1 _17726_/X sky130_fd_sc_hd__or3_1
XFILLER_76_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14938_ _18915_/Q vssd1 vssd1 vccd1 vccd1 _14939_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_75_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17042__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19711_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17657_ _17657_/A vssd1 vssd1 vccd1 vccd1 _17657_/Y sky130_fd_sc_hd__inv_2
X_14869_ _18883_/Q _13959_/X _14871_/S vssd1 vssd1 vccd1 vccd1 _14870_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16608_ _19516_/Q _16609_/C _16607_/Y vssd1 vssd1 vccd1 vccd1 _19516_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_78_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17588_ _17586_/X _17583_/Y _17587_/Y vssd1 vssd1 vccd1 vccd1 _17588_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19327_ _19375_/CLK _19327_/D vssd1 vssd1 vccd1 vccd1 _19327_/Q sky130_fd_sc_hd__dfxtp_1
X_16539_ _16540_/B _16540_/C _19494_/Q vssd1 vssd1 vccd1 vccd1 _16541_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10512__S1 _09710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_158_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19076_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09995__A _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19258_ _19384_/CLK _19258_/D vssd1 vssd1 vccd1 vccd1 _19258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17750__C1 _17831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18209_ _18213_/A _18209_/B vssd1 vssd1 vccd1 vccd1 _18210_/A sky130_fd_sc_hd__and2_1
XFILLER_163_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19189_ _19379_/CLK _19189_/D vssd1 vssd1 vccd1 vccd1 _19189_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10934__A _10934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11917__A1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15001__S _15013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13310__A _15086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10276__S0 _10274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09991__C1 _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09913_ _19195_/Q _18809_/Q _19259_/Q _18378_/Q _09904_/X _09905_/X vssd1 vssd1 vccd1
+ vccd1 _09914_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09969__S0 _10168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12342__A1 _19355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11765__A _11765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _09844_/A vssd1 vssd1 vccd1 vccd1 _09844_/X sky130_fd_sc_hd__buf_2
XFILLER_101_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09235__A _13400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09775_ _09785_/A vssd1 vssd1 vccd1 vccd1 _11389_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15671__S _15671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17033__A1 _13410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15595__A1 _12715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10503__S1 _09710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11005__A _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ _18591_/Q _18862_/Q _19086_/Q _18830_/Q _09415_/A _09443_/X vssd1 vssd1 vccd1
+ vccd1 _10550_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13358__B1 _12507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09209_ _17108_/A _11589_/B vssd1 vssd1 vccd1 vccd1 _17184_/C sky130_fd_sc_hd__nor2_1
XFILLER_136_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ _18625_/Q _18960_/Q _10481_/S vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__mux2_1
XFILLER_148_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_154_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ _12220_/A _17819_/B vssd1 vssd1 vccd1 vccd1 _12221_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15846__S _15848_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12151_ _19410_/Q _19411_/Q _12151_/C vssd1 vssd1 vccd1 vccd1 _12226_/C sky130_fd_sc_hd__and3_1
XANTENNA__10055__S _10055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10592__B1 _10074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ _11228_/A vssd1 vssd1 vccd1 vccd1 _11278_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12082_ _12020_/A _12465_/B _12081_/Y vssd1 vssd1 vccd1 vccd1 _17768_/B sky130_fd_sc_hd__a21o_2
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12333__A1 _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15910_ _15910_/A vssd1 vssd1 vccd1 vccd1 _19290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11033_ _11033_/A vssd1 vssd1 vccd1 vccd1 _11033_/X sky130_fd_sc_hd__clkbuf_4
X_16890_ _16890_/A vssd1 vssd1 vccd1 vccd1 _16915_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__14051__A _18089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12884__A2 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15841_ _15841_/A vssd1 vssd1 vccd1 vccd1 _19259_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10895__B2 _19714_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_60_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19319_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_92_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18560_ _19249_/CLK _18560_/D vssd1 vssd1 vccd1 vccd1 _18560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12984_ input32/X _12974_/A _12977_/A vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__a21o_1
X_15772_ _13602_/X _19229_/Q _15776_/S vssd1 vssd1 vccd1 vccd1 _15773_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17362_/X _17368_/A _17511_/S vssd1 vssd1 vccd1 vccd1 _17615_/B sky130_fd_sc_hd__mux2_1
XFILLER_18_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14723_ _14723_/A vssd1 vssd1 vccd1 vccd1 _18818_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11935_ _11934_/Y _11932_/Y _12100_/A vssd1 vssd1 vccd1 vccd1 _11935_/X sky130_fd_sc_hd__mux2_1
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18491_ _19006_/CLK _18491_/D vssd1 vssd1 vccd1 vccd1 _18491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10742__S1 _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17442_ _17439_/Y _17441_/Y _17500_/S vssd1 vssd1 vccd1 vccd1 _17653_/B sky130_fd_sc_hd__mux2_1
X_14654_ _14534_/X _18788_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14655_/A sky130_fd_sc_hd__mux2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _11879_/A _11793_/X _11861_/Y _11865_/X vssd1 vssd1 vccd1 vccd1 _16260_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_75_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19256_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_33_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _15089_/A vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_159_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10817_ _10817_/A vssd1 vssd1 vccd1 vccd1 _10817_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_60_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14585_ _14585_/A vssd1 vssd1 vccd1 vccd1 _14585_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17373_ _17371_/X _17372_/X _17497_/S vssd1 vssd1 vccd1 vccd1 _17552_/B sky130_fd_sc_hd__mux2_1
XANTENNA__18193__A _18234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11797_ _11795_/Y _11796_/Y _11858_/S vssd1 vssd1 vccd1 vccd1 _11797_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19112_ _19113_/CLK _19112_/D vssd1 vssd1 vccd1 vccd1 _19112_/Q sky130_fd_sc_hd__dfxtp_1
X_16324_ _19425_/Q _19424_/Q _19487_/Q _16324_/D vssd1 vssd1 vccd1 vccd1 _16333_/D
+ sky130_fd_sc_hd__and4_1
X_13536_ _18359_/Q _13535_/X _13545_/S vssd1 vssd1 vccd1 vccd1 _13537_/A sky130_fd_sc_hd__mux2_1
X_10748_ _09368_/A _10737_/X _10747_/Y _09471_/A _19717_/Q vssd1 vssd1 vccd1 vccd1
+ _10749_/B sky130_fd_sc_hd__a32o_2
XFILLER_146_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_146_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16255_ _16255_/A _16255_/B vssd1 vssd1 vccd1 vccd1 _16256_/A sky130_fd_sc_hd__or2_1
XFILLER_118_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19043_ _19205_/CLK _19043_/D vssd1 vssd1 vccd1 vccd1 _19043_/Q sky130_fd_sc_hd__dfxtp_1
X_13467_ _13467_/A vssd1 vssd1 vccd1 vccd1 _18333_/D sky130_fd_sc_hd__clkbuf_1
X_10679_ _19277_/Q _19115_/Q _18524_/Q _18294_/Q _10055_/S _10586_/X vssd1 vssd1 vccd1
+ vccd1 _10680_/B sky130_fd_sc_hd__mux4_1
XFILLER_173_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _19022_/Q _15044_/X _15206_/S vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12418_ _19422_/Q _12319_/X _12413_/X _12417_/X vssd1 vssd1 vccd1 vccd1 _12418_/X
+ sky130_fd_sc_hd__o22a_4
X_16186_ _16186_/A vssd1 vssd1 vccd1 vccd1 _19366_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11569__B _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13398_ _15565_/A vssd1 vssd1 vccd1 vccd1 _13398_/X sky130_fd_sc_hd__buf_2
XFILLER_154_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15137_ _18991_/Q _15047_/X _15145_/S vssd1 vssd1 vccd1 vccd1 _15138_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _12349_/A vssd1 vssd1 vccd1 vccd1 _17878_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_13_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19386_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_114_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15068_ _18965_/Q _15067_/X _15077_/S vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15510__A1 _15509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__A3 _12542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13276__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15057__A _15057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ _14019_/A vssd1 vssd1 vccd1 vccd1 _18534_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11585__A _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12875__A2 _12703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10430__S0 _10339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18827_ _19184_/CLK _18827_/D vssd1 vssd1 vccd1 vccd1 _18827_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold15_A hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19391_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09560_ _11022_/A vssd1 vssd1 vccd1 vccd1 _09561_/A sky130_fd_sc_hd__buf_2
XFILLER_95_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18758_ _19245_/CLK _18758_/D vssd1 vssd1 vccd1 vccd1 _18758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17015__A1 _15615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17709_ _17709_/A _17709_/B vssd1 vssd1 vccd1 vccd1 _17711_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09491_ _10721_/A vssd1 vssd1 vccd1 vccd1 _09644_/A sky130_fd_sc_hd__buf_2
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10929__A _10929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18689_ _19374_/CLK _18689_/D vssd1 vssd1 vccd1 vccd1 _18689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10733__S1 _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10648__B _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14835__S _14843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15520__A hold16/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15501__B2 _18258_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10603__S _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10877__A1 _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ _19294_/Q _19132_/Q _18541_/Q _18311_/Q _11385_/S _09785_/A vssd1 vssd1 vccd1
+ vccd1 _09827_/X sky130_fd_sc_hd__mux4_1
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10972__S1 _11266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09758_ _09758_/A vssd1 vssd1 vccd1 vccd1 _09758_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_101_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17006__A1 _12715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A1 _10680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _10414_/A vssd1 vssd1 vccd1 vccd1 _09690_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11716__A_N _11668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _18130_/A _18116_/A _12730_/C vssd1 vssd1 vccd1 vccd1 _11720_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17910__A _17910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _12372_/A _11736_/C _11649_/Y _12068_/A vssd1 vssd1 vccd1 vccd1 _11651_/X
+ sky130_fd_sc_hd__o31a_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10602_ _18621_/Q _18956_/Q _10602_/S vssd1 vssd1 vccd1 vccd1 _10602_/X sky130_fd_sc_hd__mux2_1
X_14370_ _14370_/A vssd1 vssd1 vccd1 vccd1 _18677_/D sky130_fd_sc_hd__clkbuf_1
X_11582_ _19860_/Q vssd1 vssd1 vccd1 vccd1 _18132_/A sky130_fd_sc_hd__buf_4
XFILLER_168_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13321_ _19166_/Q _13007_/X _12532_/X _19356_/Q _13320_/X vssd1 vssd1 vccd1 vccd1
+ _13321_/X sky130_fd_sc_hd__a221o_2
XFILLER_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10533_ _10535_/A _10532_/X _09821_/A vssd1 vssd1 vccd1 vccd1 _10533_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_7_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16040_ _16039_/A _16039_/C _12994_/A vssd1 vssd1 vccd1 vccd1 _16041_/B sky130_fd_sc_hd__o21ai_1
X_13252_ _13251_/X _18307_/Q _13252_/S vssd1 vssd1 vccd1 vccd1 _13253_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10464_ _18465_/Q _19056_/Q _19218_/Q _18433_/Q _10499_/S _10229_/A vssd1 vssd1 vccd1
+ vccd1 _10464_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12203_ _19349_/Q _11733_/X _12037_/X _12202_/X _12102_/X vssd1 vssd1 vccd1 vccd1
+ _12203_/X sky130_fd_sc_hd__o221a_1
XFILLER_89_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ _19444_/Q _12515_/X _13182_/X vssd1 vssd1 vccd1 vccd1 _13183_/X sky130_fd_sc_hd__o21a_1
X_10395_ _19284_/Q _19122_/Q _18531_/Q _18301_/Q _10260_/X _10436_/A vssd1 vssd1 vccd1
+ vccd1 _10395_/X sky130_fd_sc_hd__mux4_1
XANTENNA_clkbuf_leaf_26_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ _12134_/A vssd1 vssd1 vccd1 vccd1 _12134_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_124_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17991_ _17991_/A vssd1 vssd1 vccd1 vccd1 _19768_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10580__A3 _18830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11609__S _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19730_ _19734_/CLK _19730_/D vssd1 vssd1 vccd1 vccd1 _19730_/Q sky130_fd_sc_hd__dfxtp_4
X_16942_ _13404_/X _16957_/B _16941_/X _16833_/A vssd1 vssd1 vccd1 vccd1 _19631_/D
+ sky130_fd_sc_hd__a211o_1
X_12065_ _12066_/B _12065_/B vssd1 vssd1 vccd1 vccd1 _12067_/B sky130_fd_sc_hd__nor2_1
XFILLER_145_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11016_ _09366_/A _11001_/X _11015_/X _09469_/A _19712_/Q vssd1 vssd1 vccd1 vccd1
+ _11016_/X sky130_fd_sc_hd__a32o_2
XFILLER_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19661_ _19687_/CLK _19661_/D vssd1 vssd1 vccd1 vccd1 _19661_/Q sky130_fd_sc_hd__dfxtp_1
X_16873_ _16881_/A _16873_/B _16873_/C vssd1 vssd1 vccd1 vccd1 _19602_/D sky130_fd_sc_hd__nor3_1
XFILLER_78_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18188__A _18188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18612_ _19364_/CLK _18612_/D vssd1 vssd1 vccd1 vccd1 _18612_/Q sky130_fd_sc_hd__dfxtp_1
X_15824_ _13573_/X _19252_/Q _15826_/S vssd1 vssd1 vccd1 vccd1 _15825_/A sky130_fd_sc_hd__mux2_1
X_19592_ _19594_/CLK _19592_/D vssd1 vssd1 vccd1 vccd1 _19592_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16200__S _16202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18543_ _19388_/CLK _18543_/D vssd1 vssd1 vccd1 vccd1 _18543_/Q sky130_fd_sc_hd__dfxtp_1
X_15755_ _15755_/A vssd1 vssd1 vccd1 vccd1 _19221_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12967_ _13247_/S vssd1 vssd1 vccd1 vccd1 _13381_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15559__A1 _12577_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14706_ _14706_/A vssd1 vssd1 vccd1 vccd1 _18811_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17820__A _17917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ _18146_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _12159_/B sky130_fd_sc_hd__nand2_1
XFILLER_73_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18474_ _19291_/CLK _18474_/D vssd1 vssd1 vccd1 vccd1 _18474_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09365__B1_N _09468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15686_ _15686_/A vssd1 vssd1 vccd1 vccd1 _19190_/D sky130_fd_sc_hd__clkbuf_1
X_12898_ _19557_/Q _12701_/X _12897_/X _12707_/X vssd1 vssd1 vccd1 vccd1 _12898_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _17333_/X _17384_/X _17386_/X _17424_/Y vssd1 vssd1 vccd1 vccd1 _17425_/X
+ sky130_fd_sc_hd__a211o_1
X_14637_ _16301_/A vssd1 vssd1 vccd1 vccd1 _16282_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_11849_ _11849_/A vssd1 vssd1 vccd1 vccd1 _11854_/A sky130_fd_sc_hd__clkinv_2
XFILLER_61_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17356_ _17223_/X _17204_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17356_/X sky130_fd_sc_hd__mux2_1
X_14568_ _14568_/A vssd1 vssd1 vccd1 vccd1 _18761_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10399__A3 _10397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16307_ _19422_/Q _12440_/A _12413_/X _12417_/X _12556_/X vssd1 vssd1 vccd1 vccd1
+ _19422_/D sky130_fd_sc_hd__o221a_1
X_13519_ _15003_/A vssd1 vssd1 vccd1 vccd1 _13519_/X sky130_fd_sc_hd__clkbuf_2
X_14499_ _14499_/A vssd1 vssd1 vccd1 vccd1 _18733_/D sky130_fd_sc_hd__clkbuf_1
X_17287_ _17285_/X _17286_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17287_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17720__A2 _17652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19026_ _19091_/CLK _19026_/D vssd1 vssd1 vccd1 vccd1 _19026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16238_ _16238_/A vssd1 vssd1 vccd1 vccd1 _19390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16169_ _16169_/A _16169_/B vssd1 vssd1 vccd1 vccd1 _16226_/A sky130_fd_sc_hd__nand2_2
XANTENNA__16171__A _16239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19859_ _19866_/CLK _19859_/D vssd1 vssd1 vccd1 vccd1 _19859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13734__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09612_ _18479_/Q _19070_/Q _19232_/Q _18447_/Q _09599_/X _09419_/A vssd1 vssd1 vccd1
+ vccd1 _09612_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10954__S1 _09416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_clock_A clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09513__A _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ _09543_/A vssd1 vssd1 vccd1 vccd1 _09768_/A sky130_fd_sc_hd__buf_2
XANTENNA__10659__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09474_ _09474_/A _09474_/B vssd1 vssd1 vccd1 vccd1 _09474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12593__B _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11131__S1 _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10394__A _10394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11992__C1 _16109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10890__S0 _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15396__S _15400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12813__S _12887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17432__C_N _17190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17475__A1 _11639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10180_ _10181_/A _12471_/B vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__and2_1
XANTENNA__14289__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14289__B2 _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10945__S1 _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ _14550_/A vssd1 vssd1 vccd1 vccd1 _13870_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12821_ _19425_/Q _12700_/X _12820_/X vssd1 vssd1 vccd1 vccd1 _12821_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09423__A _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10569__A _10689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17640__A _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15540_ hold13/A _15540_/B vssd1 vssd1 vccd1 vccd1 _15540_/X sky130_fd_sc_hd__or2_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ _12773_/A vssd1 vssd1 vccd1 vccd1 _12752_/X sky130_fd_sc_hd__buf_2
XANTENNA__10078__A2 _10065_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11703_ _11804_/B _11703_/B _11703_/C vssd1 vssd1 vccd1 vccd1 _11703_/X sky130_fd_sc_hd__and3_1
X_15471_ _11120_/Y _12071_/X _13419_/B vssd1 vssd1 vccd1 vccd1 _15471_/Y sky130_fd_sc_hd__o21ai_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _19575_/Q _12518_/X _12682_/X _12538_/X vssd1 vssd1 vccd1 vccd1 _12683_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ _13909_/X _18699_/Q _14428_/S vssd1 vssd1 vccd1 vccd1 _14423_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11027__A1 _19109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17210_ _17440_/B _17208_/X _17501_/S vssd1 vssd1 vccd1 vccd1 _17210_/X sky130_fd_sc_hd__mux2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11634_/A _17575_/S vssd1 vssd1 vccd1 vccd1 _11681_/A sky130_fd_sc_hd__xnor2_2
XFILLER_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18190_ _18190_/A _18190_/B vssd1 vssd1 vccd1 vccd1 _18191_/A sky130_fd_sc_hd__and2_1
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _14353_/A vssd1 vssd1 vccd1 vccd1 _18669_/D sky130_fd_sc_hd__clkbuf_1
X_17141_ _18099_/A _17130_/B _17140_/X _19700_/Q vssd1 vssd1 vccd1 vccd1 _17142_/B
+ sky130_fd_sc_hd__a22o_1
X_11565_ _11565_/A vssd1 vssd1 vccd1 vccd1 _17105_/A sky130_fd_sc_hd__buf_2
XFILLER_129_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _19547_/Q _12952_/X _12953_/X _19515_/Q _13303_/X vssd1 vssd1 vccd1 vccd1
+ _13304_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17072_ _19683_/Q _15568_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17073_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10516_ _09727_/A _10509_/X _10511_/X _10515_/X _09753_/A vssd1 vssd1 vccd1 vccd1
+ _10516_/X sky130_fd_sc_hd__a311o_4
X_14284_ _14290_/A _18218_/B vssd1 vssd1 vccd1 vccd1 _14285_/A sky130_fd_sc_hd__and2_2
XANTENNA__10881__S0 _10878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16910__B1 _16344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11496_ _12322_/A vssd1 vssd1 vccd1 vccd1 _19137_/D sky130_fd_sc_hd__inv_2
XFILLER_171_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13235_ _19730_/Q _12687_/B _13306_/A vssd1 vssd1 vccd1 vccd1 _13235_/X sky130_fd_sc_hd__mux2_1
X_16023_ _16028_/B _16023_/B vssd1 vssd1 vccd1 vccd1 _16023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_155_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10447_ _11445_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _11446_/A sky130_fd_sc_hd__or2_1
XFILLER_152_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10002__A2 _09991_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11847__B _17198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13166_ _13166_/A vssd1 vssd1 vccd1 vccd1 _13166_/X sky130_fd_sc_hd__clkbuf_2
X_10378_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_152_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12117_ _12117_/A _17219_/A vssd1 vssd1 vccd1 vccd1 _12118_/B sky130_fd_sc_hd__or2_1
X_13097_ _19679_/Q _12817_/X _12680_/A _19646_/Q vssd1 vssd1 vccd1 vccd1 _13097_/X
+ sky130_fd_sc_hd__a22o_1
X_17974_ _17974_/A vssd1 vssd1 vccd1 vccd1 _19760_/D sky130_fd_sc_hd__clkbuf_1
X_19713_ _19740_/CLK _19713_/D vssd1 vssd1 vccd1 vccd1 _19713_/Q sky130_fd_sc_hd__dfxtp_4
X_16925_ input67/X _16929_/B vssd1 vssd1 vccd1 vccd1 _16925_/X sky130_fd_sc_hd__or2_1
X_12048_ _12020_/X _12464_/B _12047_/Y vssd1 vssd1 vccd1 vccd1 _12110_/A sky130_fd_sc_hd__a21o_1
XFILLER_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17026__S _17026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11863__A _16963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19644_ _19645_/CLK _19644_/D vssd1 vssd1 vccd1 vccd1 _19644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16856_ _16881_/A _16856_/B _16856_/C vssd1 vssd1 vccd1 vccd1 _19596_/D sky130_fd_sc_hd__nor3_1
XFILLER_77_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09333__A _09351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15807_ _13547_/X _19244_/Q _15815_/S vssd1 vssd1 vccd1 vccd1 _15808_/A sky130_fd_sc_hd__mux2_1
XFILLER_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19575_ _19668_/CLK _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16787_ _16790_/B _16790_/C _19570_/Q vssd1 vssd1 vccd1 vccd1 _16789_/B sky130_fd_sc_hd__a21oi_1
XFILLER_93_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13999_ _18528_/Q _13997_/X _14011_/S vssd1 vssd1 vccd1 vccd1 _14000_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11074__S _11074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18526_ _19373_/CLK _18526_/D vssd1 vssd1 vccd1 vccd1 _18526_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15738_ _15738_/A vssd1 vssd1 vccd1 vccd1 _19213_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18457_ _19306_/CLK _18457_/D vssd1 vssd1 vccd1 vccd1 _18457_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12694__A _18142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15669_ _14563_/X _19183_/Q _15671_/S vssd1 vssd1 vccd1 vccd1 _15670_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15070__A _15070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17408_ _17408_/A vssd1 vssd1 vccd1 vccd1 _17800_/A sky130_fd_sc_hd__clkbuf_2
X_09190_ _19850_/Q vssd1 vssd1 vccd1 vccd1 _09341_/A sky130_fd_sc_hd__clkbuf_2
X_18388_ _19205_/CLK _18388_/D vssd1 vssd1 vccd1 vccd1 _18388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11113__S1 _11075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17339_ _17266_/A _17231_/X _17338_/X vssd1 vssd1 vccd1 vccd1 _17340_/A sky130_fd_sc_hd__a21oi_1
XFILLER_140_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__A1 _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17709__B _17709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19009_ _19740_/CLK _19009_/D vssd1 vssd1 vccd1 vccd1 _19009_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18103__C1 _18097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10624__S0 _10055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15468__A0 _09315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13464__S _13470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10701__B1 _09760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09526_ _18638_/Q _18973_/Q _09776_/A vssd1 vssd1 vccd1 vccd1 _09527_/B sky130_fd_sc_hd__mux2_1
XFILLER_25_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09457_ _10046_/A vssd1 vssd1 vccd1 vccd1 _10236_/A sky130_fd_sc_hd__clkbuf_2
XPHY_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09389__S _09981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ _10030_/S vssd1 vssd1 vccd1 vccd1 _09981_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11350_ _11448_/A _11451_/A _11448_/C _10495_/A _11349_/X vssd1 vssd1 vccd1 vccd1
+ _11443_/C sky130_fd_sc_hd__a311o_1
XFILLER_153_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10863__S0 _10862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _09762_/A _10284_/X _10299_/X _09835_/A _10300_/Y vssd1 vssd1 vccd1 vccd1
+ _12468_/B sky130_fd_sc_hd__o32a_4
X_11281_ _11274_/Y _11276_/Y _11278_/Y _11280_/Y _10929_/A vssd1 vssd1 vccd1 vccd1
+ _11281_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13020_ _13033_/A _13020_/B _13031_/B vssd1 vssd1 vccd1 vccd1 _13020_/X sky130_fd_sc_hd__or3_1
X_10232_ _18629_/Q _18964_/Q _10367_/S vssd1 vssd1 vccd1 vccd1 _10232_/X sky130_fd_sc_hd__mux2_1
XFILLER_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09418__A _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10615__S0 _10763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11193__B1 _12445_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10163_ _19320_/Q _18732_/Q _18769_/Q _18343_/Q _09782_/A _09956_/A vssd1 vssd1 vccd1
+ vccd1 _10163_/X sky130_fd_sc_hd__mux4_1
XFILLER_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16120__A1 _19350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09137__B _19863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__S1 _10090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input37_A io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14971_ _14971_/A vssd1 vssd1 vccd1 vccd1 _18931_/D sky130_fd_sc_hd__clkbuf_1
X_10094_ _18504_/Q _18999_/Q _10094_/S vssd1 vssd1 vccd1 vccd1 _10094_/X sky130_fd_sc_hd__mux2_1
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16710_ _16715_/C _16715_/D _16709_/Y vssd1 vssd1 vccd1 vccd1 _19546_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10918__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11040__S0 _11265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13922_ _13922_/A vssd1 vssd1 vccd1 vccd1 _13935_/S sky130_fd_sc_hd__buf_4
XFILLER_47_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17690_ _19718_/Q _17688_/X _17873_/S vssd1 vssd1 vccd1 vccd1 _17691_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17620__A1 _11824_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ _16650_/B _16650_/C _14290_/A vssd1 vssd1 vccd1 vccd1 _16642_/B sky130_fd_sc_hd__o21ai_1
XFILLER_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13853_ _13853_/A vssd1 vssd1 vccd1 vccd1 _18484_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ _19701_/Q _16000_/B vssd1 vssd1 vccd1 vccd1 _13435_/B sky130_fd_sc_hd__and2_1
X_19360_ _19361_/CLK _19360_/D vssd1 vssd1 vccd1 vccd1 _19360_/Q sky130_fd_sc_hd__dfxtp_1
X_16572_ _19505_/Q _16575_/C _16546_/X vssd1 vssd1 vccd1 vccd1 _16572_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13784_ _13784_/A vssd1 vssd1 vccd1 vccd1 _18456_/D sky130_fd_sc_hd__clkbuf_1
X_10996_ _18582_/Q _18853_/Q _19077_/Q _18821_/Q _11196_/S _10990_/A vssd1 vssd1 vccd1
+ vccd1 _10996_/X sky130_fd_sc_hd__mux4_1
XFILLER_90_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09310__B1 _09309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18311_ _19326_/CLK _18311_/D vssd1 vssd1 vccd1 vccd1 _18311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15523_ _15601_/A vssd1 vssd1 vccd1 vccd1 _15543_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12735_ _18116_/A _11070_/X _12735_/S vssd1 vssd1 vccd1 vccd1 _12735_/X sky130_fd_sc_hd__mux2_1
X_19291_ _19291_/CLK _19291_/D vssd1 vssd1 vccd1 vccd1 _19291_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18242_ _18248_/A _18242_/B vssd1 vssd1 vccd1 vccd1 _18243_/A sky130_fd_sc_hd__and2_1
XFILLER_31_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _19600_/Q _12633_/X _12634_/X _19468_/Q _12665_/X vssd1 vssd1 vccd1 vccd1
+ _12667_/B sky130_fd_sc_hd__a221o_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _15454_/A vssd1 vssd1 vccd1 vccd1 _19132_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12748__A1 hold16/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ _12184_/A vssd1 vssd1 vccd1 vccd1 _13411_/A sky130_fd_sc_hd__clkbuf_2
X_14405_ _14405_/A vssd1 vssd1 vccd1 vccd1 _18691_/D sky130_fd_sc_hd__clkbuf_1
X_18173_ _18233_/A vssd1 vssd1 vccd1 vccd1 _18190_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_156_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12597_ _18234_/A vssd1 vssd1 vccd1 vccd1 _16929_/B sky130_fd_sc_hd__buf_2
XFILLER_129_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15385_ _19102_/Q _15095_/X _15387_/S vssd1 vssd1 vccd1 vccd1 _15386_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09613__A1 _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16714__A _16714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17124_ _17105_/X _17124_/B vssd1 vssd1 vccd1 vccd1 _17176_/B sky130_fd_sc_hd__and2b_1
X_14336_ _14336_/A vssd1 vssd1 vccd1 vccd1 _18661_/D sky130_fd_sc_hd__clkbuf_1
X_11548_ _12322_/A _12322_/B vssd1 vssd1 vccd1 vccd1 _11738_/A sky130_fd_sc_hd__nand2_1
XFILLER_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13549__S _13561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17055_ _19675_/Q _12651_/X _17061_/S vssd1 vssd1 vccd1 vccd1 _17056_/A sky130_fd_sc_hd__mux2_1
X_14267_ _14267_/A vssd1 vssd1 vccd1 vccd1 _18639_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10762__A _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11479_ _10082_/X _11428_/A _11428_/B vssd1 vssd1 vccd1 vccd1 _11479_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_109_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13218_ _19160_/Q _13179_/X _12958_/X _19350_/Q _13217_/X vssd1 vssd1 vccd1 vccd1
+ _13218_/X sky130_fd_sc_hd__a221o_2
X_16006_ _15998_/A _19136_/Q vssd1 vssd1 vccd1 vccd1 _16011_/C sky130_fd_sc_hd__nand2b_1
XANTENNA__10606__S0 _10763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14198_ _15317_/A _15101_/A vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__nor2_2
XFILLER_98_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12920__A1 _15493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ _13148_/X _18301_/Q _13172_/S vssd1 vssd1 vccd1 vccd1 _13150_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16111__A1 _12233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _16069_/A _19785_/Q _17957_/S vssd1 vssd1 vccd1 vccd1 _17958_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16908_ _16915_/A _16912_/C vssd1 vssd1 vccd1 vccd1 _16908_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18079__C _18099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17888_ _17406_/X _17889_/B _17887_/X _17537_/X vssd1 vssd1 vccd1 vccd1 _17888_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19627_ _19828_/CLK _19627_/D vssd1 vssd1 vccd1 vccd1 _19627_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_66_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16839_ _16839_/A vssd1 vssd1 vccd1 vccd1 _16845_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19558_ _19564_/CLK _19558_/D vssd1 vssd1 vccd1 vccd1 _19558_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12436__B1 _12230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_148_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09311_ _19707_/Q vssd1 vssd1 vccd1 vccd1 _09311_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__12987__A1 _19147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11334__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18509_ _19326_/CLK _18509_/D vssd1 vssd1 vccd1 vccd1 _18509_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12987__B2 _19337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19489_ _19619_/CLK _19489_/D vssd1 vssd1 vccd1 vccd1 _19489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10937__A _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15004__S _15013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ _12672_/A vssd1 vssd1 vccd1 vccd1 _14275_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_167_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09173_ _09134_/C _11646_/C _09327_/A vssd1 vssd1 vccd1 vccd1 _17753_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__14843__S _14843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17752__B_N _12089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09604__A1 _09434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11768__A _19397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09238__A _11560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10517__A3 _10516_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15674__S _15682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11714__A2 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17455__A _17504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17190__A _17190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10850_ _11263_/S vssd1 vssd1 vccd1 vccd1 _10962_/S sky130_fd_sc_hd__buf_4
XFILLER_71_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11325__S1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12978__A1 input31/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09557_/A _09509_/B vssd1 vssd1 vccd1 vccd1 _09509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_169_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10781_ _10639_/X _10780_/X _09484_/A vssd1 vssd1 vccd1 vccd1 _10781_/Y sky130_fd_sc_hd__o21ai_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12520_ _13009_/A vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_9_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11470__C_N _11469_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ _18100_/A _12475_/A _11542_/A vssd1 vssd1 vccd1 vccd1 _12462_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14753__S _14759_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _11402_/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11402_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15170_ _15170_/A vssd1 vssd1 vccd1 vccd1 _19006_/D sky130_fd_sc_hd__clkbuf_1
X_12382_ _19800_/Q _11418_/A _12423_/S vssd1 vssd1 vccd1 vccd1 _12383_/A sky130_fd_sc_hd__mux2_8
XFILLER_165_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14121_ _14121_/A vssd1 vssd1 vccd1 vccd1 _18575_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11333_ _10639_/X _11332_/X _09630_/X vssd1 vssd1 vccd1 vccd1 _11333_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10610__C1 _09374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11678__A _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14054__A _14122_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14352__A0 _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ _14299_/A _16169_/A vssd1 vssd1 vccd1 vccd1 _14109_/A sky130_fd_sc_hd__nand2_2
X_11264_ _11264_/A vssd1 vssd1 vccd1 vccd1 _11264_/Y sky130_fd_sc_hd__inv_2
XFILLER_153_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13003_ _19466_/Q vssd1 vssd1 vccd1 vccd1 _16450_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12902__A1 _15485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _18502_/Q _18997_/Q _10215_/S vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__mux2_1
X_18860_ _19374_/CLK _18860_/D vssd1 vssd1 vccd1 vccd1 _18860_/Q sky130_fd_sc_hd__dfxtp_1
X_11195_ _11195_/A _11195_/B vssd1 vssd1 vccd1 vccd1 _11195_/X sky130_fd_sc_hd__or2_1
XANTENNA__11261__S0 _10962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17811_ _17809_/X _17812_/B _17844_/S vssd1 vssd1 vccd1 vccd1 _17811_/X sky130_fd_sc_hd__mux2_1
XFILLER_122_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10146_ _09730_/A _10141_/X _10143_/X _10145_/X _09859_/A vssd1 vssd1 vccd1 vccd1
+ _10146_/X sky130_fd_sc_hd__a221o_1
XANTENNA__17841__A1 _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18791_ _19239_/CLK _18791_/D vssd1 vssd1 vccd1 vccd1 _18791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15852__A0 _13614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11013__S0 _11011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17742_ _17743_/A _17743_/B _17842_/S vssd1 vssd1 vccd1 vccd1 _17742_/X sky130_fd_sc_hd__mux2_1
XFILLER_153_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14954_ _18923_/Q vssd1 vssd1 vccd1 vccd1 _14955_/A sky130_fd_sc_hd__clkbuf_1
X_10077_ _19734_/Q vssd1 vssd1 vccd1 vccd1 _10077_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13905_ _14585_/A vssd1 vssd1 vccd1 vccd1 _13905_/X sky130_fd_sc_hd__buf_2
X_17673_ _17673_/A vssd1 vssd1 vccd1 vccd1 _17673_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_75_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14885_ _18890_/Q _13981_/X _14893_/S vssd1 vssd1 vccd1 vccd1 _14886_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14928__S _14930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19412_ _19699_/CLK _19412_/D vssd1 vssd1 vccd1 vccd1 _19412_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16624_ _16624_/A _16624_/B vssd1 vssd1 vccd1 vccd1 _16625_/D sky130_fd_sc_hd__or2_1
X_13836_ _13836_/A vssd1 vssd1 vccd1 vccd1 _18480_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19343_ _19349_/CLK _19343_/D vssd1 vssd1 vccd1 vccd1 _19343_/Q sky130_fd_sc_hd__dfxtp_2
X_16555_ _19498_/Q _16552_/C _16554_/Y vssd1 vssd1 vccd1 vccd1 _19498_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ _13835_/S vssd1 vssd1 vccd1 vccd1 _13776_/S sky130_fd_sc_hd__clkbuf_4
X_10979_ _10981_/A _10978_/X _09561_/A vssd1 vssd1 vccd1 vccd1 _10979_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_31_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15506_ _15629_/A vssd1 vssd1 vccd1 vccd1 _15541_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12718_ _12674_/X _12696_/X _12717_/X _12694_/X vssd1 vssd1 vccd1 vccd1 _19585_/D
+ sky130_fd_sc_hd__o22a_1
X_19274_ _19308_/CLK _19274_/D vssd1 vssd1 vccd1 vccd1 _19274_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16486_ _16486_/A vssd1 vssd1 vccd1 vccd1 _16493_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13698_ _13698_/A vssd1 vssd1 vccd1 vccd1 _18418_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15759__S _15765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18225_ _18225_/A vssd1 vssd1 vccd1 vccd1 _19859_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15437_ _15437_/A vssd1 vssd1 vccd1 vccd1 _19124_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12649_ _18262_/Q _12649_/B vssd1 vssd1 vccd1 vccd1 _12649_/X sky130_fd_sc_hd__or2_1
XFILLER_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18156_ input56/X _18155_/X _18066_/S _12657_/X _18075_/A vssd1 vssd1 vccd1 vccd1
+ _18157_/B sky130_fd_sc_hd__a32o_1
XFILLER_172_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15368_ _19094_/Q _15070_/X _15372_/S vssd1 vssd1 vccd1 vccd1 _15369_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ _17107_/A vssd1 vssd1 vccd1 vccd1 _17177_/B sky130_fd_sc_hd__clkinv_2
X_14319_ _13867_/X _18654_/Q _14321_/S vssd1 vssd1 vccd1 vccd1 _14320_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18087_ _18087_/A _18087_/B vssd1 vssd1 vccd1 vccd1 _18087_/X sky130_fd_sc_hd__or2_1
X_15299_ _15299_/A vssd1 vssd1 vccd1 vccd1 _19063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17038_ _17038_/A vssd1 vssd1 vccd1 vccd1 _19667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_74_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ _10200_/A vssd1 vssd1 vccd1 vccd1 _10197_/A sky130_fd_sc_hd__buf_2
XFILLER_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _10485_/A vssd1 vssd1 vccd1 vccd1 _10439_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15507__B hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _19006_/CLK _18989_/D vssd1 vssd1 vccd1 vccd1 _18989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17722__B _17722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15523__A _15601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13082__A0 _19721_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10667__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09225_ _11619_/A _19812_/Q vssd1 vssd1 vccd1 vccd1 _09225_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15669__S _15671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10986__A3 _10984_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16354__A _16868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09156_ _09174_/B vssd1 vssd1 vccd1 vccd1 _18102_/A sky130_fd_sc_hd__inv_2
XANTENNA__10818__S0 _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17520__A0 _19710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09087_ _09167_/A vssd1 vssd1 vccd1 vccd1 _11585_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_163_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09987__S1 _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16087__A0 _12577_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14602__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10000_ _09993_/A _09999_/X _09737_/A vssd1 vssd1 vccd1 vccd1 _10000_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09989_ _09989_/A vssd1 vssd1 vccd1 vccd1 _09989_/X sky130_fd_sc_hd__buf_4
XFILLER_130_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10341__S _10341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11951_ _12111_/A _12025_/B vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__nand2_1
XFILLER_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14748__S _14748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10902_ _11262_/A vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__buf_2
X_11882_ _12654_/B vssd1 vssd1 vccd1 vccd1 _16109_/A sky130_fd_sc_hd__clkbuf_2
X_14670_ _14557_/X _18795_/Q _14676_/S vssd1 vssd1 vccd1 vccd1 _14671_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09431__A _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11680__B _17237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10833_ _09368_/A _10821_/X _10832_/X _09471_/A _19715_/Q vssd1 vssd1 vccd1 vccd1
+ _11291_/A sky130_fd_sc_hd__a32o_2
X_13621_ _13677_/A vssd1 vssd1 vccd1 vccd1 _13690_/S sky130_fd_sc_hd__buf_6
XFILLER_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__A _10586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11172__S _11172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16340_ _19430_/Q _16340_/B _16340_/C vssd1 vssd1 vccd1 vccd1 _16341_/C sky130_fd_sc_hd__and3_1
XFILLER_25_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13552_ _18364_/Q _13551_/X _13561_/S vssd1 vssd1 vccd1 vccd1 _13553_/A sky130_fd_sc_hd__mux2_1
X_10764_ _18490_/Q _18985_/Q _10764_/S vssd1 vssd1 vccd1 vccd1 _10764_/X sky130_fd_sc_hd__mux2_1
XFILLER_34_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ _12503_/A vssd1 vssd1 vccd1 vccd1 _12503_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10831__C1 _09448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16271_ _16890_/A vssd1 vssd1 vccd1 vccd1 _18150_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14483__S _14489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13483_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13492_/S sky130_fd_sc_hd__buf_4
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10695_ _18396_/Q _18657_/Q _18556_/Q _18891_/Q _10576_/X _10577_/X vssd1 vssd1 vccd1
+ vccd1 _10695_/X sky130_fd_sc_hd__mux4_1
XFILLER_173_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18010_ _19777_/Q _11826_/A _18016_/S vssd1 vssd1 vccd1 vccd1 _18011_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15222_ _19029_/Q _15067_/X _15228_/S vssd1 vssd1 vccd1 vccd1 _15223_/A sky130_fd_sc_hd__mux2_1
X_12434_ _19423_/Q _12434_/B vssd1 vssd1 vccd1 vccd1 _12435_/B sky130_fd_sc_hd__xnor2_1
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ _15153_/A vssd1 vssd1 vccd1 vccd1 _18998_/D sky130_fd_sc_hd__clkbuf_1
X_12365_ _12365_/A vssd1 vssd1 vccd1 vccd1 _12369_/B sky130_fd_sc_hd__buf_4
XFILLER_154_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14104_ _14104_/A vssd1 vssd1 vccd1 vccd1 _18567_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11316_ _11309_/X _11311_/X _11313_/X _11315_/X _09614_/X vssd1 vssd1 vccd1 vccd1
+ _11316_/X sky130_fd_sc_hd__a221o_4
X_15084_ _18970_/Q _15083_/X _15093_/S vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12296_ _19353_/Q _11733_/X _11734_/X _12295_/X _12102_/X vssd1 vssd1 vccd1 vccd1
+ _12296_/X sky130_fd_sc_hd__o221a_1
XFILLER_99_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18912_ _19361_/CLK _18912_/D vssd1 vssd1 vccd1 vccd1 _18912_/Q sky130_fd_sc_hd__dfxtp_1
X_14035_ _14035_/A vssd1 vssd1 vccd1 vccd1 _18539_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13827__S _13831_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11247_ _18385_/Q _18646_/Q _18545_/Q _18880_/Q _11123_/A _10933_/A vssd1 vssd1 vccd1
+ vccd1 _11248_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10037__S1 _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18843_ _19390_/CLK _18843_/D vssd1 vssd1 vccd1 vccd1 _18843_/Q sky130_fd_sc_hd__dfxtp_1
X_11178_ _18580_/Q _18851_/Q _19075_/Q _18819_/Q _11127_/S _11177_/X vssd1 vssd1 vccd1
+ vccd1 _11178_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14628__A1 input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14628__B2 _09194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10129_ _10129_/A _10129_/B vssd1 vssd1 vccd1 vccd1 _10129_/Y sky130_fd_sc_hd__nor2_1
X_18774_ _19261_/CLK _18774_/D vssd1 vssd1 vccd1 vccd1 _18774_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15986_ _13599_/X _19324_/Q _15992_/S vssd1 vssd1 vccd1 vccd1 _15987_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _17724_/A _17726_/C _17724_/Y vssd1 vssd1 vccd1 vccd1 _17725_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14937_ _14937_/A vssd1 vssd1 vccd1 vccd1 _18914_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17656_ _17625_/S _17653_/X _17654_/Y _17655_/X vssd1 vssd1 vccd1 vccd1 _17656_/X
+ sky130_fd_sc_hd__a31o_1
X_14868_ _14868_/A vssd1 vssd1 vccd1 vccd1 _18882_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16607_ _16610_/A _16607_/B vssd1 vssd1 vccd1 vccd1 _16607_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13819_ _13819_/A vssd1 vssd1 vccd1 vccd1 _18472_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17587_ _17587_/A _17587_/B vssd1 vssd1 vccd1 vccd1 _17587_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14799_ _18852_/Q _13962_/X _14799_/S vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19326_ _19326_/CLK _19326_/D vssd1 vssd1 vccd1 vccd1 _19326_/Q sky130_fd_sc_hd__dfxtp_1
X_16538_ _16540_/B _16540_/C _16537_/Y vssd1 vssd1 vccd1 vccd1 _19493_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19257_ _19383_/CLK _19257_/D vssd1 vssd1 vccd1 vccd1 _19257_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16469_ _16469_/A vssd1 vssd1 vccd1 vccd1 _16474_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14393__S _14395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18208_ _18208_/A vssd1 vssd1 vccd1 vccd1 _19851_/D sky130_fd_sc_hd__clkbuf_1
X_19188_ _19378_/CLK _19188_/D vssd1 vssd1 vccd1 vccd1 _19188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18139_ _19830_/Q _18134_/X _18138_/X _18136_/X vssd1 vssd1 vccd1 vccd1 _19830_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10276__S1 _10275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__A _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10050__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09912_ _09767_/A _09890_/Y _09901_/X _09911_/Y _09813_/X vssd1 vssd1 vccd1 vccd1
+ _09912_/X sky130_fd_sc_hd__o311a_1
XFILLER_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09516__A _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09843_ _18937_/Q _18703_/Q _19385_/Q _19033_/Q _10185_/S _09714_/A vssd1 vssd1 vccd1
+ vccd1 _09843_/X sky130_fd_sc_hd__mux4_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17733__A _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _10115_/A vssd1 vssd1 vccd1 vccd1 _09785_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_85_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16349__A _16549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18230__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18230__B2 _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09251__A _16622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10959__A3 _10958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11720__S _12730_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09208_ _09208_/A vssd1 vssd1 vccd1 vccd1 _11589_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10480_ _10480_/A vssd1 vssd1 vccd1 vccd1 _10480_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09139_ _09167_/C vssd1 vssd1 vccd1 vccd1 _09338_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16812__A _16812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12150_ _12126_/A _12151_/C _19411_/Q vssd1 vssd1 vccd1 vccd1 _12150_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11101_ _11072_/A _11098_/Y _11100_/Y _11262_/A vssd1 vssd1 vccd1 vccd1 _11101_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_162_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13647__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12081_ _18112_/A _12021_/A _12022_/X vssd1 vssd1 vccd1 vccd1 _12081_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11032_ _11030_/X _11032_/B vssd1 vssd1 vccd1 vccd1 _11032_/X sky130_fd_sc_hd__and2b_1
XFILLER_77_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14051__B _14787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15840_ _13595_/X _19259_/Q _15848_/S vssd1 vssd1 vccd1 vccd1 _15841_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_9_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19374_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_58_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ _15771_/A vssd1 vssd1 vccd1 vccd1 _19228_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _12983_/A vssd1 vssd1 vccd1 vccd1 _18291_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14478__S _14478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17510_ _17508_/Y _17509_/X _17615_/A vssd1 vssd1 vccd1 vccd1 _17510_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14722_ _14528_/X _18818_/Q _14726_/S vssd1 vssd1 vccd1 vccd1 _14723_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18490_ _19081_/CLK _18490_/D vssd1 vssd1 vccd1 vccd1 _18490_/Q sky130_fd_sc_hd__dfxtp_1
X_11934_ _11969_/B _11934_/B vssd1 vssd1 vccd1 vccd1 _11934_/Y sky130_fd_sc_hd__xnor2_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_22_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17441_ _17497_/S _17249_/X _17440_/X vssd1 vssd1 vccd1 vccd1 _17441_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _14653_/A vssd1 vssd1 vccd1 vccd1 _18787_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11773_/X _11863_/X _11864_/Y _11623_/A vssd1 vssd1 vccd1 vccd1 _11865_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output106_A _17166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__C1 _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13604_ _13604_/A vssd1 vssd1 vccd1 vccd1 _18380_/D sky130_fd_sc_hd__clkbuf_1
X_10816_ _10933_/A vssd1 vssd1 vccd1 vccd1 _10817_/A sky130_fd_sc_hd__clkbuf_4
X_17372_ _17286_/X _17282_/X _17372_/S vssd1 vssd1 vccd1 vccd1 _17372_/X sky130_fd_sc_hd__mux2_1
X_14584_ _14584_/A vssd1 vssd1 vccd1 vccd1 _18766_/D sky130_fd_sc_hd__clkbuf_1
X_11796_ _11796_/A vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19111_ _19329_/CLK _19111_/D vssd1 vssd1 vccd1 vccd1 _19111_/Q sky130_fd_sc_hd__dfxtp_1
X_16323_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__buf_2
XFILLER_41_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ _15019_/A vssd1 vssd1 vccd1 vccd1 _13535_/X sky130_fd_sc_hd__buf_2
X_10747_ _10747_/A vssd1 vssd1 vccd1 vccd1 _10747_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__11630__S _12730_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19042_ _19202_/CLK _19042_/D vssd1 vssd1 vccd1 vccd1 _19042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16254_ _16254_/A vssd1 vssd1 vccd1 vccd1 _19397_/D sky130_fd_sc_hd__clkbuf_1
X_13466_ _13048_/X _18333_/Q _13470_/S vssd1 vssd1 vccd1 vccd1 _13467_/A sky130_fd_sc_hd__mux2_1
X_10678_ _19718_/Q vssd1 vssd1 vccd1 vccd1 _10678_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15205_ _15205_/A vssd1 vssd1 vccd1 vccd1 _19021_/D sky130_fd_sc_hd__clkbuf_1
X_12417_ _12130_/X _12415_/X _12416_/Y _12134_/X vssd1 vssd1 vccd1 vccd1 _12417_/X
+ sky130_fd_sc_hd__a31o_1
X_16185_ _13535_/X _19366_/Q _16191_/S vssd1 vssd1 vccd1 vccd1 _16186_/A sky130_fd_sc_hd__mux2_1
X_13397_ _13397_/A vssd1 vssd1 vccd1 vccd1 _15565_/A sky130_fd_sc_hd__clkbuf_2
X_15136_ _15158_/A vssd1 vssd1 vccd1 vccd1 _15145_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_154_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12348_ _12348_/A _12348_/B _12267_/B _12312_/Y vssd1 vssd1 vccd1 vccd1 _12363_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_126_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10583__A1 _10074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11207__S0 _11243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15067_ _15067_/A vssd1 vssd1 vccd1 vccd1 _15067_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12279_ _19416_/Q _11963_/X _12278_/X vssd1 vssd1 vccd1 vccd1 _12279_/X sky130_fd_sc_hd__o21a_2
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14018_ _18534_/Q _14017_/X _14027_/S vssd1 vssd1 vccd1 vccd1 _14019_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11585__B _18132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15772__S _15776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18826_ _19247_/CLK _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10430__S1 _10270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18757_ _19180_/CLK _18757_/D vssd1 vssd1 vccd1 vccd1 _18757_/Q sky130_fd_sc_hd__dfxtp_1
X_15969_ _15969_/A vssd1 vssd1 vccd1 vccd1 _19316_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12697__A _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15073__A _15073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17708_ _17709_/A _17709_/B _17775_/S vssd1 vssd1 vccd1 vccd1 _17708_/X sky130_fd_sc_hd__mux2_1
X_09490_ _10848_/A vssd1 vssd1 vccd1 vccd1 _10721_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_82_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18688_ _19085_/CLK _18688_/D vssd1 vssd1 vccd1 vccd1 _18688_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10194__S0 _09854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17639_ _17642_/A _17642_/B _17775_/S vssd1 vssd1 vccd1 vccd1 _17639_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16774__A1 _19565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11599__B1 _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19309_ _19309_/CLK _19309_/D vssd1 vssd1 vccd1 vccd1 _19309_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15520__B _15520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10497__S1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17723__A0 _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12260__A1 _18130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09639__S0 _10572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10574__A1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10680__A _10680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15682__S _15682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09826_ _11402_/A _09826_/B vssd1 vssd1 vccd1 vccd1 _09826_/Y sky130_fd_sc_hd__nor2_1
XFILLER_101_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09757_ _09757_/A vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12400__A _17305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09688_ _09688_/A vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_104_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16765__A1 _16772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11650_ _11652_/A vssd1 vssd1 vccd1 vccd1 _12068_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15711__A _15767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10601_ _10612_/A _10601_/B vssd1 vssd1 vccd1 vccd1 _10601_/X sky130_fd_sc_hd__or2_1
XFILLER_168_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11581_ _19861_/Q vssd1 vssd1 vccd1 vccd1 _18135_/A sky130_fd_sc_hd__buf_4
XFILLER_70_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16018__S _16024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13320_ _19692_/Q _12529_/A _12521_/A _19659_/Q vssd1 vssd1 vccd1 vccd1 _13320_/X
+ sky130_fd_sc_hd__a22o_1
X_10532_ _19313_/Q _18725_/Q _18762_/Q _18336_/Q _10481_/S _10262_/A vssd1 vssd1 vccd1
+ vccd1 _10532_/X sky130_fd_sc_hd__mux4_1
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15857__S _15865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13251_ _14598_/A vssd1 vssd1 vccd1 vccd1 _13251_/X sky130_fd_sc_hd__clkbuf_2
X_10463_ _10511_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _10463_/X sky130_fd_sc_hd__or2_1
XFILLER_109_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13200__B1 _13199_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16542__A _19495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12554__A2 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12202_ _12201_/X _12200_/Y _12341_/S vssd1 vssd1 vccd1 vccd1 _12202_/X sky130_fd_sc_hd__mux2_1
X_13182_ _19572_/Q _13006_/X _13181_/X _12538_/X vssd1 vssd1 vccd1 vccd1 _13182_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_input67_A io_irq_motor_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ _10394_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10394_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_142_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19706_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10565__B2 _19721_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _16989_/A _12156_/C vssd1 vssd1 vccd1 vccd1 _12133_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10590__A _10590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17990_ _16159_/A _19800_/Q _17990_/S vssd1 vssd1 vccd1 vccd1 _17991_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12306__A2 _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16941_ _19631_/Q _17010_/A vssd1 vssd1 vccd1 vccd1 _16941_/X sky130_fd_sc_hd__and2_1
X_12064_ _12372_/A vssd1 vssd1 vccd1 vccd1 _12369_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_132_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11015_ _11004_/X _11008_/X _11010_/X _11014_/X _09465_/A vssd1 vssd1 vccd1 vccd1
+ _11015_/X sky130_fd_sc_hd__a221o_2
X_19660_ _19660_/CLK _19660_/D vssd1 vssd1 vccd1 vccd1 _19660_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10412__S1 _10312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16872_ _16871_/A _16871_/C _19602_/Q vssd1 vssd1 vccd1 vccd1 _16873_/C sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_157_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19108_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10868__A2 _10846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18611_ _19074_/CLK _18611_/D vssd1 vssd1 vccd1 vccd1 _18611_/Q sky130_fd_sc_hd__dfxtp_1
X_15823_ _15823_/A vssd1 vssd1 vccd1 vccd1 _19251_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17650__C1 _11539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19591_ _19594_/CLK _19591_/D vssd1 vssd1 vccd1 vccd1 _19591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18542_ _19389_/CLK _18542_/D vssd1 vssd1 vccd1 vccd1 _18542_/Q sky130_fd_sc_hd__dfxtp_1
X_15754_ _13576_/X _19221_/Q _15754_/S vssd1 vssd1 vccd1 vccd1 _15755_/A sky130_fd_sc_hd__mux2_1
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12966_ _19596_/Q _12950_/X _12951_/X _19464_/Q _12965_/X vssd1 vssd1 vccd1 vccd1
+ _15505_/B sky130_fd_sc_hd__a221o_2
XFILLER_79_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10749__B _10749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _14608_/X _18811_/Q _14709_/S vssd1 vssd1 vccd1 vccd1 _14706_/A sky130_fd_sc_hd__mux2_1
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18473_ _19471_/CLK _18473_/D vssd1 vssd1 vccd1 vccd1 _18473_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17820__B _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11917_ _11950_/A _11892_/A _11950_/C _11949_/A vssd1 vssd1 vccd1 vccd1 _11923_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__16756__A1 _16760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15685_ _14585_/X _19190_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15686_/A sky130_fd_sc_hd__mux2_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _19143_/Q _12895_/X _12677_/X _19333_/Q _12896_/X vssd1 vssd1 vccd1 vccd1
+ _12897_/X sky130_fd_sc_hd__a221o_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _17390_/X _17403_/Y _17423_/X vssd1 vssd1 vccd1 vccd1 _17424_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_61_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14636_ _14636_/A vssd1 vssd1 vccd1 vccd1 _18782_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11848_ _11848_/A _11848_/B vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__or2_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ _17216_/X _17220_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17355_/X sky130_fd_sc_hd__mux2_1
X_14567_ _14566_/X _18761_/Q _14567_/S vssd1 vssd1 vccd1 vccd1 _14568_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17705__A0 _19719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11779_ _11773_/X _11777_/Y _11778_/X _11623_/A vssd1 vssd1 vccd1 vccd1 _11779_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_159_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16306_ _12391_/A _16278_/X _12393_/X _12396_/Y _16280_/X vssd1 vssd1 vccd1 vccd1
+ _19421_/D sky130_fd_sc_hd__o221a_1
XFILLER_174_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13518_ _13518_/A vssd1 vssd1 vccd1 vccd1 _18353_/D sky130_fd_sc_hd__clkbuf_1
X_17286_ _12309_/A _17563_/B _17286_/S vssd1 vssd1 vccd1 vccd1 _17286_/X sky130_fd_sc_hd__mux2_1
X_14498_ _13915_/X _18733_/Q _14500_/S vssd1 vssd1 vccd1 vccd1 _14499_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19025_ _19377_/CLK _19025_/D vssd1 vssd1 vccd1 vccd1 _19025_/Q sky130_fd_sc_hd__dfxtp_1
X_16237_ _13611_/X _19390_/Q _16239_/S vssd1 vssd1 vccd1 vccd1 _16238_/A sky130_fd_sc_hd__mux2_1
X_13449_ _13449_/A vssd1 vssd1 vccd1 vccd1 _18325_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12980__A _15025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16168_ _16168_/A vssd1 vssd1 vccd1 vccd1 _19359_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_86_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11596__A _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ _18983_/Q _15022_/X _15123_/S vssd1 vssd1 vccd1 vccd1 _15120_/A sky130_fd_sc_hd__mux2_1
X_16099_ _16107_/C _16098_/Y _13418_/A vssd1 vssd1 vccd1 vccd1 _16099_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_173_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15495__B2 hold15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10403__S1 _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19858_ _19866_/CLK _19858_/D vssd1 vssd1 vccd1 vccd1 _19858_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10005__A _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14700__A _14700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09611_ _09717_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09611_/X sky130_fd_sc_hd__or2_1
XFILLER_95_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18809_ _19391_/CLK _18809_/D vssd1 vssd1 vccd1 vccd1 _18809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19789_ _19800_/CLK _19789_/D vssd1 vssd1 vccd1 vccd1 _19789_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11535__S _11539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15007__S _15013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09542_ _09542_/A vssd1 vssd1 vccd1 vccd1 _09543_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_110_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16747__A1 _16752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ _09665_/A _09452_/X _09467_/X _09756_/A _19736_/Q vssd1 vssd1 vccd1 vccd1
+ _11418_/A sky130_fd_sc_hd__a32o_4
XANTENNA__14846__S _14854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16627__A _16659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13750__S _13758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__A2_N _12448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10890__S1 _10817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17475__A2 _17328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_74_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19382_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09809_ _10129_/A _09808_/X _09767_/X vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__o21a_1
XFILLER_101_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_89_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19618_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12820_ _19553_/Q _12701_/X _12819_/X _12644_/X vssd1 vssd1 vccd1 vccd1 _12820_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_28_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12751_/A vssd1 vssd1 vccd1 vccd1 _12773_/A sky130_fd_sc_hd__buf_4
XANTENNA__10078__A3 _10076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13660__S _13664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _11803_/A _12696_/A _11702_/C _11702_/D vssd1 vssd1 vccd1 vccd1 _11703_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_131_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_12_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _18990_/CLK sky130_fd_sc_hd__clkbuf_16
X_15470_ _15470_/A vssd1 vssd1 vccd1 vccd1 _19139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _19584_/Q _12619_/A _12678_/X _12681_/X vssd1 vssd1 vccd1 vccd1 _12682_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14421_ _14421_/A vssd1 vssd1 vccd1 vccd1 _18698_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _11670_/A _12444_/B _11632_/Y vssd1 vssd1 vccd1 vccd1 _17575_/S sky130_fd_sc_hd__o21ai_4
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17140_ _17140_/A vssd1 vssd1 vccd1 vccd1 _17140_/X sky130_fd_sc_hd__buf_2
X_14352_ _13915_/X _18669_/Q _14354_/S vssd1 vssd1 vccd1 vccd1 _14353_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12775__A2 _12773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11564_ _11577_/B _17183_/B _11564_/C _11563_/X vssd1 vssd1 vccd1 vccd1 _17177_/A
+ sky130_fd_sc_hd__or4b_4
XANTENNA__10330__S0 _10286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _19451_/Q _13005_/X _13302_/X vssd1 vssd1 vccd1 vccd1 _13303_/X sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_27_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _18975_/CLK sky130_fd_sc_hd__clkbuf_16
X_17071_ _17071_/A vssd1 vssd1 vccd1 vccd1 _19682_/D sky130_fd_sc_hd__clkbuf_1
X_10515_ _10511_/A _10512_/X _10514_/X _10243_/A vssd1 vssd1 vccd1 vccd1 _10515_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14283_ input47/X _14282_/X _14277_/X _14278_/X _18122_/A vssd1 vssd1 vccd1 vccd1
+ _18218_/B sky130_fd_sc_hd__a32o_2
XFILLER_6_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11495_ _11495_/A _11495_/B _11495_/C vssd1 vssd1 vccd1 vccd1 _12322_/A sky130_fd_sc_hd__and3_2
XFILLER_10_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10881__S1 _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13185__C1 _13184_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16022_ _16021_/A _16021_/C _16021_/B vssd1 vssd1 vccd1 vccd1 _16023_/B sky130_fd_sc_hd__o21ai_1
X_10446_ _09761_/A _10432_/X _10444_/X _09834_/A _10445_/Y vssd1 vssd1 vccd1 vccd1
+ _12465_/B sky130_fd_sc_hd__o32a_4
X_13234_ _13234_/A _13234_/B _13256_/C vssd1 vssd1 vccd1 vccd1 _13234_/X sky130_fd_sc_hd__or3_1
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__B1 _19396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12932__C1 _12584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10377_ _18930_/Q _18696_/Q _19378_/Q _19026_/Q _10260_/X _10436_/A vssd1 vssd1 vccd1
+ vccd1 _10378_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10002__A3 _10001_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13165_ _13154_/X _13163_/X _13164_/X vssd1 vssd1 vccd1 vccd1 _13165_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_3_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12116_ _12117_/A _17219_/A vssd1 vssd1 vccd1 vccd1 _12118_/A sky130_fd_sc_hd__nand2_1
XFILLER_69_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13488__A0 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13096_ _13095_/A _13111_/C _12832_/A vssd1 vssd1 vccd1 vccd1 _13096_/X sky130_fd_sc_hd__o21a_1
X_17973_ _13195_/X _19792_/Q _17979_/S vssd1 vssd1 vccd1 vccd1 _17974_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13835__S _13835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16924_ _16924_/A vssd1 vssd1 vccd1 vccd1 _19625_/D sky130_fd_sc_hd__clkbuf_1
X_19712_ _19712_/CLK _19712_/D vssd1 vssd1 vccd1 vccd1 _19712_/Q sky130_fd_sc_hd__dfxtp_4
X_12047_ _09194_/X _12021_/X _12022_/X vssd1 vssd1 vccd1 vccd1 _12047_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16211__S _16213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09614__A _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19643_ _19645_/CLK _19643_/D vssd1 vssd1 vccd1 vccd1 _19643_/Q sky130_fd_sc_hd__dfxtp_1
X_16855_ _16854_/A _16854_/C _19596_/Q vssd1 vssd1 vccd1 vccd1 _16856_/C sky130_fd_sc_hd__a21oi_1
XFILLER_120_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16977__A1 _15536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15806_ _15852_/S vssd1 vssd1 vccd1 vccd1 _15815_/S sky130_fd_sc_hd__buf_2
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19574_ _19581_/CLK _19574_/D vssd1 vssd1 vccd1 vccd1 _19574_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17831__A _17831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16786_ _16790_/B _16790_/C _16785_/Y vssd1 vssd1 vccd1 vccd1 _19569_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10149__S0 _09846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13998_ _14030_/A vssd1 vssd1 vccd1 vccd1 _14011_/S sky130_fd_sc_hd__buf_4
X_18525_ _18894_/CLK _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15737_ _13551_/X _19213_/Q _15743_/S vssd1 vssd1 vccd1 vccd1 _15738_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16729__A1 _16731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12949_ _13033_/A vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17042__S _17050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18456_ _19241_/CLK _18456_/D vssd1 vssd1 vccd1 vccd1 _18456_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15668_ _15668_/A vssd1 vssd1 vccd1 vccd1 _19182_/D sky130_fd_sc_hd__clkbuf_1
X_17407_ _17407_/A _17410_/B vssd1 vssd1 vccd1 vccd1 _17418_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17125__D_N _18140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14619_ _14619_/A vssd1 vssd1 vccd1 vccd1 _18777_/D sky130_fd_sc_hd__clkbuf_1
X_18387_ _19202_/CLK _18387_/D vssd1 vssd1 vccd1 vccd1 _18387_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15599_ _15599_/A _18276_/Q vssd1 vssd1 vccd1 vccd1 _15599_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17338_ _17241_/A _17338_/B vssd1 vssd1 vccd1 vccd1 _17338_/X sky130_fd_sc_hd__and2b_1
XFILLER_14_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10777__A1 _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17269_ _17262_/X _17267_/X _17448_/S vssd1 vssd1 vccd1 vccd1 _17269_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16182__A _16239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19008_ _19361_/CLK _19008_/D vssd1 vssd1 vccd1 vccd1 _19008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_144_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10624__S1 _11321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15468__A1 _13410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__13745__S _13747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16417__B1 _16402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11265__S _11265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10701__B2 _10700_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09525_ _10055_/S vssd1 vssd1 vccd1 vccd1 _09776_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_69_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09456_ _09998_/A _09456_/B vssd1 vssd1 vccd1 vccd1 _09456_/X sky130_fd_sc_hd__or2_1
XPHY_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10560__S0 _09415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09387_ _11297_/S vssd1 vssd1 vccd1 vccd1 _10030_/S sky130_fd_sc_hd__buf_4
XFILLER_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12757__A2 _12752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13954__A1 _13953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12824__S _13143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10863__S1 _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15200__S _15206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10300_ _19727_/Q vssd1 vssd1 vccd1 vccd1 _10300_/Y sky130_fd_sc_hd__inv_2
XFILLER_165_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11280_ _11116_/A _11279_/X _11042_/A vssd1 vssd1 vccd1 vccd1 _11280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10231_ _10419_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__or2_1
XFILLER_106_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10615__S1 _09590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10162_ _10174_/A _10162_/B vssd1 vssd1 vccd1 vccd1 _10162_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14970_ _18931_/Q vssd1 vssd1 vccd1 vccd1 _14971_/A sky130_fd_sc_hd__clkbuf_1
X_10093_ _18632_/Q _18967_/Q _10093_/S vssd1 vssd1 vccd1 vccd1 _10093_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09434__A _09434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13921_ _14601_/A vssd1 vssd1 vccd1 vccd1 _13921_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11040__S1 _11033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16640_ _16650_/B _16650_/C vssd1 vssd1 vccd1 vccd1 _16642_/A sky130_fd_sc_hd__and2_1
X_13852_ _13851_/X _18484_/Q _13855_/S vssd1 vssd1 vccd1 vccd1 _13853_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09153__B _11528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15631__A1 _15612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ _16619_/D vssd1 vssd1 vccd1 vccd1 _14715_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_76_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16571_ _19504_/Q _16569_/B _16570_/Y vssd1 vssd1 vccd1 vccd1 _19504_/D sky130_fd_sc_hd__o21a_1
XFILLER_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13783_ _12945_/X _18456_/Q _13787_/S vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__mux2_1
X_10995_ _10990_/X _10993_/X _10994_/X _11048_/A _11007_/A vssd1 vssd1 vccd1 vccd1
+ _11001_/B sky130_fd_sc_hd__o221a_1
XFILLER_43_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18310_ _19325_/CLK _18310_/D vssd1 vssd1 vccd1 vccd1 _18310_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09310__A1 _09315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15522_ _15519_/X _15520_/X _15521_/Y _15508_/X hold16/X vssd1 vssd1 vccd1 vccd1
+ _15522_/X sky130_fd_sc_hd__a32o_4
XFILLER_16_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19290_ _19290_/CLK _19290_/D vssd1 vssd1 vccd1 vccd1 _19290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12734_ _12734_/A vssd1 vssd1 vccd1 vccd1 _18254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18241_ input55/X _14274_/X _18229_/X _18234_/X _17125_/A vssd1 vssd1 vccd1 vccd1
+ _18242_/B sky130_fd_sc_hd__a32o_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _19132_/Q _15089_/X _15455_/S vssd1 vssd1 vccd1 vccd1 _15454_/A sky130_fd_sc_hd__mux2_1
X_12665_ _19532_/Q _12583_/X _12635_/X _19500_/Q _12664_/X vssd1 vssd1 vccd1 vccd1
+ _12665_/X sky130_fd_sc_hd__a221o_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404_ _13883_/X _18691_/Q _14406_/S vssd1 vssd1 vccd1 vccd1 _14405_/A sky130_fd_sc_hd__mux2_1
X_11616_ _16000_/B vssd1 vssd1 vccd1 vccd1 _12184_/A sky130_fd_sc_hd__clkbuf_2
X_18172_ _18172_/A vssd1 vssd1 vccd1 vccd1 _18233_/A sky130_fd_sc_hd__buf_2
X_15384_ _15384_/A vssd1 vssd1 vccd1 vccd1 _19101_/D sky130_fd_sc_hd__clkbuf_1
X_12596_ _14623_/A vssd1 vssd1 vccd1 vccd1 _18234_/A sky130_fd_sc_hd__buf_2
XFILLER_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10759__A1 _09597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17123_ _12482_/A _17114_/X _12021_/X _17119_/X _17122_/X vssd1 vssd1 vccd1 vccd1
+ _17130_/C sky130_fd_sc_hd__a2111o_1
XFILLER_129_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14335_ _13889_/X _18661_/Q _14343_/S vssd1 vssd1 vccd1 vccd1 _14336_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _11623_/A vssd1 vssd1 vccd1 vccd1 _12134_/A sky130_fd_sc_hd__buf_2
XFILLER_117_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15110__S _15112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17054_ _17054_/A vssd1 vssd1 vccd1 vccd1 _19674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output98_A _11765_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14266_ _18639_/Q _14045_/X _14268_/S vssd1 vssd1 vccd1 vccd1 _14267_/A sky130_fd_sc_hd__mux2_1
X_11478_ _10089_/A _11429_/X _11430_/X _11431_/Y _11477_/X vssd1 vssd1 vccd1 vccd1
+ _11478_/X sky130_fd_sc_hd__a221o_1
XFILLER_171_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16005_ _16005_/A vssd1 vssd1 vccd1 vccd1 _19330_/D sky130_fd_sc_hd__clkbuf_1
X_13217_ _19686_/Q _13008_/X _12680_/X _19653_/Q vssd1 vssd1 vccd1 vccd1 _13217_/X
+ sky130_fd_sc_hd__a22o_1
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10429_/Y sky130_fd_sc_hd__nor2_1
X_14197_ _14642_/D _14197_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _15101_/A sky130_fd_sc_hd__or3_2
XANTENNA__10606__S1 _09590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ _14579_/A vssd1 vssd1 vccd1 vccd1 _13148_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_111_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16111__A2 _15582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13565__S _13577_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13079_ _19438_/Q _12636_/X _13078_/X vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__o21a_1
XFILLER_111_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17956_ _17956_/A vssd1 vssd1 vccd1 vccd1 _19752_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16907_ _16907_/A vssd1 vssd1 vccd1 vccd1 _16912_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17887_ _11512_/B _17885_/B _17462_/X _17886_/X vssd1 vssd1 vccd1 vccd1 _17887_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15780__S _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19626_ _19663_/CLK _19626_/D vssd1 vssd1 vccd1 vccd1 _19626_/Q sky130_fd_sc_hd__dfxtp_2
X_16838_ _16838_/A _16838_/B _16838_/C vssd1 vssd1 vccd1 vccd1 _19590_/D sky130_fd_sc_hd__nor3_1
XFILLER_65_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10790__S0 _10692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12436__A1 _19359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16769_ _16778_/C _16772_/C _16772_/D vssd1 vssd1 vccd1 vccd1 _16770_/C sky130_fd_sc_hd__and3_1
X_19557_ _19828_/CLK _19557_/D vssd1 vssd1 vccd1 vccd1 _19557_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09310_ _09315_/B _09306_/A _09309_/X vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_70_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18508_ _18987_/CLK _18508_/D vssd1 vssd1 vccd1 vccd1 _18508_/Q sky130_fd_sc_hd__dfxtp_1
X_19488_ _19619_/CLK _19488_/D vssd1 vssd1 vccd1 vccd1 _19488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ _09241_/A _17133_/A vssd1 vssd1 vccd1 vccd1 _12672_/A sky130_fd_sc_hd__or2_1
X_18439_ _19471_/CLK _18439_/D vssd1 vssd1 vccd1 vccd1 _18439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09172_ _18083_/A _18081_/A _09172_/C _09176_/A vssd1 vssd1 vccd1 vccd1 _09327_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__17678__A2 _17680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09519__A _09519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15955__S _15959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09238__B _18083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11175__A1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16638__B1 _12556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13475__S _13481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12599__B _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10686__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11883__C1 _16109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17190__B _17432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09508_ _18941_/Q _18707_/Q _19389_/Q _19037_/Q _10518_/S _10261_/A vssd1 vssd1 vccd1
+ vccd1 _09509_/B sky130_fd_sc_hd__mux4_1
XFILLER_25_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ _18458_/Q _19049_/Q _19211_/Q _18426_/Q _09519_/A _09506_/A vssd1 vssd1 vccd1
+ vccd1 _10780_/X sky130_fd_sc_hd__mux4_1
XFILLER_13_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17366__A1 _17294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _18606_/Q _18877_/Q _19101_/Q _18845_/Q _10496_/A _09671_/A vssd1 vssd1 vccd1
+ vccd1 _09439_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10339__S _10339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11024__A _11024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12450_/A _12450_/B vssd1 vssd1 vccd1 vccd1 _12450_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17118__A1 _18100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11401_ _18480_/Q _19071_/Q _19233_/Q _18448_/Q _09815_/X _09788_/A vssd1 vssd1 vccd1
+ vccd1 _11402_/B sky130_fd_sc_hd__mux4_1
X_12381_ _17899_/A _12381_/B vssd1 vssd1 vccd1 vccd1 _12385_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11572__A2_N _11918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14120_ _13937_/X _18575_/Q _14122_/S vssd1 vssd1 vccd1 vccd1 _14121_/A sky130_fd_sc_hd__mux2_1
X_11332_ _19311_/Q _18723_/Q _18760_/Q _18334_/Q _10579_/X _10705_/A vssd1 vssd1 vccd1
+ vccd1 _11332_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09429__A _18782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15865__S _15865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14051_ _18089_/A _14787_/B vssd1 vssd1 vccd1 vccd1 _16169_/A sky130_fd_sc_hd__nor2_4
XFILLER_141_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11263_ _18481_/Q _18976_/Q _11263_/S vssd1 vssd1 vccd1 vccd1 _11264_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11166__A1 _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13002_ _19598_/Q vssd1 vssd1 vccd1 vccd1 _16862_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10214_ _10214_/A _10214_/B vssd1 vssd1 vccd1 vccd1 _10214_/Y sky130_fd_sc_hd__nor2_1
XFILLER_134_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11194_ _18913_/Q _18679_/Q _19361_/Q _19009_/Q _11243_/S _11177_/A vssd1 vssd1 vccd1
+ vccd1 _11195_/B sky130_fd_sc_hd__mux4_1
XFILLER_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11261__S1 _11220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10145_ _10105_/A _10144_/X _09857_/X vssd1 vssd1 vccd1 vccd1 _10145_/X sky130_fd_sc_hd__o21a_1
X_17810_ _17810_/A _17810_/B vssd1 vssd1 vccd1 vccd1 _17812_/B sky130_fd_sc_hd__nand2_1
X_18790_ _19241_/CLK _18790_/D vssd1 vssd1 vccd1 vccd1 _18790_/Q sky130_fd_sc_hd__dfxtp_1
X_17741_ _17717_/S _17740_/Y _17402_/A vssd1 vssd1 vccd1 vccd1 _17741_/X sky130_fd_sc_hd__a21o_1
XFILLER_130_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14953_ _14953_/A vssd1 vssd1 vccd1 vccd1 _18922_/D sky130_fd_sc_hd__clkbuf_1
X_10076_ _10067_/Y _10069_/Y _10071_/Y _10075_/Y _09829_/A vssd1 vssd1 vccd1 vccd1
+ _10076_/X sky130_fd_sc_hd__o221a_2
XFILLER_130_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11013__S1 _11012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ _13904_/A vssd1 vssd1 vccd1 vccd1 _18500_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17672_ _17672_/A vssd1 vssd1 vccd1 vccd1 _17673_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14884_ _14930_/S vssd1 vssd1 vccd1 vccd1 _14893_/S sky130_fd_sc_hd__buf_2
XFILLER_48_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16623_ _16623_/A _16623_/B _19816_/Q _19815_/Q vssd1 vssd1 vccd1 vccd1 _16624_/B
+ sky130_fd_sc_hd__or4_1
X_19411_ _19649_/CLK _19411_/D vssd1 vssd1 vccd1 vccd1 _19411_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13835_ _13386_/X _18480_/Q _13835_/S vssd1 vssd1 vccd1 vccd1 _13836_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16554_ _16570_/A _16559_/C vssd1 vssd1 vccd1 vccd1 _16554_/Y sky130_fd_sc_hd__nor2_1
X_19342_ _19759_/CLK _19342_/D vssd1 vssd1 vccd1 vccd1 _19342_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ _13822_/A vssd1 vssd1 vccd1 vccd1 _13835_/S sky130_fd_sc_hd__buf_6
X_10978_ _19304_/Q _18716_/Q _18753_/Q _18327_/Q _10852_/S _10837_/A vssd1 vssd1 vccd1
+ vccd1 _10978_/X sky130_fd_sc_hd__mux4_1
X_15505_ hold12/A _15505_/B vssd1 vssd1 vccd1 vccd1 _15505_/X sky130_fd_sc_hd__or2_1
X_12717_ _19587_/Q _12716_/X _14518_/B vssd1 vssd1 vccd1 vccd1 _12717_/X sky130_fd_sc_hd__mux2_1
X_19273_ _19305_/CLK _19273_/D vssd1 vssd1 vccd1 vccd1 _19273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16485_ _16485_/A _16485_/B _16485_/C vssd1 vssd1 vccd1 vccd1 _19479_/D sky130_fd_sc_hd__nor3_1
X_13697_ _12828_/X _18418_/Q _13703_/S vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16725__A _16754_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18224_ _18224_/A _18224_/B vssd1 vssd1 vccd1 vccd1 _18225_/A sky130_fd_sc_hd__and2_1
XFILLER_30_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15436_ _19124_/Q _15063_/X _15444_/S vssd1 vssd1 vccd1 vccd1 _15437_/A sky130_fd_sc_hd__mux2_1
X_12648_ _19599_/Q _12633_/X _12634_/X _19467_/Q _12647_/X vssd1 vssd1 vccd1 vccd1
+ _12649_/B sky130_fd_sc_hd__a221o_2
XFILLER_50_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18155_ _18197_/A vssd1 vssd1 vccd1 vccd1 _18155_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15367_ _15367_/A vssd1 vssd1 vccd1 vccd1 _19093_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12579_ _19682_/Q _12601_/A _12566_/X _19346_/Q vssd1 vssd1 vccd1 vccd1 _12579_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_11_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17106_ _17124_/B _17105_/X _11556_/B _17108_/B _11508_/A vssd1 vssd1 vccd1 vccd1
+ _17107_/A sky130_fd_sc_hd__o221a_1
XFILLER_129_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09339__A _18122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14318_ _14318_/A vssd1 vssd1 vccd1 vccd1 _18653_/D sky130_fd_sc_hd__clkbuf_1
X_18086_ _18134_/A vssd1 vssd1 vccd1 vccd1 _18086_/X sky130_fd_sc_hd__buf_2
XFILLER_172_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15298_ _14595_/X _19063_/Q _15300_/S vssd1 vssd1 vccd1 vccd1 _15299_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17037_ _19667_/Q _16935_/A _17039_/S vssd1 vssd1 vccd1 vccd1 _17038_/A sky130_fd_sc_hd__mux2_1
X_14249_ _18631_/Q _14020_/X _14253_/S vssd1 vssd1 vccd1 vccd1 _14250_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_17_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11157__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17293__A0 _12405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13295__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15076__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _10277_/A vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__clkbuf_2
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _19098_/CLK _18988_/D vssd1 vssd1 vccd1 vccd1 _18988_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17939_ _17939_/A vssd1 vssd1 vccd1 vccd1 _19744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19609_ _19618_/CLK _19609_/D vssd1 vssd1 vccd1 vccd1 _19609_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12409__A1 _12391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14854__S _14854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16635__A _16666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ _19857_/Q vssd1 vssd1 vccd1 vccd1 _11619_/A sky130_fd_sc_hd__buf_2
XFILLER_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16308__C1 _12556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12042__C1 _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ _17166_/B _11577_/B _17166_/C vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__or3_2
XANTENNA__10818__S1 _10817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09086_ _19849_/Q _19848_/Q vssd1 vssd1 vccd1 vccd1 _09167_/A sky130_fd_sc_hd__or2_1
XFILLER_174_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15685__S _15693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15531__A0 _19719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13994__A _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12403__A _17907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ _10612_/A _09988_/B vssd1 vssd1 vccd1 vccd1 _09988_/X sky130_fd_sc_hd__or2_1
XFILLER_103_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11019__A _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ _11950_/A _17662_/A _11950_/C _17680_/A vssd1 vssd1 vccd1 vccd1 _12025_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_85_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10754__S0 _10650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09712__A _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ _10968_/A vssd1 vssd1 vccd1 vccd1 _11262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ _11880_/Y _11877_/Y _14275_/B vssd1 vssd1 vccd1 vccd1 _11881_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10858__A _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ _15926_/A _14299_/A vssd1 vssd1 vccd1 vccd1 _13677_/A sky130_fd_sc_hd__nand2_4
XFILLER_26_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13234__A _13234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10832_ _09432_/A _10823_/X _10827_/X _10831_/X _11307_/A vssd1 vssd1 vccd1 vccd1
+ _10832_/X sky130_fd_sc_hd__a311o_2
XANTENNA__13073__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13551_ _15035_/A vssd1 vssd1 vccd1 vccd1 _13551_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12820__A1 _19553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14764__S _14770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10763_ _18618_/Q _18953_/Q _10763_/S vssd1 vssd1 vccd1 vccd1 _10763_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _13356_/B vssd1 vssd1 vccd1 vccd1 _12503_/A sky130_fd_sc_hd__buf_2
XFILLER_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16270_ _11969_/C _12319_/X _11974_/X _16269_/X vssd1 vssd1 vccd1 vccd1 _19404_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13482_ _13482_/A vssd1 vssd1 vccd1 vccd1 _18340_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10694_ _09547_/X _10691_/Y _10693_/Y _09644_/A vssd1 vssd1 vccd1 vccd1 _10694_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_12_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15221_ _15221_/A vssd1 vssd1 vccd1 vccd1 _19028_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11689__A _19331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ _12432_/A _12432_/B _12369_/A vssd1 vssd1 vccd1 vccd1 _12433_/Y sky130_fd_sc_hd__a21boi_2
XFILLER_139_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14065__A _14122_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15152_ _18998_/Q _15070_/X _15156_/S vssd1 vssd1 vccd1 vccd1 _15153_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ _12388_/B _12364_/B vssd1 vssd1 vccd1 vccd1 _12365_/A sky130_fd_sc_hd__and2_1
XFILLER_165_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14103_ _13912_/X _18567_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _14104_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11315_ _11309_/A _11314_/X _09602_/X vssd1 vssd1 vccd1 vccd1 _11315_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15083_ _15083_/A vssd1 vssd1 vccd1 vccd1 _15083_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16280__A _18136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12295_ _12294_/Y _12291_/Y _12341_/S vssd1 vssd1 vccd1 vccd1 _12295_/X sky130_fd_sc_hd__mux2_1
XFILLER_107_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14034_ _18539_/Q _14033_/X _14043_/S vssd1 vssd1 vccd1 vccd1 _14035_/A sky130_fd_sc_hd__mux2_1
X_18911_ _19297_/CLK _18911_/D vssd1 vssd1 vccd1 vccd1 _18911_/Q sky130_fd_sc_hd__dfxtp_1
X_11246_ _18577_/Q _18848_/Q _19072_/Q _18816_/Q _09410_/A _11124_/X vssd1 vssd1 vccd1
+ vccd1 _11246_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17275__A0 _17810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18842_ _19386_/CLK _18842_/D vssd1 vssd1 vccd1 vccd1 _18842_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11177_ _11177_/A vssd1 vssd1 vccd1 vccd1 _11177_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10128_ _18472_/Q _19063_/Q _19225_/Q _18440_/Q _09786_/A _10169_/A vssd1 vssd1 vccd1
+ vccd1 _10129_/B sky130_fd_sc_hd__mux4_1
X_18773_ _19324_/CLK _18773_/D vssd1 vssd1 vccd1 vccd1 _18773_/Q sky130_fd_sc_hd__dfxtp_1
X_15985_ _15985_/A vssd1 vssd1 vccd1 vccd1 _19323_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17724_ _17724_/A _17724_/B vssd1 vssd1 vccd1 vccd1 _17724_/Y sky130_fd_sc_hd__nand2_1
X_10059_ _10640_/A vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__buf_4
X_14936_ _18914_/Q vssd1 vssd1 vccd1 vccd1 _14937_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_76_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11311__A1 _09597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15589__A0 _19729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14867_ _18882_/Q _13956_/X _14871_/S vssd1 vssd1 vccd1 vccd1 _14868_/A sky130_fd_sc_hd__mux2_1
X_17655_ _17535_/B _17655_/B vssd1 vssd1 vccd1 vccd1 _17655_/X sky130_fd_sc_hd__and2b_1
XFILLER_35_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16606_ _19516_/Q _16609_/C vssd1 vssd1 vccd1 vccd1 _16607_/B sky130_fd_sc_hd__and2_1
X_13818_ _13240_/X _18472_/Q _13820_/S vssd1 vssd1 vccd1 vccd1 _13819_/A sky130_fd_sc_hd__mux2_1
XFILLER_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17586_ _17603_/A vssd1 vssd1 vccd1 vccd1 _17586_/X sky130_fd_sc_hd__clkbuf_2
X_14798_ _14798_/A vssd1 vssd1 vccd1 vccd1 _18851_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16537_ _16540_/B _16540_/C _16489_/X vssd1 vssd1 vccd1 vccd1 _16537_/Y sky130_fd_sc_hd__a21oi_1
X_19325_ _19325_/CLK _19325_/D vssd1 vssd1 vccd1 vccd1 _19325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14674__S _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ _13749_/A vssd1 vssd1 vccd1 vccd1 _13758_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17050__S _17050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11170__S0 _11011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16468_ _16485_/A _16468_/B _16468_/C vssd1 vssd1 vccd1 vccd1 _19473_/D sky130_fd_sc_hd__nor3_1
X_19256_ _19256_/CLK _19256_/D vssd1 vssd1 vccd1 vccd1 _19256_/Q sky130_fd_sc_hd__dfxtp_1
X_18207_ _18213_/A _18207_/B vssd1 vssd1 vccd1 vccd1 _18208_/A sky130_fd_sc_hd__and2_1
X_15419_ _15419_/A vssd1 vssd1 vccd1 vccd1 _19116_/D sky130_fd_sc_hd__clkbuf_1
X_19187_ _19315_/CLK _19187_/D vssd1 vssd1 vccd1 vccd1 _19187_/Q sky130_fd_sc_hd__dfxtp_1
X_16399_ _19449_/Q _16399_/B vssd1 vssd1 vccd1 vccd1 _16406_/C sky130_fd_sc_hd__and2_1
XFILLER_157_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18138_ _18138_/A _18146_/B vssd1 vssd1 vccd1 vccd1 _18138_/X sky130_fd_sc_hd__or2_1
XFILLER_117_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10050__A1 _09665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18069_ _18150_/A _18069_/B vssd1 vssd1 vccd1 vccd1 _18070_/A sky130_fd_sc_hd__or2_1
XFILLER_105_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09991__A1 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10050__B2 _19734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09911_ _10174_/A _09906_/X _09910_/X vssd1 vssd1 vccd1 vccd1 _09911_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10338__C1 _09831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09842_ _10138_/A _09840_/X _10195_/A vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__a21o_1
XFILLER_98_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09773_/A vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__buf_2
XFILLER_112_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15534__A hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_clock clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__17569__A1 _19712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09532__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10678__A _19718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11161__S0 _09496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09207_ _09207_/A _11567_/A _11526_/A vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__or3b_4
XFILLER_120_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09138_ _19862_/Q _19861_/Q _19860_/Q vssd1 vssd1 vccd1 vccd1 _09167_/C sky130_fd_sc_hd__or3_2
XFILLER_108_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12117__B _17219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ _11100_/A _11100_/B vssd1 vssd1 vccd1 vccd1 _11100_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_192_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__A _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12080_ _12066_/B _11963_/X _12073_/Y _12079_/Y vssd1 vssd1 vccd1 vccd1 _12080_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_78_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11031_ _18486_/Q _18981_/Q _11151_/S vssd1 vssd1 vccd1 vccd1 _11032_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13818__A0 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14759__S _14759_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15770_ _13599_/X _19228_/Q _15776_/S vssd1 vssd1 vccd1 vccd1 _15771_/A sky130_fd_sc_hd__mux2_1
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12981_/X _18291_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12983_/A sky130_fd_sc_hd__mux2_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input12_A io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14721_ _14721_/A vssd1 vssd1 vccd1 vccd1 _18817_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ _19403_/Q vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17440_ _17446_/S _17440_/B vssd1 vssd1 vccd1 vccd1 _17440_/X sky130_fd_sc_hd__or2_1
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14531_/X _18787_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14653_/A sky130_fd_sc_hd__mux2_1
X_11864_ _16963_/A _11886_/C vssd1 vssd1 vccd1 vccd1 _11864_/Y sky130_fd_sc_hd__nand2_1
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13046__A1 _11538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13603_ _18380_/Q _13602_/X _13609_/S vssd1 vssd1 vccd1 vccd1 _13604_/A sky130_fd_sc_hd__mux2_1
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _18780_/Q vssd1 vssd1 vccd1 vccd1 _10933_/A sky130_fd_sc_hd__clkbuf_2
X_17371_ _17283_/X _17270_/X _17372_/S vssd1 vssd1 vccd1 vccd1 _17371_/X sky130_fd_sc_hd__mux2_1
X_14583_ _14582_/X _18766_/Q _14583_/S vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14494__S _14500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11795_ _11826_/A _12098_/C vssd1 vssd1 vccd1 vccd1 _11795_/Y sky130_fd_sc_hd__xnor2_1
X_16322_ _16341_/A _16322_/B _16322_/C vssd1 vssd1 vccd1 vccd1 _19424_/D sky130_fd_sc_hd__nor3_1
XANTENNA__09588__S _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19110_ _19329_/CLK _19110_/D vssd1 vssd1 vccd1 vccd1 _19110_/Q sky130_fd_sc_hd__dfxtp_1
X_13534_ _13534_/A vssd1 vssd1 vccd1 vccd1 _18358_/D sky130_fd_sc_hd__clkbuf_1
X_10746_ _10739_/Y _10741_/Y _10743_/Y _10745_/Y _11307_/A vssd1 vssd1 vccd1 vccd1
+ _10747_/A sky130_fd_sc_hd__o221a_1
XFILLER_40_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19041_ _19235_/CLK _19041_/D vssd1 vssd1 vccd1 vccd1 _19041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16253_ _16255_/A _16253_/B vssd1 vssd1 vccd1 vccd1 _16254_/A sky130_fd_sc_hd__or2_1
XANTENNA__15743__A0 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ _13465_/A vssd1 vssd1 vccd1 vccd1 _18332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10677_ _10677_/A vssd1 vssd1 vccd1 vccd1 _11456_/A sky130_fd_sc_hd__inv_2
XFILLER_139_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15204_ _19021_/Q _15041_/X _15206_/S vssd1 vssd1 vccd1 vccd1 _15205_/A sky130_fd_sc_hd__mux2_1
X_12416_ _17020_/A _12416_/B vssd1 vssd1 vccd1 vccd1 _12416_/Y sky130_fd_sc_hd__nand2_1
XFILLER_173_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16184_ _16184_/A vssd1 vssd1 vccd1 vccd1 _19365_/D sky130_fd_sc_hd__clkbuf_1
X_13396_ _13396_/A vssd1 vssd1 vccd1 vccd1 _18315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15135_ _15135_/A vssd1 vssd1 vccd1 vccd1 _18990_/D sky130_fd_sc_hd__clkbuf_1
X_12347_ _12347_/A _12347_/B vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__nand2_1
XFILLER_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11780__A1 _19397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output80_A _12123_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15066_ _15066_/A vssd1 vssd1 vccd1 vccd1 _18964_/D sky130_fd_sc_hd__clkbuf_1
X_12278_ _12071_/X _12273_/X _12274_/X _12277_/X _12134_/A vssd1 vssd1 vccd1 vccd1
+ _12278_/X sky130_fd_sc_hd__a311o_1
XANTENNA__11207__S1 _11177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14017_ _14589_/A vssd1 vssd1 vccd1 vccd1 _14017_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11229_ _19299_/Q _18711_/Q _18748_/Q _18322_/Q _10969_/A _09511_/A vssd1 vssd1 vccd1
+ vccd1 _11229_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18825_ _19308_/CLK _18825_/D vssd1 vssd1 vccd1 vccd1 _18825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16471__A1 _19474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18756_ _19307_/CLK _18756_/D vssd1 vssd1 vccd1 vccd1 _18756_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15968_ _13573_/X _19316_/Q _15970_/S vssd1 vssd1 vccd1 vccd1 _15969_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10718__S0 _09645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17707_ _17392_/X _17444_/A _17402_/X vssd1 vssd1 vccd1 vccd1 _17707_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14919_ _14919_/A vssd1 vssd1 vccd1 vccd1 _18905_/D sky130_fd_sc_hd__clkbuf_1
X_15899_ _15899_/A vssd1 vssd1 vccd1 vccd1 _19285_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10498__A _10509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18687_ _19081_/CLK _18687_/D vssd1 vssd1 vccd1 vccd1 _18687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10194__S1 _09676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17638_ _17479_/X _17574_/A _17483_/X vssd1 vssd1 vccd1 vccd1 _17827_/B sky130_fd_sc_hd__a21oi_2
XFILLER_24_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17971__A1 _19791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17569_ _19712_/Q _09322_/X _17567_/X _17568_/Y vssd1 vssd1 vccd1 vccd1 _19712_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11599__A1 _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19308_ _19308_/CLK _19308_/D vssd1 vssd1 vccd1 vccd1 _19308_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13602__A _15086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17723__A1 _17722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19239_ _19239_/CLK _19239_/D vssd1 vssd1 vccd1 vccd1 _19239_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11122__A _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09639__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11771__A1 _11765_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09527__A _10347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input4_A io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09825_ _18477_/Q _19068_/Q _19230_/Q _18445_/Q _09815_/X _09799_/X vssd1 vssd1 vccd1
+ vccd1 _09826_/B sky130_fd_sc_hd__mux4_1
XFILLER_171_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09756_ _09756_/A vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__buf_2
XFILLER_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09687_ _09687_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _09687_/X sky130_fd_sc_hd__and2_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_139_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10600_ _18924_/Q _18690_/Q _19372_/Q _19020_/Q _10546_/S _09419_/A vssd1 vssd1 vccd1
+ vccd1 _10601_/B sky130_fd_sc_hd__mux4_1
XFILLER_23_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ _12442_/B vssd1 vssd1 vccd1 vccd1 _11580_/Y sky130_fd_sc_hd__inv_2
XFILLER_70_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10531_ _10531_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10531_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_129_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13250_ _15076_/A vssd1 vssd1 vccd1 vccd1 _14598_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10462_ _19314_/Q _18726_/Q _18763_/Q _18337_/Q _10499_/S _10311_/A vssd1 vssd1 vccd1
+ vccd1 _10463_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16542__B _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13658__S _13664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ _19413_/Q _12201_/B vssd1 vssd1 vccd1 vccd1 _12201_/X sky130_fd_sc_hd__xor2_1
XFILLER_136_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13181_ _19158_/Q _13179_/X _12958_/X _19348_/Q _13180_/X vssd1 vssd1 vccd1 vccd1
+ _13181_/X sky130_fd_sc_hd__a221o_2
XFILLER_164_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10393_ _18467_/Q _19058_/Q _19220_/Q _18435_/Q _10274_/X _10275_/X vssd1 vssd1 vccd1
+ vccd1 _10394_/B sky130_fd_sc_hd__mux4_1
XFILLER_135_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10871__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10565__A2 _10555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12132_ _16989_/A _12156_/C vssd1 vssd1 vccd1 vccd1 _12132_/X sky130_fd_sc_hd__or2_1
XFILLER_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16940_ _16946_/A vssd1 vssd1 vccd1 vccd1 _17010_/A sky130_fd_sc_hd__clkbuf_2
X_12063_ _12435_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ _11171_/A _11013_/X _09447_/A vssd1 vssd1 vccd1 vccd1 _11014_/X sky130_fd_sc_hd__o21a_1
XFILLER_78_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14489__S _14489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16871_ _16871_/A _19602_/Q _16871_/C vssd1 vssd1 vccd1 vccd1 _16873_/B sky130_fd_sc_hd__and3_1
XANTENNA__10868__A3 _10866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12798__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18610_ _19361_/CLK _18610_/D vssd1 vssd1 vccd1 vccd1 _18610_/Q sky130_fd_sc_hd__dfxtp_1
X_15822_ _13570_/X _19251_/Q _15826_/S vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__mux2_1
X_19590_ _19688_/CLK _19590_/D vssd1 vssd1 vccd1 vccd1 _19590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09172__A _18083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15753_ _15753_/A vssd1 vssd1 vccd1 vccd1 _19220_/D sky130_fd_sc_hd__clkbuf_1
X_18541_ _19325_/CLK _18541_/D vssd1 vssd1 vccd1 vccd1 _18541_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12965_ _19528_/Q _12952_/X _12953_/X _16551_/B _12964_/X vssd1 vssd1 vccd1 vccd1
+ _12965_/X sky130_fd_sc_hd__a221o_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ _12134_/A _11911_/Y _11914_/X _11915_/X vssd1 vssd1 vccd1 vccd1 _16264_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_46_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14704_ _14704_/A vssd1 vssd1 vccd1 vccd1 _18810_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18472_ _19382_/CLK _18472_/D vssd1 vssd1 vccd1 vccd1 _18472_/Q sky130_fd_sc_hd__dfxtp_1
X_15684_ _15695_/A vssd1 vssd1 vccd1 vccd1 _15693_/S sky130_fd_sc_hd__buf_4
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ _19669_/Q _12817_/X _12680_/A _19636_/Q vssd1 vssd1 vccd1 vccd1 _12896_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17953__A1 _19783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ _17414_/X _17418_/Y _17420_/X _17733_/A vssd1 vssd1 vccd1 vccd1 _17423_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14635_ _14635_/A _18211_/B vssd1 vssd1 vccd1 vccd1 _14636_/A sky130_fd_sc_hd__and2_1
XFILLER_127_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _11847_/A _17198_/A vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__nor2_1
XANTENNA__16209__S _16213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14518__A _16833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11125__S0 _11173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13422__A _16109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14566_ _14566_/A vssd1 vssd1 vccd1 vccd1 _14566_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17354_ _17498_/B _17353_/X _17501_/S vssd1 vssd1 vccd1 vccd1 _17548_/B sky130_fd_sc_hd__mux2_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ _16953_/A _11778_/B _11778_/C vssd1 vssd1 vccd1 vccd1 _11778_/X sky130_fd_sc_hd__or3_1
XANTENNA__17705__A1 _17704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16305_ _12366_/Y _12134_/X _12375_/X _16914_/A vssd1 vssd1 vccd1 vccd1 _19420_/D
+ sky130_fd_sc_hd__a211oi_1
X_13517_ _18353_/Q _13509_/X _13529_/S vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__mux2_1
X_17285_ _12349_/A _17252_/X _17286_/S vssd1 vssd1 vccd1 vccd1 _17285_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10729_ _18619_/Q _18954_/Q _10729_/S vssd1 vssd1 vccd1 vccd1 _10729_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14497_ _14497_/A vssd1 vssd1 vccd1 vccd1 _18732_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12038__A _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19024_ _19376_/CLK _19024_/D vssd1 vssd1 vccd1 vccd1 _19024_/Q sky130_fd_sc_hd__dfxtp_1
X_16236_ _16236_/A vssd1 vssd1 vccd1 vccd1 _19389_/D sky130_fd_sc_hd__clkbuf_1
X_13448_ _12886_/X _18325_/Q _13448_/S vssd1 vssd1 vccd1 vccd1 _13449_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_174_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13568__S _13577_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _16166_/X _19359_/Q _16167_/S vssd1 vssd1 vccd1 vccd1 _16168_/A sky130_fd_sc_hd__mux2_1
X_13379_ _19551_/Q _13004_/X _13054_/X _19519_/Q _13378_/X vssd1 vssd1 vccd1 vccd1
+ _13379_/X sky130_fd_sc_hd__a221o_1
XFILLER_154_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15118_ _15118_/A vssd1 vssd1 vccd1 vccd1 _18982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16098_ _19758_/Q _16098_/B vssd1 vssd1 vccd1 vccd1 _16098_/Y sky130_fd_sc_hd__nand2_1
XFILLER_141_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15049_ _18959_/Q _15047_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15050_/A sky130_fd_sc_hd__mux2_1
XFILLER_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19857_ _19866_/CLK _19857_/D vssd1 vssd1 vccd1 vccd1 _19857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09610_ _19296_/Q _19134_/Q _18543_/Q _18313_/Q _09599_/X _09977_/A vssd1 vssd1 vccd1
+ vccd1 _09611_/B sky130_fd_sc_hd__mux4_1
X_18808_ _19384_/CLK _18808_/D vssd1 vssd1 vccd1 vccd1 _18808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19788_ _19800_/CLK _19788_/D vssd1 vssd1 vccd1 vccd1 _19788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09541_ _09541_/A vssd1 vssd1 vccd1 vccd1 _09542_/A sky130_fd_sc_hd__buf_4
X_18739_ _19375_/CLK _18739_/D vssd1 vssd1 vccd1 vccd1 _18739_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12220__B _17819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16908__A _16915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09472_ _09472_/A vssd1 vssd1 vccd1 vccd1 _09756_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_140_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15955__A0 _13554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10956__A _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11992__A1 _19341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _18987_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_165_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__A0 _19714_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_65_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15693__S _15693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09808_ _18605_/Q _18876_/Q _19100_/Q _18844_/Q _11387_/A _09785_/A vssd1 vssd1 vccd1
+ vccd1 _09808_/X sky130_fd_sc_hd__mux4_1
XFILLER_47_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09739_ _09857_/A vssd1 vssd1 vccd1 vccd1 _09740_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13941__S _13941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ _18263_/Q _12744_/X _10648_/A _12747_/X vssd1 vssd1 vccd1 vccd1 _18263_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _16619_/B _12621_/B vssd1 vssd1 vccd1 vccd1 _11702_/C sky130_fd_sc_hd__or2_1
XANTENNA__10483__A1 _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15946__A0 _13541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12681_ _19687_/Q _12659_/X _12680_/X _19654_/Q vssd1 vssd1 vccd1 vccd1 _12681_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14420_ _13905_/X _18698_/Q _14428_/S vssd1 vssd1 vccd1 vccd1 _14421_/A sky130_fd_sc_hd__mux2_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _09207_/X _11630_/X _11631_/X vssd1 vssd1 vccd1 vccd1 _11632_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_168_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14351_ _14351_/A vssd1 vssd1 vccd1 vccd1 _18668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11563_ _11565_/A _11487_/S _09146_/C _11646_/B _11559_/A vssd1 vssd1 vccd1 vccd1
+ _11563_/X sky130_fd_sc_hd__a2111o_1
XFILLER_129_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ hold22/A _13006_/X _13301_/X _13012_/X vssd1 vssd1 vccd1 vccd1 _13302_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10330__S1 _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17070_ _19682_/Q _12593_/B _17072_/S vssd1 vssd1 vccd1 vccd1 _17071_/A sky130_fd_sc_hd__mux2_1
X_10514_ _10514_/A _10514_/B vssd1 vssd1 vccd1 vccd1 _10514_/X sky130_fd_sc_hd__or2_1
X_14282_ _18197_/A vssd1 vssd1 vccd1 vccd1 _14282_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _11490_/X _11481_/X _11492_/Y _11493_/X vssd1 vssd1 vccd1 vccd1 _11495_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16272__B _16272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16021_ _16021_/A _16021_/B _16021_/C vssd1 vssd1 vccd1 vccd1 _16028_/B sky130_fd_sc_hd__or3_1
X_13233_ _19762_/Q _13233_/B vssd1 vssd1 vccd1 vccd1 _13256_/C sky130_fd_sc_hd__and2_1
XFILLER_143_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10445_ _19724_/Q vssd1 vssd1 vccd1 vccd1 _10445_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11735__A1 _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12932__B1 _12606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16123__A0 _12689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ _13164_/A vssd1 vssd1 vccd1 vccd1 _13164_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_156_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10376_ _09666_/A _10364_/X _10375_/X _09757_/A _19725_/Q vssd1 vssd1 vccd1 vccd1
+ _10401_/A sky130_fd_sc_hd__a32o_4
XFILLER_112_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output166_A _12441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12115_ _19789_/Q _10401_/A _12423_/S vssd1 vssd1 vccd1 vccd1 _17219_/A sky130_fd_sc_hd__mux2_2
XFILLER_152_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13095_ _13095_/A _13111_/C vssd1 vssd1 vccd1 vccd1 _13095_/Y sky130_fd_sc_hd__nand2_1
X_17972_ _17972_/A vssd1 vssd1 vccd1 vccd1 _19759_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14801__A _14858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19711_ _19711_/CLK _19711_/D vssd1 vssd1 vccd1 vccd1 _19711_/Q sky130_fd_sc_hd__dfxtp_4
X_16923_ _19625_/Q _16932_/A _17026_/S vssd1 vssd1 vccd1 vccd1 _16924_/A sky130_fd_sc_hd__mux2_1
X_12046_ _12066_/A _12078_/A _12042_/X _12045_/Y vssd1 vssd1 vccd1 vccd1 _16276_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12160__A1 _09351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15108__S _15112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19642_ _19645_/CLK _19642_/D vssd1 vssd1 vccd1 vccd1 _19642_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16854_ _16854_/A _19596_/Q _16854_/C vssd1 vssd1 vccd1 vccd1 _16856_/B sky130_fd_sc_hd__and3_1
XANTENNA__12321__A _12321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15805_ _15805_/A vssd1 vssd1 vccd1 vccd1 _19243_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19573_ _19668_/CLK _19573_/D vssd1 vssd1 vccd1 vccd1 _19573_/Q sky130_fd_sc_hd__dfxtp_1
X_16785_ _16790_/B _16790_/C _16764_/X vssd1 vssd1 vccd1 vccd1 _16785_/Y sky130_fd_sc_hd__a21oi_1
X_13997_ _14569_/A vssd1 vssd1 vccd1 vccd1 _13997_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__18179__B2 _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10149__S1 _09871_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18524_ _19278_/CLK _18524_/D vssd1 vssd1 vccd1 vccd1 _18524_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15736_ _15736_/A vssd1 vssd1 vccd1 vccd1 _19212_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12948_ _13065_/A vssd1 vssd1 vccd1 vccd1 _13033_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15937__A0 _13528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18455_ _19241_/CLK _18455_/D vssd1 vssd1 vccd1 vccd1 _18455_/Q sky130_fd_sc_hd__dfxtp_1
X_12879_ _16650_/B _12782_/X _12699_/X _19492_/Q _12878_/X vssd1 vssd1 vccd1 vccd1
+ _12879_/X sky130_fd_sc_hd__a221o_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15667_ _14560_/X _19182_/Q _15671_/S vssd1 vssd1 vccd1 vccd1 _15668_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17406_ _17844_/S vssd1 vssd1 vccd1 vccd1 _17406_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14618_ _14617_/X _18777_/Q _14621_/S vssd1 vssd1 vccd1 vccd1 _14619_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13412__A1 _13410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15598_ _18276_/Q _15598_/B vssd1 vssd1 vccd1 vccd1 _15598_/X sky130_fd_sc_hd__or2_1
XFILLER_21_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18386_ _19235_/CLK _18386_/D vssd1 vssd1 vccd1 vccd1 _18386_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15778__S _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14549_ _14549_/A vssd1 vssd1 vccd1 vccd1 _18755_/D sky130_fd_sc_hd__clkbuf_1
X_17337_ _17305_/A _17372_/S _17305_/B vssd1 vssd1 vccd1 vccd1 _17337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_147_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17268_ _17501_/S vssd1 vssd1 vccd1 vccd1 _17448_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_146_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19007_ _19731_/CLK _19007_/D vssd1 vssd1 vccd1 vccd1 _19007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_161_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16219_ _16219_/A vssd1 vssd1 vccd1 vccd1 _19381_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15079__A _15079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17199_ _17630_/B _12245_/A _17251_/S vssd1 vssd1 vccd1 vccd1 _17199_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11726__A1 _11070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09805__A _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__clkbuf_2
XFILLER_111_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14428__A0 _13918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10450__S _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10701__A2 _09833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17090__A1 _15615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12439__C1 _12230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11492__D _11492_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09524_ _11320_/S vssd1 vssd1 vccd1 vccd1 _10055_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_65_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_141_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19800_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_169_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09950__S0 _10112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09455_ _19327_/Q _18739_/Q _18776_/Q _18350_/Q _10496_/A _09390_/A vssd1 vssd1 vccd1
+ vccd1 _09456_/B sky130_fd_sc_hd__mux4_1
XFILLER_80_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10560__S1 _09443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09386_ _09598_/A vssd1 vssd1 vccd1 vccd1 _11297_/S sky130_fd_sc_hd__buf_2
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18064__S _18066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_156_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19301_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10230_ _18932_/Q _18698_/Q _19380_/Q _19028_/Q _10315_/S _10229_/X vssd1 vssd1 vccd1
+ vccd1 _10231_/B sky130_fd_sc_hd__mux4_2
XFILLER_145_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17853__A0 _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ _19192_/Q _18806_/Q _19256_/Q _18375_/Q _09904_/X _09888_/X vssd1 vssd1 vccd1
+ vccd1 _10162_/B sky130_fd_sc_hd__mux4_1
XFILLER_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10092_ _10148_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__or2_1
XFILLER_120_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13920_ _13920_/A vssd1 vssd1 vccd1 vccd1 _18505_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17081__A1 _12689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13851_ _14531_/A vssd1 vssd1 vccd1 vccd1 _13851_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13671__S _13675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12802_ _19812_/Q vssd1 vssd1 vccd1 vccd1 _16619_/D sky130_fd_sc_hd__buf_6
X_16570_ _16570_/A _16575_/C vssd1 vssd1 vccd1 vccd1 _16570_/Y sky130_fd_sc_hd__nor2_1
X_13782_ _13782_/A vssd1 vssd1 vccd1 vccd1 _18455_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17908__A1 _11512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ _18917_/Q _18683_/Q _19365_/Q _19013_/Q _11050_/S _10934_/A vssd1 vssd1 vccd1
+ vccd1 _10994_/X sky130_fd_sc_hd__mux4_1
XFILLER_76_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_109_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19671_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09450__A _09450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15521_ _15541_/A hold16/A vssd1 vssd1 vccd1 vccd1 _15521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_15_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12733_ _18254_/Q _12732_/X _17520_/S vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__mux2_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__A _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18240_ _18240_/A vssd1 vssd1 vccd1 vccd1 _19863_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15452_ _15452_/A vssd1 vssd1 vccd1 vccd1 _19131_/D sky130_fd_sc_hd__clkbuf_1
X_12664_ _19436_/Q _12636_/X _12663_/X vssd1 vssd1 vccd1 vccd1 _12664_/X sky130_fd_sc_hd__o21a_1
XFILLER_15_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14403_/A vssd1 vssd1 vccd1 vccd1 _18690_/D sky130_fd_sc_hd__clkbuf_1
X_11615_ _12093_/A vssd1 vssd1 vccd1 vccd1 _12078_/A sky130_fd_sc_hd__clkbuf_2
X_18171_ _18171_/A vssd1 vssd1 vccd1 vccd1 _19841_/D sky130_fd_sc_hd__clkbuf_1
X_15383_ _19101_/Q _15092_/X _15383_/S vssd1 vssd1 vccd1 vccd1 _15384_/A sky130_fd_sc_hd__mux2_1
XFILLER_169_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _14275_/A vssd1 vssd1 vccd1 vccd1 _14623_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14334_ _14356_/A vssd1 vssd1 vccd1 vccd1 _14343_/S sky130_fd_sc_hd__buf_4
X_17122_ _17122_/A _17122_/B _17122_/C _17122_/D vssd1 vssd1 vccd1 vccd1 _17122_/X
+ sky130_fd_sc_hd__or4_1
X_11546_ _14272_/A _12672_/A vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__or2_2
XFILLER_129_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17053_ _19674_/Q _15522_/X _17061_/S vssd1 vssd1 vccd1 vccd1 _17054_/A sky130_fd_sc_hd__mux2_1
X_14265_ _14265_/A vssd1 vssd1 vccd1 vccd1 _18638_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ _11432_/X _11433_/Y _11434_/X _11435_/Y _11476_/X vssd1 vssd1 vccd1 vccd1
+ _11477_/X sky130_fd_sc_hd__a221o_1
X_16004_ _15999_/Y _19330_/Q _16025_/S vssd1 vssd1 vccd1 vccd1 _16005_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11220__A _11220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ _19478_/Q vssd1 vssd1 vccd1 vccd1 _16483_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10428_ _19283_/Q _19121_/Q _18530_/Q _18300_/Q _10381_/S _09886_/A vssd1 vssd1 vccd1
+ vccd1 _10429_/B sky130_fd_sc_hd__mux4_1
XFILLER_125_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14196_ _14196_/A vssd1 vssd1 vccd1 vccd1 _18608_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ _15057_/A vssd1 vssd1 vccd1 vccd1 _14579_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10359_ _10237_/X _10358_/X _09727_/A vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16222__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10392__B1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13078_ _16782_/C _12638_/X _13077_/X _12644_/X vssd1 vssd1 vccd1 vccd1 _13078_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17955_ _19752_/Q _19784_/Q _17957_/S vssd1 vssd1 vccd1 vccd1 _17956_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13147__A _15057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16906_ _16914_/A _16906_/B _16906_/C vssd1 vssd1 vccd1 vccd1 _19614_/D sky130_fd_sc_hd__nor3_1
X_12029_ _12031_/A _17211_/A vssd1 vssd1 vccd1 vccd1 _12030_/A sky130_fd_sc_hd__nand2_1
XFILLER_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17886_ _17907_/A _17886_/B vssd1 vssd1 vccd1 vccd1 _17886_/X sky130_fd_sc_hd__or2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17072__A1 _15568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19625_ _19663_/CLK _19625_/D vssd1 vssd1 vccd1 vccd1 _19625_/Q sky130_fd_sc_hd__dfxtp_1
X_16837_ _16836_/A _16836_/B _19590_/Q vssd1 vssd1 vccd1 vccd1 _16838_/C sky130_fd_sc_hd__a21oi_1
XFILLER_65_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13581__S _13593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11890__A _18144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10790__S1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19556_ _19828_/CLK _19556_/D vssd1 vssd1 vccd1 vccd1 _19556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16768_ _16778_/C _16780_/C vssd1 vssd1 vccd1 vccd1 _16770_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18021__A0 _19782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18507_ _19098_/CLK _18507_/D vssd1 vssd1 vccd1 vccd1 _18507_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_13_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ _13525_/X _19205_/Q _15721_/S vssd1 vssd1 vccd1 vccd1 _15720_/A sky130_fd_sc_hd__mux2_1
X_19487_ _19594_/CLK _19487_/D vssd1 vssd1 vccd1 vccd1 _19487_/Q sky130_fd_sc_hd__dfxtp_1
X_16699_ _19542_/Q _16704_/D _16698_/Y vssd1 vssd1 vccd1 vccd1 _19542_/D sky130_fd_sc_hd__o21a_1
X_09240_ _09206_/X _09231_/X _09235_/X _11943_/A _12159_/A vssd1 vssd1 vccd1 vccd1
+ _17133_/A sky130_fd_sc_hd__o2111a_4
X_18438_ _19619_/CLK _18438_/D vssd1 vssd1 vccd1 vccd1 _18438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19471_/CLK sky130_fd_sc_hd__clkbuf_16
X_09171_ _11513_/A _09171_/B vssd1 vssd1 vccd1 vccd1 _11646_/C sky130_fd_sc_hd__nand2_1
X_18369_ _19250_/CLK _18369_/D vssd1 vssd1 vccd1 vccd1 _18369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16193__A _16239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_88_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19607_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12226__A _19412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09999__S0 _09850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13756__S _13758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_11_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19098_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09535__A _10590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12599__C _12606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10686__A1 _10590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10230__S0 _10315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14587__S _14599_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19388_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09507_ _09507_/A vssd1 vssd1 vccd1 vccd1 _10261_/A sky130_fd_sc_hd__buf_2
XFILLER_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _10614_/A vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__clkbuf_2
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16574__B1 _19506_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09369_ _09369_/A vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_138_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15211__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11400_ _11404_/A _11400_/B vssd1 vssd1 vccd1 vccd1 _11400_/Y sky130_fd_sc_hd__nor2_1
X_12380_ _17404_/A _17886_/B _12356_/B vssd1 vssd1 vccd1 vccd1 _12381_/B sky130_fd_sc_hd__a21boi_2
XFILLER_166_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ _11331_/A _11331_/B vssd1 vssd1 vccd1 vccd1 _11331_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10610__A1 _09995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16831__A _16833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14050_ _14050_/A vssd1 vssd1 vccd1 vccd1 _18544_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11262_ _11262_/A _11262_/B vssd1 vssd1 vccd1 vccd1 _11262_/Y sky130_fd_sc_hd__nor2_1
XFILLER_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ _13001_/A vssd1 vssd1 vccd1 vccd1 _18292_/D sky130_fd_sc_hd__clkbuf_1
X_10213_ _18933_/Q _18699_/Q _19381_/Q _19029_/Q _09955_/S _09954_/A vssd1 vssd1 vccd1
+ vccd1 _10214_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11193_ _12444_/B _11284_/A _12445_/B _11192_/Y vssd1 vssd1 vccd1 vccd1 _11464_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_79_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input42_A io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__A _10042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10144_ _18599_/Q _18870_/Q _19094_/Q _18838_/Q _10094_/S _10090_/X vssd1 vssd1 vccd1
+ vccd1 _10144_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12115__A1 _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15881__S _15887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17740_ _17740_/A vssd1 vssd1 vccd1 vccd1 _17740_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14952_ _18922_/Q vssd1 vssd1 vccd1 vccd1 _14953_/A sky130_fd_sc_hd__clkbuf_1
X_10075_ _10684_/A _10072_/X _10074_/X vssd1 vssd1 vccd1 vccd1 _10075_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_87_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13903_ _13902_/X _18500_/Q _13903_/S vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17671_ _10703_/Y _17652_/X _17670_/X vssd1 vssd1 vccd1 vccd1 _19717_/D sky130_fd_sc_hd__a21oi_1
XFILLER_130_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14883_ _14883_/A vssd1 vssd1 vccd1 vccd1 _18889_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19410_ _19802_/CLK _19410_/D vssd1 vssd1 vccd1 vccd1 _19410_/Q sky130_fd_sc_hd__dfxtp_1
X_16622_ _16622_/A _16622_/B _16622_/C _16621_/X vssd1 vssd1 vccd1 vccd1 _16625_/C
+ sky130_fd_sc_hd__or4b_1
X_13834_ _13834_/A vssd1 vssd1 vccd1 vccd1 _18479_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13615__A1 _13614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09180__A _18102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ _19759_/CLK _19341_/D vssd1 vssd1 vccd1 vccd1 _19341_/Q sky130_fd_sc_hd__dfxtp_2
X_16553_ _19498_/Q _19497_/Q _19496_/Q _16553_/D vssd1 vssd1 vccd1 vccd1 _16559_/C
+ sky130_fd_sc_hd__and4_1
X_13765_ _15926_/A _15710_/A vssd1 vssd1 vccd1 vccd1 _13822_/A sky130_fd_sc_hd__nand2_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10977_ _10977_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10977_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_187_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15504_ _15504_/A vssd1 vssd1 vccd1 vccd1 _19145_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12716_ _12715_/X _12696_/X _12716_/S vssd1 vssd1 vccd1 vccd1 _12716_/X sky130_fd_sc_hd__mux2_1
X_19272_ _19272_/CLK _19272_/D vssd1 vssd1 vccd1 vccd1 _19272_/Q sky130_fd_sc_hd__dfxtp_1
X_16484_ _16483_/B _16483_/C _19479_/Q vssd1 vssd1 vccd1 vccd1 _16485_/C sky130_fd_sc_hd__a21oi_1
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13696_ _13696_/A vssd1 vssd1 vccd1 vccd1 _18417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18223_ _18223_/A vssd1 vssd1 vccd1 vccd1 _19858_/D sky130_fd_sc_hd__clkbuf_1
X_12647_ _19531_/Q _12583_/X _12635_/X hold3/A _12646_/X vssd1 vssd1 vccd1 vccd1 _12647_/X
+ sky130_fd_sc_hd__a221o_2
X_15435_ _15446_/A vssd1 vssd1 vccd1 vccd1 _15444_/S sky130_fd_sc_hd__buf_4
XFILLER_157_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15366_ _19093_/Q _15067_/X _15372_/S vssd1 vssd1 vccd1 vccd1 _15367_/A sky130_fd_sc_hd__mux2_1
X_18154_ _18154_/A vssd1 vssd1 vccd1 vccd1 _19836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12578_ _19622_/Q _12556_/X _12498_/Y _12577_/X vssd1 vssd1 vccd1 vccd1 _19622_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17105_ _17105_/A _17117_/B vssd1 vssd1 vccd1 vccd1 _17105_/X sky130_fd_sc_hd__or2_1
X_14317_ _13864_/X _18653_/Q _14321_/S vssd1 vssd1 vccd1 vccd1 _14318_/A sky130_fd_sc_hd__mux2_1
X_11529_ _11525_/A _09158_/A _17114_/C _17122_/C _11559_/A vssd1 vssd1 vccd1 vccd1
+ _17174_/B sky130_fd_sc_hd__a32o_1
X_18085_ _19809_/Q _12627_/X _18083_/X _18084_/X vssd1 vssd1 vccd1 vccd1 _19809_/D
+ sky130_fd_sc_hd__o211a_1
X_15297_ _15297_/A vssd1 vssd1 vccd1 vccd1 _19062_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16741__A _19557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17036_ _17036_/A vssd1 vssd1 vccd1 vccd1 _19666_/D sky130_fd_sc_hd__clkbuf_1
X_14248_ _14248_/A vssd1 vssd1 vccd1 vccd1 _18630_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17048__S _17050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09755__C1 _09754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ _14179_/A vssd1 vssd1 vccd1 vccd1 _18600_/D sky130_fd_sc_hd__clkbuf_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10460__S0 _10499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18987_ _18987_/CLK _18987_/D vssd1 vssd1 vccd1 vccd1 _18987_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15791__S _15793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _16021_/A _19776_/Q _17946_/S vssd1 vssd1 vccd1 vccd1 _17939_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17869_ _17413_/A _17866_/X _17868_/Y _17494_/X vssd1 vssd1 vccd1 vccd1 _17869_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19608_ _19618_/CLK _19608_/D vssd1 vssd1 vccd1 vccd1 _19608_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13605__A _15089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15092__A _15092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19539_ _19540_/CLK _19539_/D vssd1 vssd1 vccd1 vccd1 _19539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09286__A1 _12543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15359__A1 _15057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09223_ _09474_/A _09223_/B _09474_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__or3_1
XFILLER_167_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10840__A1 _19112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09154_ _09154_/A _09211_/A _09211_/B vssd1 vssd1 vccd1 vccd1 _17166_/C sky130_fd_sc_hd__and3_1
XFILLER_147_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_10_0_clock clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__15966__S _15970_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09085_ _17121_/A _17124_/B vssd1 vssd1 vccd1 vccd1 _12482_/B sky130_fd_sc_hd__nor2_8
XFILLER_162_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15531__A1 _12669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13486__S _13492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11795__A _11826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17808__B1 _17807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12896__A2 _12817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ _18411_/Q _18672_/Q _18571_/Q _18906_/Q _09599_/X _09977_/A vssd1 vssd1 vccd1
+ vccd1 _09988_/B sky130_fd_sc_hd__mux4_1
XFILLER_77_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10754__S1 _11298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ _10965_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15206__S _15206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14110__S _14118_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11880_ _11880_/A _11969_/D vssd1 vssd1 vccd1 vccd1 _11880_/Y sky130_fd_sc_hd__nor2_1
XFILLER_72_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10831_ _09596_/A _10828_/X _10830_/X _09448_/A vssd1 vssd1 vccd1 vccd1 _10831_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13073__A2 _12974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13550_ _13550_/A vssd1 vssd1 vccd1 vccd1 _18363_/D sky130_fd_sc_hd__clkbuf_1
X_10762_ _11309_/A _10762_/B vssd1 vssd1 vccd1 vccd1 _10762_/X sky130_fd_sc_hd__or2_1
XFILLER_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12501_ _13260_/A vssd1 vssd1 vccd1 vccd1 _12501_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10831__A1 _09596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13481_ _13171_/X _18340_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _13482_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10693_ _10693_/A _10693_/B vssd1 vssd1 vccd1 vccd1 _10693_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15220_ _19028_/Q _15063_/X _15228_/S vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13250__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12432_ _12432_/A _12432_/B vssd1 vssd1 vccd1 vccd1 _12432_/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _15151_/A vssd1 vssd1 vccd1 vccd1 _18997_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12363_ _12363_/A _12363_/B _12363_/C vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__nand3_1
XFILLER_154_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14102_ _14102_/A vssd1 vssd1 vccd1 vccd1 _18566_/D sky130_fd_sc_hd__clkbuf_1
X_11314_ _19279_/Q _19117_/Q _18526_/Q _18296_/Q _10030_/S _10669_/A vssd1 vssd1 vccd1
+ vccd1 _11314_/X sky130_fd_sc_hd__mux4_1
X_15082_ _15082_/A vssd1 vssd1 vccd1 vccd1 _18969_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15522__B2 hold16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _12294_/A _12339_/C vssd1 vssd1 vccd1 vccd1 _12294_/Y sky130_fd_sc_hd__nor2_1
X_18910_ _19296_/CLK _18910_/D vssd1 vssd1 vccd1 vccd1 _18910_/Q sky130_fd_sc_hd__dfxtp_1
X_14033_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14033_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11245_ _11138_/A _11240_/X _11242_/X _11244_/X vssd1 vssd1 vccd1 vccd1 _11245_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17275__A1 _17662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18841_ _19391_/CLK _18841_/D vssd1 vssd1 vccd1 vccd1 _18841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13409__B _18252_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _18780_/Q vssd1 vssd1 vccd1 vccd1 _11177_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_122_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10127_ _10129_/A _10126_/X _09823_/X vssd1 vssd1 vccd1 vccd1 _10127_/Y sky130_fd_sc_hd__o21ai_1
X_18772_ _19385_/CLK _18772_/D vssd1 vssd1 vccd1 vccd1 _18772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15984_ _13595_/X _19323_/Q _15992_/S vssd1 vssd1 vccd1 vccd1 _15985_/A sky130_fd_sc_hd__mux2_1
X_17723_ _17722_/A _17722_/B _17832_/S vssd1 vssd1 vccd1 vccd1 _17724_/B sky130_fd_sc_hd__mux2_1
X_14935_ _14935_/A vssd1 vssd1 vccd1 vccd1 _18913_/D sky130_fd_sc_hd__clkbuf_1
X_10058_ _10056_/A _10054_/Y _10056_/Y _10689_/A vssd1 vssd1 vccd1 vccd1 _10058_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15589__A1 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17654_ _17654_/A _17654_/B vssd1 vssd1 vccd1 vccd1 _17654_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14866_ _14866_/A vssd1 vssd1 vccd1 vccd1 _18881_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16605_ _16660_/A _16605_/B _16609_/C vssd1 vssd1 vccd1 vccd1 _19515_/D sky130_fd_sc_hd__nor3_1
XFILLER_51_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13817_ _13817_/A vssd1 vssd1 vccd1 vccd1 _18471_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17585_ _17582_/X _17583_/Y _17855_/S vssd1 vssd1 vccd1 vccd1 _17585_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14797_ _18851_/Q _13959_/X _14799_/S vssd1 vssd1 vccd1 vccd1 _14798_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15640__A _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19324_ _19324_/CLK _19324_/D vssd1 vssd1 vccd1 vccd1 _19324_/Q sky130_fd_sc_hd__dfxtp_1
X_16536_ _19492_/Q _16530_/C _16535_/Y vssd1 vssd1 vccd1 vccd1 _19492_/D sky130_fd_sc_hd__o21a_1
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13748_ _13748_/A vssd1 vssd1 vccd1 vccd1 _18441_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11170__S1 _11012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19255_ _19502_/CLK _19255_/D vssd1 vssd1 vccd1 vccd1 _19255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16467_ _16466_/B _16466_/C _19473_/Q vssd1 vssd1 vccd1 vccd1 _16468_/C sky130_fd_sc_hd__a21oi_1
XFILLER_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13679_ _13679_/A vssd1 vssd1 vccd1 vccd1 _18410_/D sky130_fd_sc_hd__clkbuf_1
X_18206_ _18206_/A vssd1 vssd1 vccd1 vccd1 _19850_/D sky130_fd_sc_hd__clkbuf_1
X_15418_ _19116_/Q _15038_/X _15422_/S vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__mux2_1
X_19186_ _19250_/CLK _19186_/D vssd1 vssd1 vccd1 vccd1 _19186_/Q sky130_fd_sc_hd__dfxtp_1
X_16398_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16427_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_163_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10035__C1 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18137_ _19829_/Q _18134_/X _18135_/X _18136_/X vssd1 vssd1 vccd1 vccd1 _19829_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14690__S _14698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15349_ _15349_/A vssd1 vssd1 vccd1 vccd1 _19085_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10050__A2 _10040_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18068_ _09236_/D _19803_/Q _18121_/A vssd1 vssd1 vccd1 vccd1 _18069_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10681__S0 _10566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17019_ _15625_/X _17010_/X _17018_/X _17008_/X vssd1 vssd1 vccd1 vccd1 _19660_/D
+ sky130_fd_sc_hd__o211a_1
X_09910_ _09968_/A _09908_/X _09909_/X vssd1 vssd1 vccd1 vccd1 _09910_/X sky130_fd_sc_hd__o21a_1
XFILLER_144_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09841_ _09866_/A vssd1 vssd1 vccd1 vccd1 _10195_/A sky130_fd_sc_hd__buf_2
XFILLER_98_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09891_/A vssd1 vssd1 vccd1 vccd1 _09773_/A sky130_fd_sc_hd__buf_2
XFILLER_98_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09813__A _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15534__B _15534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17569__A2 _09322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14865__S _14871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09206_ _11567_/A _11678_/A _09205_/X vssd1 vssd1 vccd1 vccd1 _09206_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10026__C1 _09811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ _19864_/Q _19863_/Q _19865_/Q vssd1 vssd1 vccd1 vccd1 _09167_/B sky130_fd_sc_hd__or3b_1
XANTENNA__15696__S _15704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10672__S0 _10729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_135_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10633__S _10633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14105__S _14107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11030_ _11033_/A vssd1 vssd1 vccd1 vccd1 _11030_/X sky130_fd_sc_hd__buf_2
XANTENNA__10424__S0 _10381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17009__A1 _15600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09723__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _14547_/A vssd1 vssd1 vccd1 vccd1 _12981_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10869__A _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10727__S1 _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14525_/X _18817_/Q _14726_/S vssd1 vssd1 vccd1 vccd1 _14721_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _11932_/A vssd1 vssd1 vccd1 vccd1 _11932_/Y sky130_fd_sc_hd__clkinv_4
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ _16963_/A _11886_/C vssd1 vssd1 vccd1 vccd1 _11863_/X sky130_fd_sc_hd__or2_1
XFILLER_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14651_ _14651_/A vssd1 vssd1 vccd1 vccd1 _18786_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14775__S _14781_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _10878_/A vssd1 vssd1 vccd1 vccd1 _11049_/S sky130_fd_sc_hd__buf_4
XANTENNA__11057__A1 _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13602_ _15086_/A vssd1 vssd1 vccd1 vccd1 _13602_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17364_/Y _17369_/X _17615_/A vssd1 vssd1 vccd1 vccd1 _17370_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14582_ _14582_/A vssd1 vssd1 vccd1 vccd1 _14582_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11794_ _11794_/A vssd1 vssd1 vccd1 vccd1 _11794_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_14_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16321_ _19424_/Q _16321_/B _16504_/B vssd1 vssd1 vccd1 vccd1 _16322_/C sky130_fd_sc_hd__and3_1
XFILLER_9_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13533_ _18358_/Q _13531_/X _13545_/S vssd1 vssd1 vccd1 vccd1 _13534_/A sky130_fd_sc_hd__mux2_1
X_10745_ _11305_/A _10744_/X _09448_/A vssd1 vssd1 vccd1 vccd1 _10745_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14076__A _14122_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19040_ _19202_/CLK _19040_/D vssd1 vssd1 vccd1 vccd1 _19040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_158_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16252_ _16252_/A vssd1 vssd1 vccd1 vccd1 _19396_/D sky130_fd_sc_hd__clkbuf_1
X_13464_ _13038_/X _18332_/Q _13470_/S vssd1 vssd1 vccd1 vccd1 _13465_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10676_ _09368_/A _10663_/X _10675_/X _09471_/A _19718_/Q vssd1 vssd1 vccd1 vccd1
+ _10677_/A sky130_fd_sc_hd__a32o_1
XFILLER_167_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12415_ _17020_/A _12416_/B vssd1 vssd1 vccd1 vccd1 _12415_/X sky130_fd_sc_hd__or2_1
X_15203_ _15203_/A vssd1 vssd1 vccd1 vccd1 _19020_/D sky130_fd_sc_hd__clkbuf_1
X_13395_ _11801_/B _18315_/Q _13424_/S vssd1 vssd1 vccd1 vccd1 _13396_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16183_ _13531_/X _19365_/Q _16191_/S vssd1 vssd1 vccd1 vccd1 _16184_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12346_ _19419_/Q _11640_/X _12342_/X _12345_/Y vssd1 vssd1 vccd1 vccd1 _16302_/B
+ sky130_fd_sc_hd__o22a_4
X_15134_ _18990_/Q _15044_/X _15134_/S vssd1 vssd1 vccd1 vccd1 _15135_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09973__A2 _09962_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15065_ _18964_/Q _15063_/X _15077_/S vssd1 vssd1 vccd1 vccd1 _15066_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14015__S _14027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ _17005_/A _12298_/C _12276_/Y vssd1 vssd1 vccd1 vccd1 _12277_/X sky130_fd_sc_hd__o21a_1
XFILLER_114_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14016_ _14016_/A vssd1 vssd1 vccd1 vccd1 _18533_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17248__A1 _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _11228_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11228_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_output73_A _11932_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18824_ _18824_/CLK _18824_/D vssd1 vssd1 vccd1 vccd1 _18824_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11159_ _19173_/Q _18787_/Q _19237_/Q _18356_/Q _10904_/X _11033_/X vssd1 vssd1 vccd1
+ vccd1 _11160_/B sky130_fd_sc_hd__mux4_1
XFILLER_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18755_ _19307_/CLK _18755_/D vssd1 vssd1 vccd1 vccd1 _18755_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15967_ _15967_/A vssd1 vssd1 vccd1 vccd1 _19315_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17706_ _17706_/A vssd1 vssd1 vccd1 vccd1 _19719_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14918_ _18905_/Q _14029_/X _14926_/S vssd1 vssd1 vccd1 vccd1 _14919_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18686_ _19369_/CLK _18686_/D vssd1 vssd1 vccd1 vccd1 _18686_/Q sky130_fd_sc_hd__dfxtp_1
X_15898_ _19285_/Q _14582_/A _15898_/S vssd1 vssd1 vccd1 vccd1 _15899_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17637_ _19715_/Q _17570_/X _17636_/X vssd1 vssd1 vccd1 vccd1 _19715_/D sky130_fd_sc_hd__o21a_1
XFILLER_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14685__S _14687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14849_ _14849_/A vssd1 vssd1 vccd1 vccd1 _18874_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17568_ _11765_/A _17328_/B _09322_/X vssd1 vssd1 vccd1 vccd1 _17568_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19307_ _19307_/CLK _19307_/D vssd1 vssd1 vccd1 vccd1 _19307_/Q sky130_fd_sc_hd__dfxtp_1
X_16519_ _16520_/B _16915_/B _19488_/Q vssd1 vssd1 vccd1 vccd1 _16521_/B sky130_fd_sc_hd__a21oi_1
XFILLER_149_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17499_ _17448_/S _17347_/Y _17498_/Y vssd1 vssd1 vccd1 vccd1 _17499_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_149_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19238_ _19302_/CLK _19238_/D vssd1 vssd1 vccd1 vccd1 _19238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13745__A0 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12218__B _12219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19169_ _19660_/CLK _19169_/D vssd1 vssd1 vccd1 vccd1 _19169_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10019__A _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11646__D_N _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09824_ _11402_/A _09819_/X _09823_/X vssd1 vssd1 vccd1 vccd1 _09824_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_150_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10731__B1 _09596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09755_ _09730_/X _09745_/X _09747_/X _09751_/X _09754_/X vssd1 vssd1 vccd1 vccd1
+ _09755_/X sky130_fd_sc_hd__a311o_1
XFILLER_100_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10689__A _10689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_104_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09686_ _18637_/Q _18972_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__mux2_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17411__A1 _17907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15280__A _15302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_61_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12787__A1 _16731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_168_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10530_ _19185_/Q _18799_/Q _19249_/Q _18368_/Q _10433_/S _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10531_/B sky130_fd_sc_hd__mux4_1
XFILLER_11_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11313__A _11313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10461_ _10461_/A _10461_/B vssd1 vssd1 vccd1 vccd1 _10461_/X sky130_fd_sc_hd__or2_1
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _12200_/A vssd1 vssd1 vccd1 vccd1 _12200_/Y sky130_fd_sc_hd__clkinv_2
X_13180_ _19684_/Q _12659_/X _12680_/X _19651_/Q vssd1 vssd1 vccd1 vccd1 _13180_/X
+ sky130_fd_sc_hd__a22o_1
X_10392_ _10394_/A _10391_/X _09822_/A vssd1 vssd1 vccd1 vccd1 _10392_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_136_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15489__A0 _19712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12131_ _19649_/Q vssd1 vssd1 vccd1 vccd1 _16989_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10565__A3 _10564_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12062_ _12175_/A vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_78_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11013_ _19271_/Q _19109_/Q _18518_/Q _18288_/Q _11011_/X _11012_/X vssd1 vssd1 vccd1
+ vccd1 _11013_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16870_ _16871_/A _16871_/C _16869_/Y vssd1 vssd1 vccd1 vccd1 _19601_/D sky130_fd_sc_hd__o21a_1
XFILLER_104_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15821_ _15821_/A vssd1 vssd1 vccd1 vccd1 _19250_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18540_ _19387_/CLK _18540_/D vssd1 vssd1 vccd1 vccd1 _18540_/Q sky130_fd_sc_hd__dfxtp_1
X_15752_ _13573_/X _19220_/Q _15754_/S vssd1 vssd1 vccd1 vccd1 _15753_/A sky130_fd_sc_hd__mux2_1
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09172__B _18081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12964_ _12957_/X _12959_/X _12961_/X _12962_/X _16351_/B vssd1 vssd1 vccd1 vccd1
+ _12964_/X sky130_fd_sc_hd__o32a_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14703_ _14605_/X _18810_/Q _14709_/S vssd1 vssd1 vccd1 vccd1 _14704_/A sky130_fd_sc_hd__mux2_1
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ _11915_/A _12093_/A vssd1 vssd1 vccd1 vccd1 _11915_/X sky130_fd_sc_hd__or2_1
X_18471_ _19471_/CLK _18471_/D vssd1 vssd1 vccd1 vccd1 _18471_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15683_ _15683_/A vssd1 vssd1 vccd1 vccd1 _19189_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A vssd1 vssd1 vccd1 vccd1 _12895_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17422_ _17422_/A vssd1 vssd1 vccd1 vccd1 _17733_/A sky130_fd_sc_hd__buf_2
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14634_ input43/X _18148_/A _14293_/X _14623_/X _18114_/A vssd1 vssd1 vccd1 vccd1
+ _18211_/B sky130_fd_sc_hd__a32o_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11847_/A _17198_/A vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__and2_1
XFILLER_54_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11125__S1 _11124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13422__B _13422_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17353_ _17206_/X _17197_/X _17356_/S vssd1 vssd1 vccd1 vccd1 _17353_/X sky130_fd_sc_hd__mux2_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11778_/B _11778_/C _16953_/A vssd1 vssd1 vccd1 vccd1 _11777_/Y sky130_fd_sc_hd__o21ai_1
X_14565_ _14565_/A vssd1 vssd1 vccd1 vccd1 _18760_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _18079_/B vssd1 vssd1 vccd1 vccd1 _16914_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_119_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13516_ _13615_/S vssd1 vssd1 vccd1 vccd1 _13529_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_41_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10728_ _10769_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10728_/X sky130_fd_sc_hd__or2_1
X_17284_ _17282_/X _17283_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17284_/X sky130_fd_sc_hd__mux2_1
X_14496_ _13912_/X _18732_/Q _14500_/S vssd1 vssd1 vccd1 vccd1 _14497_/A sky130_fd_sc_hd__mux2_1
X_19023_ _19119_/CLK _19023_/D vssd1 vssd1 vccd1 vccd1 _19023_/Q sky130_fd_sc_hd__dfxtp_1
X_16235_ _13608_/X _19389_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16236_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13447_ _13447_/A vssd1 vssd1 vccd1 vccd1 _18324_/D sky130_fd_sc_hd__clkbuf_1
X_10659_ _10667_/A _10659_/B vssd1 vssd1 vccd1 vccd1 _10659_/X sky130_fd_sc_hd__or2_1
XFILLER_155_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13378_ _19455_/Q _12962_/X _13377_/X vssd1 vssd1 vccd1 vccd1 _13378_/X sky130_fd_sc_hd__o21a_1
XFILLER_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16166_ _12130_/X _16165_/Y _13430_/B vssd1 vssd1 vccd1 vccd1 _16166_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10636__S0 _10022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11753__A2 _11752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ _18982_/Q _15019_/X _15123_/S vssd1 vssd1 vccd1 vccd1 _15118_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ _18138_/A _11516_/X _12302_/X vssd1 vssd1 vccd1 vccd1 _12329_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_173_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16097_ _19758_/Q _16098_/B vssd1 vssd1 vccd1 vccd1 _16107_/C sky130_fd_sc_hd__or2_1
XFILLER_130_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15048_ _15080_/A vssd1 vssd1 vccd1 vccd1 _15061_/S sky130_fd_sc_hd__buf_2
XFILLER_170_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13584__S _13593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12702__A1 _19162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12702__B2 _19352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19856_ _19866_/CLK _19856_/D vssd1 vssd1 vccd1 vccd1 _19856_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11061__S0 _11011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18807_ _19383_/CLK _18807_/D vssd1 vssd1 vccd1 vccd1 _18807_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold13_A hold13/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19787_ _19800_/CLK _19787_/D vssd1 vssd1 vccd1 vccd1 _19787_/Q sky130_fd_sc_hd__dfxtp_1
X_16999_ _15582_/X _16997_/X _16998_/X _16995_/X vssd1 vssd1 vccd1 vccd1 _19652_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09540_ _10855_/A vssd1 vssd1 vccd1 vccd1 _09541_/A sky130_fd_sc_hd__clkbuf_2
X_18738_ _19264_/CLK _18738_/D vssd1 vssd1 vccd1 vccd1 _18738_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10302__A _10303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09471_ _09471_/A vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18669_ _18902_/CLK _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10492__A2 _10478_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14391__A0 _13864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11787__B _17247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09538__A _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__A1 _15499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09807_ _09968_/A vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__buf_2
XFILLER_87_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09738_ _10243_/A vssd1 vssd1 vccd1 vccd1 _09857_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09548__S1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10468__C1 _09753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09669_ _09669_/A vssd1 vssd1 vccd1 vccd1 _09670_/A sky130_fd_sc_hd__buf_4
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11700_ _12974_/A _11700_/B vssd1 vssd1 vccd1 vccd1 _11703_/B sky130_fd_sc_hd__nand2_2
X_12680_ _12680_/A vssd1 vssd1 vccd1 vccd1 _12680_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _19844_/Q _11721_/S _11596_/A _11755_/A vssd1 vssd1 vccd1 vccd1 _11631_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12139__A _17790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14350_ _13912_/X _18668_/Q _14354_/S vssd1 vssd1 vccd1 vccd1 _14351_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11562_ _11562_/A _11562_/B _11562_/C _17169_/A vssd1 vssd1 vccd1 vccd1 _11713_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_128_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13669__S _13675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ _19165_/Q _13179_/X _12566_/X _19355_/Q _13300_/X vssd1 vssd1 vccd1 vccd1
+ _13301_/X sky130_fd_sc_hd__a221o_2
X_10513_ _19281_/Q _19119_/Q _18528_/Q _18298_/Q _09980_/S _10310_/A vssd1 vssd1 vccd1
+ vccd1 _10514_/B sky130_fd_sc_hd__mux4_1
X_14281_ _14281_/A vssd1 vssd1 vccd1 vccd1 _18641_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10882__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11493_ _11412_/A _11492_/D _18100_/A _17117_/A _11491_/B vssd1 vssd1 vccd1 vccd1
+ _11493_/X sky130_fd_sc_hd__a2111o_1
X_16020_ _16020_/A vssd1 vssd1 vccd1 vccd1 _19333_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14382__A0 _13851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13232_ _16126_/A _13233_/B vssd1 vssd1 vccd1 vccd1 _13234_/B sky130_fd_sc_hd__nor2_1
X_10444_ _10297_/X _10437_/X _10439_/Y _10443_/Y _09812_/A vssd1 vssd1 vccd1 vccd1
+ _10444_/X sky130_fd_sc_hd__o311a_4
XANTENNA__09448__A _09448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10093__S _10093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ _19726_/Q _15566_/B _13360_/S vssd1 vssd1 vccd1 vccd1 _13163_/X sky130_fd_sc_hd__mux2_1
X_10375_ _09844_/A _10366_/X _10370_/X _10374_/X _09669_/A vssd1 vssd1 vccd1 vccd1
+ _10375_/X sky130_fd_sc_hd__a311o_4
XFILLER_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12114_ _12143_/S vssd1 vssd1 vccd1 vccd1 _12423_/S sky130_fd_sc_hd__buf_2
XFILLER_123_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13094_ _19754_/Q vssd1 vssd1 vccd1 vccd1 _13095_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_17971_ _16107_/A _19791_/Q _17979_/S vssd1 vssd1 vccd1 vccd1 _17972_/A sky130_fd_sc_hd__mux2_1
XFILLER_151_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output159_A _16298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19710_ _19740_/CLK _19710_/D vssd1 vssd1 vccd1 vccd1 _19710_/Q sky130_fd_sc_hd__dfxtp_4
X_16922_ _16922_/A vssd1 vssd1 vccd1 vccd1 _19624_/D sky130_fd_sc_hd__clkbuf_1
X_12045_ _16114_/A _12043_/Y _12105_/C _11835_/X vssd1 vssd1 vccd1 vccd1 _12045_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_111_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19641_ _19645_/CLK _19641_/D vssd1 vssd1 vccd1 vccd1 _19641_/Q sky130_fd_sc_hd__dfxtp_1
X_16853_ _16854_/A _16854_/C _16852_/Y vssd1 vssd1 vccd1 vccd1 _19595_/D sky130_fd_sc_hd__o21a_1
XFILLER_66_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15804_ _13544_/X _19243_/Q _15804_/S vssd1 vssd1 vccd1 vccd1 _15805_/A sky130_fd_sc_hd__mux2_1
X_19572_ _19668_/CLK _19572_/D vssd1 vssd1 vccd1 vccd1 _19572_/Q sky130_fd_sc_hd__dfxtp_1
X_16784_ _19568_/Q _16788_/D _16783_/Y vssd1 vssd1 vccd1 vccd1 _19568_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13996_ _13996_/A vssd1 vssd1 vccd1 vccd1 _18527_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10459__C1 _09669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18523_ _19370_/CLK _18523_/D vssd1 vssd1 vccd1 vccd1 _18523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15735_ _13547_/X _19212_/Q _15743_/S vssd1 vssd1 vccd1 vccd1 _15736_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12947_ _12947_/A vssd1 vssd1 vccd1 vccd1 _18290_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13433__A _13619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18454_ _19239_/CLK _18454_/D vssd1 vssd1 vccd1 vccd1 _18454_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15666_ _15666_/A vssd1 vssd1 vccd1 vccd1 _19181_/D sky130_fd_sc_hd__clkbuf_1
X_12878_ _19428_/Q _12700_/X _12877_/X vssd1 vssd1 vccd1 vccd1 _12878_/X sky130_fd_sc_hd__o21a_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17584_/A vssd1 vssd1 vccd1 vccd1 _17844_/S sky130_fd_sc_hd__buf_2
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14617_ _14617_/A vssd1 vssd1 vccd1 vccd1 _14617_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11829_ _19335_/Q _11766_/X _11734_/X _11828_/X _11691_/X vssd1 vssd1 vccd1 vccd1
+ _11829_/X sky130_fd_sc_hd__o221a_1
X_18385_ _19203_/CLK _18385_/D vssd1 vssd1 vccd1 vccd1 _18385_/Q sky130_fd_sc_hd__dfxtp_1
X_15597_ _15597_/A vssd1 vssd1 vccd1 vccd1 _19162_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09616__B2 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12620__A0 _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__A2 _10212_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17336_ _17336_/A vssd1 vssd1 vccd1 vccd1 _17372_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14548_ _14547_/X _18755_/Q _14551_/S vssd1 vssd1 vccd1 vccd1 _14549_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17267_ _17264_/X _17265_/X _17375_/S vssd1 vssd1 vccd1 vccd1 _17267_/X sky130_fd_sc_hd__mux2_1
X_14479_ _14479_/A vssd1 vssd1 vccd1 vccd1 _18724_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19006_ _19006_/CLK _19006_/D vssd1 vssd1 vccd1 vccd1 _19006_/Q sky130_fd_sc_hd__dfxtp_1
X_16218_ _13583_/X _19381_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16219_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09358__A _12751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17198_ _17198_/A vssd1 vssd1 vccd1 vccd1 _17630_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__18103__A2 _18086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11099__S _11265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16149_ _19767_/Q _16150_/B vssd1 vssd1 vccd1 vccd1 _16159_/C sky130_fd_sc_hd__or2_1
XFILLER_170_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17862__A1 _12291_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15095__A _15095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13608__A _15092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14203__S _14209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19839_ _19846_/CLK _19839_/D vssd1 vssd1 vccd1 vccd1 _19839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16919__A _16919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09821__A _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09523_ _10579_/A vssd1 vssd1 vccd1 vccd1 _11320_/S sky130_fd_sc_hd__buf_2
XFILLER_71_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09454_ _10514_/A _09454_/B vssd1 vssd1 vccd1 vccd1 _09454_/X sky130_fd_sc_hd__or2_1
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09385_ _09396_/A vssd1 vssd1 vccd1 vccd1 _09598_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16105__A1 _19348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17485__A _17485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10160_ _09890_/A _10159_/X _09909_/X vssd1 vssd1 vccd1 vccd1 _10160_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17853__A1 _17856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15209__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11025__S0 _10969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10091_ _18935_/Q _18701_/Q _19383_/Q _19031_/Q _10094_/S _10090_/X vssd1 vssd1 vccd1
+ vccd1 _10092_/B sky130_fd_sc_hd__mux4_1
XFILLER_126_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12422__A _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15616__A0 _19734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13850_ _13850_/A vssd1 vssd1 vccd1 vccd1 _18483_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ _14519_/A vssd1 vssd1 vccd1 vccd1 _12801_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__15631__A3 _09234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13781_ _12924_/X _18455_/Q _13787_/S vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__mux2_1
X_10993_ _11242_/A _10992_/X _11257_/A vssd1 vssd1 vccd1 vccd1 _10993_/X sky130_fd_sc_hd__a21o_1
XFILLER_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15520_ hold16/A _15520_/B vssd1 vssd1 vccd1 vccd1 _15520_/X sky130_fd_sc_hd__or2_1
XFILLER_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18030__A1 _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _18114_/A _11677_/X _12735_/S vssd1 vssd1 vccd1 vccd1 _12732_/X sky130_fd_sc_hd__mux2_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10596__B _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15879__S _15887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _19131_/Q _15086_/X _15455_/S vssd1 vssd1 vccd1 vccd1 _15452_/A sky130_fd_sc_hd__mux2_1
X_12663_ _16778_/C _12638_/X _12662_/X _12644_/X vssd1 vssd1 vccd1 vccd1 _12663_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14783__S _14785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _13880_/X _18690_/Q _14406_/S vssd1 vssd1 vccd1 vccd1 _14403_/A sky130_fd_sc_hd__mux2_1
X_11614_ _11887_/A vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18170_ _18170_/A _18170_/B vssd1 vssd1 vccd1 vccd1 _18171_/A sky130_fd_sc_hd__and2_1
X_15382_ _15382_/A vssd1 vssd1 vccd1 vccd1 _19100_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12594_ _19621_/Q _12556_/X _12498_/Y _12593_/X vssd1 vssd1 vccd1 vccd1 _19621_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_129_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17121_ _17121_/A _17121_/B vssd1 vssd1 vccd1 vccd1 _17122_/D sky130_fd_sc_hd__nor2_1
X_14333_ _14333_/A vssd1 vssd1 vccd1 vccd1 _18660_/D sky130_fd_sc_hd__clkbuf_1
X_11545_ input66/X vssd1 vssd1 vccd1 vccd1 _14272_/A sky130_fd_sc_hd__clkinv_2
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11501__A _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__B2 _19347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17052_ _17098_/S vssd1 vssd1 vccd1 vccd1 _17061_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__09178__A _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11476_ _11436_/X _11437_/Y _11438_/X _11439_/Y _11475_/X vssd1 vssd1 vccd1 vccd1
+ _11476_/X sky130_fd_sc_hd__a221o_1
X_14264_ _18638_/Q _14042_/X _14264_/S vssd1 vssd1 vccd1 vccd1 _14265_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16003_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16025_/S sky130_fd_sc_hd__buf_2
XFILLER_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12905__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ _19610_/Q vssd1 vssd1 vccd1 vccd1 _16896_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10427_ _10471_/A _10426_/X _09821_/A vssd1 vssd1 vccd1 vccd1 _10427_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12905__B2 _12798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14195_ _18608_/Q _14048_/X _14195_/S vssd1 vssd1 vccd1 vccd1 _14196_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14107__A0 _13918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14812__A _14858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_183_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _19316_/Q _18728_/Q _18765_/Q _18339_/Q _09700_/A _10238_/X vssd1 vssd1 vccd1
+ vccd1 _10358_/X sky130_fd_sc_hd__mux4_2
X_13146_ _13051_/X _13144_/X _13145_/X vssd1 vssd1 vccd1 vccd1 _15057_/A sky130_fd_sc_hd__o21a_4
XANTENNA__10392__A1 _10394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _19152_/Q _12895_/X _12677_/X _19342_/Q _13076_/X vssd1 vssd1 vccd1 vccd1
+ _13077_/X sky130_fd_sc_hd__a221o_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17954_ _17954_/A vssd1 vssd1 vccd1 vccd1 _19751_/D sky130_fd_sc_hd__clkbuf_1
X_10289_ _10289_/A vssd1 vssd1 vccd1 vccd1 _10535_/A sky130_fd_sc_hd__buf_2
XANTENNA__12332__A _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16905_ _16904_/A _16904_/C _19614_/Q vssd1 vssd1 vccd1 vccd1 _16906_/C sky130_fd_sc_hd__a21oi_1
X_12028_ _19786_/Q _11347_/A _12028_/S vssd1 vssd1 vccd1 vccd1 _17211_/A sky130_fd_sc_hd__mux2_2
XFILLER_111_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17885_ _17886_/B _17885_/B vssd1 vssd1 vccd1 vccd1 _17889_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16739__A _16762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13862__S _13871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19624_ _19671_/CLK _19624_/D vssd1 vssd1 vccd1 vccd1 _19624_/Q sky130_fd_sc_hd__dfxtp_1
X_16836_ _16836_/A _16836_/B _19590_/Q vssd1 vssd1 vccd1 vccd1 _16838_/B sky130_fd_sc_hd__and3_1
XFILLER_38_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19085_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_66_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19555_ _19828_/CLK _19555_/D vssd1 vssd1 vccd1 vccd1 _19555_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11890__B _11890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16767_ _19563_/Q _19562_/Q _16767_/C vssd1 vssd1 vccd1 vccd1 _16780_/C sky130_fd_sc_hd__and3_1
XFILLER_47_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13979_ _18522_/Q _13978_/X _13979_/S vssd1 vssd1 vccd1 vccd1 _13980_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18021__A1 _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18506_ _19385_/CLK _18506_/D vssd1 vssd1 vccd1 vccd1 _18506_/Q sky130_fd_sc_hd__dfxtp_1
X_15718_ _15718_/A vssd1 vssd1 vccd1 vccd1 _19204_/D sky130_fd_sc_hd__clkbuf_1
X_19486_ _19491_/CLK _19486_/D vssd1 vssd1 vccd1 vccd1 _19486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16698_ _16707_/A _16706_/D vssd1 vssd1 vccd1 vccd1 _16698_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18437_ _19287_/CLK _18437_/D vssd1 vssd1 vccd1 vccd1 _18437_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15789__S _15793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15649_ _14534_/X _19174_/Q _15649_/S vssd1 vssd1 vccd1 vccd1 _15650_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09170_ _09186_/A vssd1 vssd1 vccd1 vccd1 _11513_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18368_ _19249_/CLK _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17319_ _17404_/A _17319_/B _17319_/C vssd1 vssd1 vccd1 vccd1 _17659_/A sky130_fd_sc_hd__and3_1
XANTENNA__11947__A2 _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18299_ _19314_/CLK _18299_/D vssd1 vssd1 vccd1 vccd1 _18299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14346__A0 _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__A _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12226__B _19413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18088__A1 _14787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11255__S0 _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10027__A _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09999__S1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16099__B1 _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12242__A _17305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13772__S _13776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15553__A _15603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10230__S1 _10229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A1 _19337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09506_ _09506_/A vssd1 vssd1 vccd1 vccd1 _09507_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__18012__A1 _19399_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11635__A1 _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09437_ _10743_/A vssd1 vssd1 vccd1 vccd1 _10614_/A sky130_fd_sc_hd__clkbuf_4
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09368_ _09368_/A vssd1 vssd1 vccd1 vccd1 _09369_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09299_ _09284_/X _09292_/Y _11805_/C _11698_/B _19697_/Q vssd1 vssd1 vccd1 vccd1
+ _09299_/X sky130_fd_sc_hd__a2111o_1
XFILLER_138_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11330_ _19183_/Q _18797_/Q _19247_/Q _18366_/Q _10692_/S _09628_/X vssd1 vssd1 vccd1
+ vccd1 _11331_/B sky130_fd_sc_hd__mux4_2
XANTENNA__11321__A _11321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11261_ _18912_/Q _18678_/Q _19360_/Q _19008_/Q _10962_/S _11220_/A vssd1 vssd1 vccd1
+ vccd1 _11262_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11246__S0 _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18104__A _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10212_ _10205_/Y _10207_/Y _10209_/Y _10211_/Y _09831_/A vssd1 vssd1 vccd1 vccd1
+ _10212_/X sky130_fd_sc_hd__o221a_2
XFILLER_122_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13000_ _12999_/X _18292_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _13001_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09726__A _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _09367_/A _11182_/X _11191_/X _09470_/A _19710_/Q vssd1 vssd1 vccd1 vccd1
+ _11192_/Y sky130_fd_sc_hd__a32oi_2
XFILLER_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10143_ _10148_/A _10143_/B vssd1 vssd1 vccd1 vccd1 _10143_/X sky130_fd_sc_hd__or2_1
XFILLER_43_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input35_A io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _10074_/A vssd1 vssd1 vccd1 vccd1 _10074_/X sky130_fd_sc_hd__clkbuf_4
X_14951_ _14951_/A vssd1 vssd1 vccd1 vccd1 _18921_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17662__B _17662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13682__S _13686_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ _14582_/A vssd1 vssd1 vccd1 vccd1 _13902_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17670_ _11904_/A _17328_/B _17669_/X _17831_/A vssd1 vssd1 vccd1 vccd1 _17670_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_75_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14882_ _18889_/Q _13978_/X _14882_/S vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__mux2_1
X_16621_ _19809_/Q _19807_/Q _19804_/Q _19803_/Q vssd1 vssd1 vccd1 vccd1 _16621_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09461__A _10042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13833_ _13367_/X _18479_/Q _13835_/S vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13076__B1 _12704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19340_ _19356_/CLK _19340_/D vssd1 vssd1 vccd1 vccd1 _19340_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18003__A1 _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16552_ _16585_/A _16552_/B _16552_/C vssd1 vssd1 vccd1 vccd1 _19497_/D sky130_fd_sc_hd__nor3_1
XFILLER_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13764_ _13947_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _15710_/A sky130_fd_sc_hd__nor2_2
XANTENNA__10400__A _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16014__A0 _15481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10976_ _19176_/Q _18790_/Q _19240_/Q _18359_/Q _10862_/X _09513_/A vssd1 vssd1 vccd1
+ vccd1 _10977_/B sky130_fd_sc_hd__mux4_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15503_ _15502_/X _19145_/Q _15517_/S vssd1 vssd1 vccd1 vccd1 _15504_/A sky130_fd_sc_hd__mux2_1
X_12715_ _12544_/X _12712_/X _12713_/Y _15549_/A _18275_/Q vssd1 vssd1 vccd1 vccd1
+ _12715_/X sky130_fd_sc_hd__a32o_4
X_19271_ _19271_/CLK _19271_/D vssd1 vssd1 vccd1 vccd1 _19271_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16483_ _19479_/Q _16483_/B _16483_/C vssd1 vssd1 vccd1 vccd1 _16485_/B sky130_fd_sc_hd__and3_1
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13695_ _12801_/X _18417_/Q _13703_/S vssd1 vssd1 vccd1 vccd1 _13696_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13379__A1 _19551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18222_ _18224_/A _18222_/B vssd1 vssd1 vccd1 vccd1 _18223_/A sky130_fd_sc_hd__and2_1
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15434_ _15434_/A vssd1 vssd1 vccd1 vccd1 _19123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12646_ _19435_/Q _12636_/X _12645_/X vssd1 vssd1 vccd1 vccd1 _12646_/X sky130_fd_sc_hd__o21a_1
XFILLER_169_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13430__B _13430_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18153_ _18163_/A _18153_/B vssd1 vssd1 vccd1 vccd1 _18154_/A sky130_fd_sc_hd__or2_1
XFILLER_50_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15365_ _15365_/A vssd1 vssd1 vccd1 vccd1 _19092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10546__S _10546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ _17026_/S _12577_/B vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__and2_1
XANTENNA__14018__S _14027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17104_ _19696_/Q _12674_/A _18091_/B _11557_/D _17142_/A vssd1 vssd1 vccd1 vccd1
+ _19696_/D sky130_fd_sc_hd__o221a_1
X_14316_ _14316_/A vssd1 vssd1 vccd1 vccd1 _18652_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18084_ _18097_/A vssd1 vssd1 vccd1 vccd1 _18084_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_117_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _11528_/A _11528_/B _11528_/C vssd1 vssd1 vccd1 vccd1 _17122_/C sky130_fd_sc_hd__and3_2
X_15296_ _14592_/X _19062_/Q _15300_/S vssd1 vssd1 vccd1 vccd1 _15297_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16741__B _16752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17035_ _19666_/Q _13418_/B _17039_/S vssd1 vssd1 vccd1 vccd1 _17036_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14247_ _18630_/Q _14017_/X _14253_/S vssd1 vssd1 vccd1 vccd1 _14248_/A sky130_fd_sc_hd__mux2_1
X_11459_ _11462_/A _11459_/B vssd1 vssd1 vccd1 vccd1 _11460_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16233__S _16235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12354__A2 _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ _18600_/Q _14023_/X _14180_/S vssd1 vssd1 vccd1 vccd1 _14179_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_140_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19786_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_125_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ _16091_/A _13127_/B _13113_/C vssd1 vssd1 vccd1 vccd1 _13130_/B sky130_fd_sc_hd__o21ai_1
XFILLER_140_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _19006_/CLK _18986_/D vssd1 vssd1 vccd1 vccd1 _18986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14500__A0 _13918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _17937_/A vssd1 vssd1 vccd1 vccd1 _17946_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_155_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19302_/CLK sky130_fd_sc_hd__clkbuf_16
X_17868_ _17490_/X _17865_/Y _17867_/Y vssd1 vssd1 vccd1 vccd1 _17868_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_27_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19607_ _19607_/CLK _19607_/D vssd1 vssd1 vccd1 vccd1 _19607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ hold22/A _16821_/C _16818_/X vssd1 vssd1 vccd1 vccd1 _19579_/D sky130_fd_sc_hd__o21ba_1
XANTENNA__16619__D _16619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17799_ _17802_/A _17802_/B vssd1 vssd1 vccd1 vccd1 _17800_/B sky130_fd_sc_hd__and2_1
XFILLER_93_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19538_ _19540_/CLK _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10310__A _10310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09286__A2 _13400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19469_ _19471_/CLK _19469_/D vssd1 vssd1 vccd1 vccd1 _19469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14717__A _14785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ _19859_/Q _13619_/A _13944_/A _09331_/A _09221_/X vssd1 vssd1 vccd1 vccd1
+ _09474_/B sky130_fd_sc_hd__a221o_1
XANTENNA__13621__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09153_ _11528_/A _11528_/B _09176_/B vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__and3_1
XANTENNA__12042__A1 _19343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16932__A _16932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09084_ _09174_/A _19847_/Q vssd1 vssd1 vccd1 vccd1 _17124_/B sky130_fd_sc_hd__or2_4
XFILLER_135_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_174_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13542__A1 _13541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_108_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19830_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_122_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09546__A _10680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09986_ _10769_/A vssd1 vssd1 vccd1 vccd1 _10612_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09980__S _09980_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13058__B1 _13057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11069__C1 _09465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_131_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ _10951_/A _10830_/B vssd1 vssd1 vccd1 vccd1 _10830_/X sky130_fd_sc_hd__or2_1
XFILLER_44_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10761_ _18921_/Q _18687_/Q _19369_/Q _19017_/Q _10660_/X _10655_/X vssd1 vssd1 vccd1
+ vccd1 _10762_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15222__S _15228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10292__B1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12500_ _12697_/A vssd1 vssd1 vccd1 vccd1 _13260_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__13531__A _15015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13480_ _13480_/A vssd1 vssd1 vccd1 vccd1 _18339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10692_ _18620_/Q _18955_/Q _10692_/S vssd1 vssd1 vccd1 vccd1 _10693_/B sky130_fd_sc_hd__mux2_1
XFILLER_139_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ _12430_/A _12430_/B _12430_/C vssd1 vssd1 vccd1 vccd1 _12432_/B sky130_fd_sc_hd__a21o_2
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10044__B1 _09434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15150_ _18997_/Q _15067_/X _15156_/S vssd1 vssd1 vccd1 vccd1 _15151_/A sky130_fd_sc_hd__mux2_1
X_12362_ _12363_/A _12363_/B _12363_/C vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__a21o_1
XFILLER_165_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14101_ _13909_/X _18566_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _14102_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11313_ _11313_/A _11313_/B vssd1 vssd1 vccd1 vccd1 _11313_/X sky130_fd_sc_hd__or2_1
X_15081_ _18969_/Q _15079_/X _15093_/S vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__mux2_1
X_12293_ _19417_/Q _12293_/B vssd1 vssd1 vccd1 vccd1 _12339_/C sky130_fd_sc_hd__and2_1
XFILLER_153_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13533__A1 _13531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ _11005_/X _11243_/X _11257_/A vssd1 vssd1 vccd1 vccd1 _11244_/X sky130_fd_sc_hd__a21o_1
X_14032_ _14032_/A vssd1 vssd1 vccd1 vccd1 _18538_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_56_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15892__S _15898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11197__S _11241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18840_ _19384_/CLK _18840_/D vssd1 vssd1 vccd1 vccd1 _18840_/Q sky130_fd_sc_hd__dfxtp_1
X_11175_ _09394_/A _11172_/X _11174_/X _11188_/A vssd1 vssd1 vccd1 vccd1 _11175_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_72_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19320_/CLK sky130_fd_sc_hd__clkbuf_16
X_10126_ _19321_/Q _18733_/Q _18770_/Q _18344_/Q _09918_/X _09900_/A vssd1 vssd1 vccd1
+ vccd1 _10126_/X sky130_fd_sc_hd__mux4_1
X_18771_ _19384_/CLK _18771_/D vssd1 vssd1 vccd1 vccd1 _18771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15983_ _15983_/A vssd1 vssd1 vccd1 vccd1 _15992_/S sky130_fd_sc_hd__buf_4
XFILLER_79_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17722_ _17722_/A _17722_/B vssd1 vssd1 vccd1 vccd1 _17726_/C sky130_fd_sc_hd__and2_1
X_14934_ _18913_/Q vssd1 vssd1 vccd1 vccd1 _14935_/A sky130_fd_sc_hd__clkbuf_1
X_10057_ _10721_/A vssd1 vssd1 vccd1 vccd1 _10689_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_76_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17653_ _17653_/A _17653_/B vssd1 vssd1 vccd1 vccd1 _17653_/X sky130_fd_sc_hd__or2_1
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14865_ _18881_/Q _13953_/X _14871_/S vssd1 vssd1 vccd1 vccd1 _14866_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_87_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19594_/CLK sky130_fd_sc_hd__clkbuf_16
X_16604_ _19515_/Q _19514_/Q _16604_/C vssd1 vssd1 vccd1 vccd1 _16609_/C sky130_fd_sc_hd__and3_1
X_13816_ _13228_/X _18471_/Q _13820_/S vssd1 vssd1 vccd1 vccd1 _13817_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17584_ _17584_/A vssd1 vssd1 vccd1 vccd1 _17855_/S sky130_fd_sc_hd__clkbuf_2
X_14796_ _14796_/A vssd1 vssd1 vccd1 vccd1 _18850_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16736__B _16736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19323_ _19385_/CLK _19323_/D vssd1 vssd1 vccd1 vccd1 _19323_/Q sky130_fd_sc_hd__dfxtp_1
X_16535_ _16570_/A _16540_/C vssd1 vssd1 vccd1 vccd1 _16535_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16538__A1 _16540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ _13251_/X _18441_/Q _13747_/S vssd1 vssd1 vccd1 vccd1 _13748_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17735__A0 _19721_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10959_ _09367_/A _10949_/X _10958_/X _09470_/A _19713_/Q vssd1 vssd1 vccd1 vccd1
+ _11288_/A sky130_fd_sc_hd__a32o_2
X_19254_ _19380_/CLK _19254_/D vssd1 vssd1 vccd1 vccd1 _19254_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_10_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19086_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16466_ _19473_/Q _16466_/B _16466_/C vssd1 vssd1 vccd1 vccd1 _16468_/B sky130_fd_sc_hd__and3_1
X_13678_ _13274_/X _18410_/Q _13686_/S vssd1 vssd1 vccd1 vccd1 _13679_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_opt_3_0_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18205_ _18213_/A _18205_/B vssd1 vssd1 vccd1 vccd1 _18206_/A sky130_fd_sc_hd__and2_1
XFILLER_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15417_ _15417_/A vssd1 vssd1 vccd1 vccd1 _19115_/D sky130_fd_sc_hd__clkbuf_1
X_12629_ _16245_/A vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__buf_2
X_19185_ _19249_/CLK _19185_/D vssd1 vssd1 vccd1 vccd1 _19185_/Q sky130_fd_sc_hd__dfxtp_1
X_16397_ _16442_/A _16397_/B _16399_/B vssd1 vssd1 vccd1 vccd1 _19448_/D sky130_fd_sc_hd__nor3_1
XFILLER_157_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18136_ _18136_/A vssd1 vssd1 vccd1 vccd1 _18136_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15348_ _19085_/Q _15041_/X _15350_/S vssd1 vssd1 vccd1 vccd1 _15349_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11783__B1 _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19326_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13587__S _13593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18067_ _18067_/A vssd1 vssd1 vccd1 vccd1 _19802_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14272__A _14272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15279_ _15279_/A vssd1 vssd1 vccd1 vccd1 _19054_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10050__A3 _10049_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17018_ _19660_/Q _17024_/B vssd1 vssd1 vccd1 vccd1 _17018_/X sky130_fd_sc_hd__or2_1
XFILLER_99_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09366__A _09366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09840_ _18506_/Q _19001_/Q _09840_/S vssd1 vssd1 vccd1 vccd1 _09840_/X sky130_fd_sc_hd__mux2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _10382_/A vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__buf_2
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _19385_/CLK _18969_/D vssd1 vssd1 vccd1 vccd1 _18969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15307__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12520__A _13009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11838__B2 _19863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10040__A _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14447__A _14515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15042__S _15045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15977__S _15981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09205_ _09341_/A _09193_/X _09198_/X _09204_/X vssd1 vssd1 vccd1 vccd1 _09205_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_147_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09136_ _19848_/Q _19849_/Q vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__or2b_1
XFILLER_163_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13497__S _13503_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10672__S1 _10655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09276__A _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10329__B2 _19726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clock clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09969_ _19290_/Q _19128_/Q _18537_/Q _18307_/Q _10168_/S _10218_/A vssd1 vssd1 vccd1
+ vccd1 _09969_/X sky130_fd_sc_hd__mux4_1
XANTENNA__15217__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11829__A1 _19335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ _15025_/A vssd1 vssd1 vccd1 vccd1 _14547_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10869__B _12453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _11931_/A _11931_/B vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__xor2_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13960__S _13963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14528_/X _18786_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14651_/A sky130_fd_sc_hd__mux2_1
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11862_ _19639_/Q vssd1 vssd1 vccd1 vccd1 _16963_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13601_ _13601_/A vssd1 vssd1 vccd1 vccd1 _18379_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10813_ _11011_/A vssd1 vssd1 vccd1 vccd1 _10878_/A sky130_fd_sc_hd__buf_2
XANTENNA__12254__A1 _12252_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14581_ _14581_/A vssd1 vssd1 vccd1 vccd1 _18765_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _12093_/A vssd1 vssd1 vccd1 vccd1 _11793_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16320_ _16321_/B _16504_/B _19424_/Q vssd1 vssd1 vccd1 vccd1 _16322_/B sky130_fd_sc_hd__a21oi_1
X_13532_ _13615_/S vssd1 vssd1 vccd1 vccd1 _13545_/S sky130_fd_sc_hd__buf_2
XFILLER_159_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10744_ _19276_/Q _19114_/Q _18523_/Q _18293_/Q _10654_/A _09442_/A vssd1 vssd1 vccd1
+ vccd1 _10744_/X sky130_fd_sc_hd__mux4_1
XFILLER_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10360__S0 _09700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16251_ _16255_/A _16251_/B vssd1 vssd1 vccd1 vccd1 _16252_/A sky130_fd_sc_hd__or2_1
XANTENNA__15887__S _15887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ _13463_/A vssd1 vssd1 vccd1 vccd1 _18331_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14791__S _14799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10675_ _09989_/X _10665_/X _10667_/X _09374_/A _10674_/X vssd1 vssd1 vccd1 vccd1
+ _10675_/X sky130_fd_sc_hd__a311o_4
X_15202_ _19020_/Q _15038_/X _15206_/S vssd1 vssd1 vccd1 vccd1 _15203_/A sky130_fd_sc_hd__mux2_1
X_12414_ _19661_/Q vssd1 vssd1 vccd1 vccd1 _17020_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_127_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16182_ _16239_/S vssd1 vssd1 vccd1 vccd1 _16191_/S sky130_fd_sc_hd__buf_2
X_13394_ _13431_/S vssd1 vssd1 vccd1 vccd1 _13424_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_127_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15133_ _15133_/A vssd1 vssd1 vccd1 vccd1 _18989_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12345_ _12394_/C _12344_/Y _11665_/X vssd1 vssd1 vccd1 vccd1 _12345_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10824__S _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09973__A3 _09971_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15064_ _15080_/A vssd1 vssd1 vccd1 vccd1 _15077_/S sky130_fd_sc_hd__buf_4
XFILLER_153_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12276_ _17005_/A _12298_/C _15632_/S vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_107_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14015_ _18533_/Q _14013_/X _14027_/S vssd1 vssd1 vccd1 vccd1 _14016_/A sky130_fd_sc_hd__mux2_1
X_11227_ _19171_/Q _18785_/Q _19235_/Q _18354_/Q _11074_/S _10971_/A vssd1 vssd1 vccd1
+ vccd1 _11228_/B sky130_fd_sc_hd__mux4_2
XFILLER_96_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09914__A _10174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18823_ _19271_/CLK _18823_/D vssd1 vssd1 vccd1 vccd1 _18823_/Q sky130_fd_sc_hd__dfxtp_1
X_11158_ _10915_/X _11153_/X _11155_/Y _11157_/Y _09553_/A vssd1 vssd1 vccd1 vccd1
+ _11158_/X sky130_fd_sc_hd__o221a_1
XFILLER_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _09732_/A _10106_/X _10108_/X _09740_/X vssd1 vssd1 vccd1 vccd1 _10109_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13436__A _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15966_ _13570_/X _19315_/Q _15970_/S vssd1 vssd1 vccd1 vccd1 _15967_/A sky130_fd_sc_hd__mux2_1
X_18754_ _19305_/CLK _18754_/D vssd1 vssd1 vccd1 vccd1 _18754_/Q sky130_fd_sc_hd__dfxtp_1
X_11089_ _11160_/A _11089_/B vssd1 vssd1 vccd1 vccd1 _11089_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14031__S _14043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17705_ _19719_/Q _17704_/X _17873_/S vssd1 vssd1 vccd1 vccd1 _17706_/A sky130_fd_sc_hd__mux2_1
X_14917_ _14917_/A vssd1 vssd1 vccd1 vccd1 _14926_/S sky130_fd_sc_hd__buf_4
XFILLER_76_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15897_ _15897_/A vssd1 vssd1 vccd1 vccd1 _19284_/D sky130_fd_sc_hd__clkbuf_1
X_18685_ _19365_/CLK _18685_/D vssd1 vssd1 vccd1 vccd1 _18685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15651__A _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17636_ _11855_/Y _17427_/X _17635_/X _09359_/X vssd1 vssd1 vccd1 vccd1 _17636_/X
+ sky130_fd_sc_hd__a211o_1
X_14848_ _18874_/Q _14033_/X _14854_/S vssd1 vssd1 vccd1 vccd1 _14849_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15431__A1 _15057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17567_ _17434_/X _17555_/X _17566_/X _17473_/X vssd1 vssd1 vccd1 vccd1 _17567_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10795__A _19716_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14779_ _14611_/X _18844_/Q _14781_/S vssd1 vssd1 vccd1 vccd1 _14780_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16518_ _16522_/D vssd1 vssd1 vccd1 vccd1 _16915_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10256__B1 _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19306_ _19306_/CLK _19306_/D vssd1 vssd1 vccd1 vccd1 _19306_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_143_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17498_ _17511_/S _17498_/B vssd1 vssd1 vccd1 vccd1 _17498_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09661__A2 _09642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16449_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19237_ _19237_/CLK _19237_/D vssd1 vssd1 vccd1 vccd1 _19237_/Q sky130_fd_sc_hd__dfxtp_1
X_19168_ _19694_/CLK _19168_/D vssd1 vssd1 vccd1 vccd1 _19168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11756__B1 _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18119_ _09351_/A _18091_/B _18118_/Y _18110_/X vssd1 vssd1 vccd1 vccd1 _19823_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19099_ _19387_/CLK _19099_/D vssd1 vssd1 vccd1 vccd1 _19099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09823_ _09823_/A vssd1 vssd1 vccd1 vccd1 _09823_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17644__C1 _17532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10731__A1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09754_ _09754_/A vssd1 vssd1 vccd1 vccd1 _09754_/X sky130_fd_sc_hd__buf_2
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14876__S _14882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ _10093_/S vssd1 vssd1 vccd1 vccd1 _11375_/S sky130_fd_sc_hd__buf_2
XFILLER_104_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12236__A1 _12233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10460_ _19186_/Q _18800_/Q _19250_/Q _18369_/Q _10499_/S _10311_/A vssd1 vssd1 vccd1
+ vccd1 _10461_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ _17120_/B _17120_/C _17120_/D vssd1 vssd1 vccd1 vccd1 _09120_/A sky130_fd_sc_hd__and3_1
XFILLER_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10391_ _19316_/Q _18728_/Q _18765_/Q _18339_/Q _10260_/X _10436_/A vssd1 vssd1 vccd1
+ vccd1 _10391_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14116__S _14118_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15489__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12130_ _16162_/S vssd1 vssd1 vccd1 vccd1 _12130_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_163_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12144__B _17222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12061_ _19408_/Q vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__buf_2
XANTENNA__18112__A _18112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16438__B1 _16402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11012_ _11012_/A vssd1 vssd1 vccd1 vccd1 _11012_/X sky130_fd_sc_hd__buf_2
XANTENNA__11514__A3 _17112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15820_ _13567_/X _19250_/Q _15826_/S vssd1 vssd1 vccd1 vccd1 _15821_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15751_/A vssd1 vssd1 vccd1 vccd1 _19219_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12963_ _19432_/Q vssd1 vssd1 vccd1 vccd1 _16351_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09172__C _09172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09876__C1 _09754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13690__S _13690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14702_ _14702_/A vssd1 vssd1 vccd1 vccd1 _18809_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18470_ _19491_/CLK _18470_/D vssd1 vssd1 vccd1 vccd1 _18470_/Q sky130_fd_sc_hd__dfxtp_1
X_11914_ _16967_/A _11939_/C _11913_/Y vssd1 vssd1 vccd1 vccd1 _11914_/X sky130_fd_sc_hd__o21a_1
X_15682_ _14582_/X _19189_/Q _15682_/S vssd1 vssd1 vccd1 vccd1 _15683_/A sky130_fd_sc_hd__mux2_1
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ _19429_/Q vssd1 vssd1 vccd1 vccd1 _16340_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16286__B _16286_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17421_ _17541_/A vssd1 vssd1 vccd1 vccd1 _17422_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14633_ _14633_/A vssd1 vssd1 vccd1 vccd1 _18781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _19779_/Q _11291_/A _11925_/S vssd1 vssd1 vccd1 vccd1 _17198_/A sky130_fd_sc_hd__mux2_2
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output104_A _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17352_ _17199_/X _17246_/X _17367_/S vssd1 vssd1 vccd1 vccd1 _17498_/B sky130_fd_sc_hd__mux2_1
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14564_ _14563_/X _18760_/Q _14567_/S vssd1 vssd1 vccd1 vccd1 _14565_/A sky130_fd_sc_hd__mux2_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11776_ _19636_/Q vssd1 vssd1 vccd1 vccd1 _16953_/A sky130_fd_sc_hd__inv_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16303_/A vssd1 vssd1 vccd1 vccd1 _19419_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ _13596_/A vssd1 vssd1 vccd1 vccd1 _13615_/S sky130_fd_sc_hd__buf_6
XFILLER_159_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17283_ _12289_/A _17605_/B _17283_/S vssd1 vssd1 vccd1 vccd1 _17283_/X sky130_fd_sc_hd__mux2_1
X_10727_ _18922_/Q _18688_/Q _19370_/Q _19018_/Q _11299_/S _09590_/A vssd1 vssd1 vccd1
+ vccd1 _10728_/B sky130_fd_sc_hd__mux4_1
X_14495_ _14495_/A vssd1 vssd1 vccd1 vccd1 _18731_/D sky130_fd_sc_hd__clkbuf_1
X_19022_ _19086_/CLK _19022_/D vssd1 vssd1 vccd1 vccd1 _19022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16234_ _16234_/A vssd1 vssd1 vccd1 vccd1 _19388_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09909__A _09909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13446_ _12865_/X _18324_/Q _13448_/S vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10658_ _19277_/Q _19115_/Q _18524_/Q _18294_/Q _10650_/X _11298_/A vssd1 vssd1 vccd1
+ vccd1 _10659_/B sky130_fd_sc_hd__mux4_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16165_ _19770_/Q _16165_/B vssd1 vssd1 vccd1 vccd1 _16165_/Y sky130_fd_sc_hd__xnor2_1
X_13377_ _19583_/Q _13055_/X _13376_/X _13265_/X vssd1 vssd1 vccd1 vccd1 _13377_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10636__S1 _10567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10589_ _18463_/Q _19054_/Q _19216_/Q _18431_/Q _10017_/S _10577_/X vssd1 vssd1 vccd1
+ vccd1 _10590_/B sky130_fd_sc_hd__mux4_2
XFILLER_6_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15116_ _15116_/A vssd1 vssd1 vccd1 vccd1 _18981_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12328_ _12321_/A _12319_/X _12324_/X _12327_/Y vssd1 vssd1 vccd1 vccd1 _12328_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_115_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16096_ _16096_/A vssd1 vssd1 vccd1 vccd1 _19346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13865__S _13871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15047_ _15047_/A vssd1 vssd1 vccd1 vccd1 _15047_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12259_ _19415_/Q _12093_/X _12255_/X _12258_/Y vssd1 vssd1 vccd1 vccd1 _16295_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__16429__B1 _16402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11893__B _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09644__A _09644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19855_ _19865_/CLK _19855_/D vssd1 vssd1 vccd1 vccd1 _19855_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11061__S1 _11012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18806_ _19471_/CLK _18806_/D vssd1 vssd1 vccd1 vccd1 _18806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13166__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19786_ _19786_/CLK _19786_/D vssd1 vssd1 vccd1 vccd1 _19786_/Q sky130_fd_sc_hd__dfxtp_1
X_16998_ _19652_/Q _16998_/B vssd1 vssd1 vccd1 vccd1 _16998_/X sky130_fd_sc_hd__or2_1
XFILLER_23_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18737_ _19387_/CLK _18737_/D vssd1 vssd1 vccd1 vccd1 _18737_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14696__S _14698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15949_ _15949_/A vssd1 vssd1 vccd1 vccd1 _19307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16477__A _16868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10302__B _12468_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__B1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09470_ _09470_/A vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18668_ _19088_/CLK _18668_/D vssd1 vssd1 vccd1 vccd1 _18668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17619_ _17571_/A _17618_/X _17477_/X vssd1 vssd1 vccd1 vccd1 _17619_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10492__A3 _10490_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10729__S _10729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18599_ _18902_/CLK _18599_/D vssd1 vssd1 vccd1 vccd1 _18599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_178_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11414__A _11416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10324__S0 _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15320__S _15328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12245__A _12245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09554__A _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10165__C1 _09831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15990__S _15992_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ _10209_/A vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__buf_2
XFILLER_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09737_ _09737_/A vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15291__A _15302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09668_ _10040_/A vssd1 vssd1 vccd1 vccd1 _09669_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_131_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _10654_/A vssd1 vssd1 vccd1 vccd1 _09599_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _11619_/A _18112_/A _12730_/C vssd1 vssd1 vccd1 vccd1 _11630_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11561_ _11566_/A _18102_/A _17122_/C _17175_/D vssd1 vssd1 vccd1 vccd1 _17169_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18107__A _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ _19691_/Q _13008_/X _13009_/X _19658_/Q vssd1 vssd1 vccd1 vccd1 _13300_/X
+ sky130_fd_sc_hd__a22o_1
X_10512_ _18464_/Q _19055_/Q _19217_/Q _18432_/Q _10496_/X _09710_/A vssd1 vssd1 vccd1
+ vccd1 _10512_/X sky130_fd_sc_hd__mux4_1
XFILLER_155_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09729__A _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14280_ _14290_/A _18216_/B vssd1 vssd1 vccd1 vccd1 _14281_/A sky130_fd_sc_hd__and2_2
XFILLER_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11492_ _17120_/D _11492_/B _11492_/C _11492_/D vssd1 vssd1 vccd1 vccd1 _11492_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_171_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _19762_/Q vssd1 vssd1 vccd1 vccd1 _16126_/A sky130_fd_sc_hd__clkbuf_2
X_10443_ _10439_/A _10440_/X _10442_/X vssd1 vssd1 vccd1 vccd1 _10443_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_137_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12393__B1 _11686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13162_ _16887_/A _12501_/X _12503_/X _16474_/A _13161_/X vssd1 vssd1 vccd1 vccd1
+ _15566_/B sky130_fd_sc_hd__a221o_2
XANTENNA_input65_A io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _10237_/X _10371_/X _10373_/X _10243_/X vssd1 vssd1 vccd1 vccd1 _10374_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_163_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12113_ _17779_/A _12113_/B vssd1 vssd1 vccd1 vccd1 _12117_/A sky130_fd_sc_hd__xor2_1
XFILLER_124_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13093_ input7/X _12974_/A _12977_/A vssd1 vssd1 vccd1 vccd1 _13105_/A sky130_fd_sc_hd__a21o_1
X_17970_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17979_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16921_ _19624_/Q _16920_/X _16921_/S vssd1 vssd1 vccd1 vccd1 _16922_/A sky130_fd_sc_hd__mux2_1
X_12044_ _19646_/Q _19645_/Q _12044_/C vssd1 vssd1 vccd1 vccd1 _12105_/C sky130_fd_sc_hd__and3_1
X_19640_ _19669_/CLK _19640_/D vssd1 vssd1 vccd1 vccd1 _19640_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_5_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16852_ _16854_/A _16854_/C _16812_/X vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__a21oi_1
X_15803_ _15803_/A vssd1 vssd1 vccd1 vccd1 _19242_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19571_ _19668_/CLK _19571_/D vssd1 vssd1 vccd1 vccd1 _19571_/Q sky130_fd_sc_hd__dfxtp_1
X_16783_ _16840_/A _16790_/C vssd1 vssd1 vccd1 vccd1 _16783_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13995_ _18527_/Q _13994_/X _13995_/S vssd1 vssd1 vccd1 vccd1 _13996_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09313__A1 _19708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15734_ _15780_/S vssd1 vssd1 vccd1 vccd1 _15743_/S sky130_fd_sc_hd__buf_2
X_18522_ _19081_/CLK _18522_/D vssd1 vssd1 vccd1 vccd1 _18522_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12946_ _12945_/X _18290_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12947_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15665_ _14557_/X _19181_/Q _15671_/S vssd1 vssd1 vccd1 vccd1 _15666_/A sky130_fd_sc_hd__mux2_1
X_18453_ _19302_/CLK _18453_/D vssd1 vssd1 vccd1 vccd1 _18453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12975__D input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ _16752_/D _12701_/X _12876_/X _12707_/X vssd1 vssd1 vccd1 vccd1 _12877_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17404_/A _17404_/B _17404_/C vssd1 vssd1 vccd1 vccd1 _17584_/A sky130_fd_sc_hd__nor3_2
XFILLER_60_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14616_ _14616_/A vssd1 vssd1 vccd1 vccd1 _18776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14070__A0 _13864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18384_ _19071_/CLK _18384_/D vssd1 vssd1 vccd1 vccd1 _18384_/Q sky130_fd_sc_hd__dfxtp_1
X_11828_ _11827_/Y _11824_/Y _14275_/B vssd1 vssd1 vccd1 vccd1 _11828_/X sky130_fd_sc_hd__mux2_1
X_15596_ _15595_/X _19162_/Q _15596_/S vssd1 vssd1 vccd1 vccd1 _15597_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10306__S0 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09616__A2 _09604_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17524_/S vssd1 vssd1 vccd1 vccd1 _17461_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14547_ _14547_/A vssd1 vssd1 vccd1 vccd1 _14547_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10226__A3 _10224_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11759_ _19776_/Q _11016_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _17250_/A sky130_fd_sc_hd__mux2_4
XFILLER_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17266_ _17266_/A vssd1 vssd1 vccd1 vccd1 _17375_/S sky130_fd_sc_hd__clkbuf_2
X_14478_ _13886_/X _18724_/Q _14478_/S vssd1 vssd1 vccd1 vccd1 _14479_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16217_ _16217_/A vssd1 vssd1 vccd1 vccd1 _19380_/D sky130_fd_sc_hd__clkbuf_1
X_19005_ _19292_/CLK _19005_/D vssd1 vssd1 vccd1 vccd1 _19005_/Q sky130_fd_sc_hd__dfxtp_1
X_13429_ _16162_/S _17023_/A vssd1 vssd1 vccd1 vccd1 _13430_/B sky130_fd_sc_hd__nor2_2
XANTENNA__17856__A _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12065__A _12066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17197_ _17642_/B _12219_/A _17251_/S vssd1 vssd1 vccd1 vccd1 _17197_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16760__A _19561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16148_ _16148_/A vssd1 vssd1 vccd1 vccd1 _19355_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16079_ _19755_/Q _16080_/B vssd1 vssd1 vccd1 vccd1 _16091_/C sky130_fd_sc_hd__or2_1
XANTENNA__14280__A _14290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09374__A _09374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19838_ _19838_/CLK _19838_/D vssd1 vssd1 vccd1 vccd1 _19838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15625__A1 _15612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput1 io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_2
X_19769_ _19799_/CLK _19769_/D vssd1 vssd1 vccd1 vccd1 _19769_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09522_ _10854_/S vssd1 vssd1 vccd1 vccd1 _10579_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15315__S _15315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ _19199_/Q _18813_/Q _19263_/Q _18382_/Q _10496_/A _09390_/A vssd1 vssd1 vccd1
+ vccd1 _09454_/B sky130_fd_sc_hd__mux4_1
XFILLER_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16935__A _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14061__A0 _13851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09384_ _11050_/S vssd1 vssd1 vccd1 vccd1 _09396_/A sky130_fd_sc_hd__buf_2
XFILLER_33_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12914__A2 _12817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11273__S1 _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12703__A _13008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09131__B1_N input33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10090_ _10090_/A vssd1 vssd1 vccd1 vccd1 _10090_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12678__A1 _19161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11025__S1 _11266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12678__B2 _19351_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15616__A1 _15615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16813__B1 _16812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12800_ _14996_/A vssd1 vssd1 vccd1 vccd1 _14519_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_56_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13780_ _13780_/A vssd1 vssd1 vccd1 vccd1 _18454_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10992_ _18486_/Q _18981_/Q _11243_/S vssd1 vssd1 vccd1 vccd1 _10992_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12731_ _18253_/Q _12727_/X _11284_/A _12747_/A _12730_/X vssd1 vssd1 vccd1 vccd1
+ _18253_/D sky130_fd_sc_hd__a221o_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15450_ _15450_/A vssd1 vssd1 vccd1 vccd1 _19130_/D sky130_fd_sc_hd__clkbuf_1
X_12662_ _19676_/Q _12659_/X _12565_/A _16974_/A _12661_/X vssd1 vssd1 vccd1 vccd1
+ _12662_/X sky130_fd_sc_hd__a221o_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14401_ _14401_/A vssd1 vssd1 vccd1 vccd1 _18689_/D sky130_fd_sc_hd__clkbuf_1
X_11613_ _14272_/A _14275_/A vssd1 vssd1 vccd1 vccd1 _11887_/A sky130_fd_sc_hd__nor2_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15381_ _19100_/Q _15089_/X _15383_/S vssd1 vssd1 vccd1 vccd1 _15382_/A sky130_fd_sc_hd__mux2_1
X_12593_ _17026_/S _12593_/B vssd1 vssd1 vccd1 vccd1 _12593_/X sky130_fd_sc_hd__and2_1
XFILLER_129_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17120_ _17120_/A _17120_/B _17120_/C _17120_/D vssd1 vssd1 vccd1 vccd1 _17122_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_156_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14332_ _13886_/X _18660_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14333_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11544_ _12447_/A _17133_/A vssd1 vssd1 vccd1 vccd1 _11544_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17051_ _17051_/A vssd1 vssd1 vccd1 vccd1 _19673_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15552__A0 _19722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ _14263_/A vssd1 vssd1 vccd1 vccd1 _18637_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11475_ _11440_/X _11441_/Y _11442_/X _11443_/Y _11474_/X vssd1 vssd1 vccd1 vccd1
+ _11475_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11169__A1 _09477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16002_ _16146_/A vssd1 vssd1 vccd1 vccd1 _16119_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11169__B2 _11168_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ _13234_/A _13214_/B _13233_/B vssd1 vssd1 vccd1 vccd1 _13214_/X sky130_fd_sc_hd__or3_1
X_10426_ _19315_/Q _18727_/Q _18764_/Q _18338_/Q _10339_/S _10270_/A vssd1 vssd1 vccd1
+ vccd1 _10426_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12905__A2 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14194_ _14194_/A vssd1 vssd1 vccd1 vccd1 _18607_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_100_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10916__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_126_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13145_ input10/X _13117_/X _13120_/X vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__a21o_1
X_10357_ _10419_/A _10357_/B vssd1 vssd1 vccd1 vccd1 _10357_/X sky130_fd_sc_hd__or2_1
XANTENNA__14304__S _14310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _19678_/Q _12703_/X _12704_/X _16978_/A vssd1 vssd1 vccd1 vccd1 _13076_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17953_ _16055_/B _19783_/Q _17957_/S vssd1 vssd1 vccd1 vccd1 _17954_/A sky130_fd_sc_hd__mux2_1
X_10288_ _10390_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10288_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12669__B2 _18263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16904_ _16904_/A _19614_/Q _16904_/C vssd1 vssd1 vccd1 vccd1 _16906_/B sky130_fd_sc_hd__and3_1
X_12027_ _12140_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12031_/A sky130_fd_sc_hd__xnor2_1
XFILLER_78_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10133__A _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17884_ _19734_/Q _17831_/X _17883_/X vssd1 vssd1 vccd1 vccd1 _19734_/D sky130_fd_sc_hd__o21a_1
X_19623_ _19669_/CLK _19623_/D vssd1 vssd1 vccd1 vccd1 _19623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16835_ _16836_/A _16836_/B _16834_/Y vssd1 vssd1 vccd1 vccd1 _19589_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19554_ _19828_/CLK _19554_/D vssd1 vssd1 vccd1 vccd1 _19554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16766_ _16772_/C _16772_/D _16765_/Y vssd1 vssd1 vccd1 vccd1 _19563_/D sky130_fd_sc_hd__o21a_1
X_13978_ _14550_/A vssd1 vssd1 vccd1 vccd1 _13978_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18505_ _18902_/CLK _18505_/D vssd1 vssd1 vccd1 vccd1 _18505_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15717_ _13522_/X _19204_/Q _15721_/S vssd1 vssd1 vccd1 vccd1 _15718_/A sky130_fd_sc_hd__mux2_1
X_12929_ _12929_/A _12971_/B vssd1 vssd1 vccd1 vccd1 _12929_/Y sky130_fd_sc_hd__nor2_1
X_16697_ _19542_/Q _19541_/Q _16697_/C _16697_/D vssd1 vssd1 vccd1 vccd1 _16706_/D
+ sky130_fd_sc_hd__and4_1
X_19485_ _19491_/CLK _19485_/D vssd1 vssd1 vccd1 vccd1 _19485_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18436_ _19124_/CLK _18436_/D vssd1 vssd1 vccd1 vccd1 _18436_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15648_ _15648_/A vssd1 vssd1 vccd1 vccd1 _19173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15791__A0 _13525_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15579_ _15579_/A vssd1 vssd1 vccd1 vccd1 _19158_/D sky130_fd_sc_hd__clkbuf_1
X_18367_ _19184_/CLK _18367_/D vssd1 vssd1 vccd1 vccd1 _18367_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10604__B1 _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17318_ _17415_/A vssd1 vssd1 vccd1 vccd1 _17319_/C sky130_fd_sc_hd__clkinv_2
XFILLER_159_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18298_ _19282_/CLK _18298_/D vssd1 vssd1 vccd1 vccd1 _18298_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15543__A0 _19721_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11411__B _12482_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17249_ _17246_/X _17346_/B _17266_/A vssd1 vssd1 vccd1 vccd1 _17249_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18088__A2 _18086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11255__S1 _11124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13619__A _13619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12523__A _13391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15045__S _15045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09505_ _10640_/A vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_53_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17220__A0 _17709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09436_ _09596_/A vssd1 vssd1 vccd1 vccd1 _10743_/A sky130_fd_sc_hd__clkbuf_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ _09367_/A vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_166_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09298_ _09295_/X _09296_/X _09297_/X _19620_/Q vssd1 vssd1 vccd1 vccd1 _11698_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_21_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09439__S1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11260_ _09366_/A _11250_/X _11259_/X _09469_/A _19707_/Q vssd1 vssd1 vccd1 vccd1
+ _11260_/X sky130_fd_sc_hd__a32o_2
XFILLER_137_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11246__S1 _11124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14632__B _18209_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _10214_/A _10210_/X _09909_/A vssd1 vssd1 vccd1 vccd1 _10211_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17826__A2 _17648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11191_ _11184_/X _11186_/X _11188_/X _11190_/X _09465_/A vssd1 vssd1 vccd1 vccd1
+ _11191_/X sky130_fd_sc_hd__a221o_2
XFILLER_122_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10142_ _18407_/Q _18668_/Q _18567_/Q _18902_/Q _09930_/S _09871_/X vssd1 vssd1 vccd1
+ vccd1 _10143_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13963__S _13963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ _10073_/A vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__buf_2
X_14950_ _18921_/Q vssd1 vssd1 vccd1 vccd1 _14951_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10757__S0 _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13901_ _13901_/A vssd1 vssd1 vccd1 vccd1 _18499_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09742__A _09859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input28_A io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14881_ _14881_/A vssd1 vssd1 vccd1 vccd1 _18888_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16620_ _19808_/Q _19806_/Q _19805_/Q vssd1 vssd1 vccd1 vccd1 _16622_/C sky130_fd_sc_hd__or3_1
X_13832_ _13832_/A vssd1 vssd1 vccd1 vccd1 _18478_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16551_ _19497_/Q _16551_/B _16551_/C vssd1 vssd1 vccd1 vccd1 _16552_/C sky130_fd_sc_hd__and3_1
XANTENNA__11087__B1 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13763_ _13763_/A vssd1 vssd1 vccd1 vccd1 _18448_/D sky130_fd_sc_hd__clkbuf_1
X_10975_ _09482_/A _10961_/Y _10966_/X _10974_/Y _09658_/A vssd1 vssd1 vccd1 vccd1
+ _10975_/X sky130_fd_sc_hd__o311a_1
XFILLER_44_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16575__A _19506_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10400__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A vssd1 vssd1 vccd1 vccd1 _15549_/A sky130_fd_sc_hd__buf_2
X_15502_ _19714_/Q _16919_/A _15516_/S vssd1 vssd1 vccd1 vccd1 _15502_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16482_ _16483_/B _16483_/C _16481_/Y vssd1 vssd1 vccd1 vccd1 _19478_/D sky130_fd_sc_hd__o21a_1
X_19270_ _19301_/CLK _19270_/D vssd1 vssd1 vccd1 vccd1 _19270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_71_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13694_ _13762_/S vssd1 vssd1 vccd1 vccd1 _13703_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15433_ _19123_/Q _15060_/X _15433_/S vssd1 vssd1 vccd1 vccd1 _15434_/A sky130_fd_sc_hd__mux2_1
X_18221_ _18221_/A vssd1 vssd1 vccd1 vccd1 _19857_/D sky130_fd_sc_hd__clkbuf_1
X_12645_ _16772_/C _12638_/X _12643_/X _12644_/X vssd1 vssd1 vccd1 vccd1 _12645_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12587__B1 _13356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15364_ _19092_/Q _15063_/X _15372_/S vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__mux2_1
X_18152_ _09236_/C _12674_/A _18148_/Y input45/X vssd1 vssd1 vccd1 vccd1 _18153_/B
+ sky130_fd_sc_hd__o22a_1
X_12576_ _12557_/X _12572_/X _12574_/Y _12575_/X _18268_/Q vssd1 vssd1 vccd1 vccd1
+ _12577_/B sky130_fd_sc_hd__a32o_4
XFILLER_129_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17103_ _17163_/A vssd1 vssd1 vccd1 vccd1 _17142_/A sky130_fd_sc_hd__clkbuf_2
X_14315_ _13861_/X _18652_/Q _14321_/S vssd1 vssd1 vccd1 vccd1 _14316_/A sky130_fd_sc_hd__mux2_1
X_18083_ _18083_/A _18087_/B vssd1 vssd1 vccd1 vccd1 _18083_/X sky130_fd_sc_hd__or2_1
X_11527_ _17121_/B _11574_/B _12475_/A vssd1 vssd1 vccd1 vccd1 _11564_/C sky130_fd_sc_hd__o21ai_1
X_15295_ _15295_/A vssd1 vssd1 vccd1 vccd1 _19061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17034_ _17034_/A vssd1 vssd1 vccd1 vccd1 _19665_/D sky130_fd_sc_hd__clkbuf_1
X_14246_ _14246_/A vssd1 vssd1 vccd1 vccd1 _18629_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output96_A _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ _11456_/X _11295_/Y _11457_/X vssd1 vssd1 vccd1 vccd1 _11458_/X sky130_fd_sc_hd__o21a_1
X_10409_ _10461_/A _10409_/B vssd1 vssd1 vccd1 vccd1 _10409_/X sky130_fd_sc_hd__or2_1
XANTENNA__13439__A _13507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14177_ _14177_/A vssd1 vssd1 vccd1 vccd1 _18599_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14034__S _14043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11389_ _11389_/A _11389_/B vssd1 vssd1 vccd1 vccd1 _11389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_140_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10996__S0 _11196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ _19756_/Q vssd1 vssd1 vccd1 vccd1 _16091_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _19367_/CLK _18985_/D vssd1 vssd1 vccd1 vccd1 _18985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10770__C1 _09602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _19437_/Q _13005_/X _13058_/X vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__o21a_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _17936_/A vssd1 vssd1 vccd1 vccd1 _19743_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17867_ _17867_/A _17867_/B vssd1 vssd1 vccd1 vccd1 _17867_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_2_2_0_clock clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_5_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19606_ _19607_/CLK _19606_/D vssd1 vssd1 vccd1 vccd1 _19606_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16818_ hold22/A _19578_/Q _16816_/B _16810_/C _18163_/A vssd1 vssd1 vccd1 vccd1
+ _16818_/X sky130_fd_sc_hd__a41o_1
XANTENNA__13067__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17798_ _17802_/A _17802_/B _17842_/S vssd1 vssd1 vccd1 vccd1 _17798_/X sky130_fd_sc_hd__mux2_1
XFILLER_54_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19537_ _19540_/CLK _19537_/D vssd1 vssd1 vccd1 vccd1 _19537_/Q sky130_fd_sc_hd__dfxtp_1
X_16749_ _19557_/Q _19556_/Q _19553_/Q _19552_/Q vssd1 vssd1 vccd1 vccd1 _16750_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19468_ _19603_/CLK _19468_/D vssd1 vssd1 vccd1 vccd1 _19468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ _11618_/A _19813_/Q vssd1 vssd1 vccd1 vccd1 _09221_/X sky130_fd_sc_hd__xor2_1
X_18419_ _19202_/CLK _18419_/D vssd1 vssd1 vccd1 vccd1 _18419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19399_ _19838_/CLK _19399_/D vssd1 vssd1 vccd1 vccd1 _19399_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__14209__S _14209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _19866_/Q _19841_/Q _19840_/Q _19839_/Q vssd1 vssd1 vccd1 vccd1 _09176_/B
+ sky130_fd_sc_hd__and4bb_2
XFILLER_148_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15516__A0 _19716_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09083_ _19849_/Q vssd1 vssd1 vccd1 vccd1 _09174_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10038__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput70 reset vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_6
XFILLER_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17808__A2 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12253__A _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12750__B1 _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ _18603_/Q _18874_/Q _19098_/Q _18842_/Q _10602_/S _09977_/X vssd1 vssd1 vccd1
+ vccd1 _09985_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13058__A1 _19565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17184__D_N _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10760_ _09434_/A _10753_/X _10755_/X _10759_/X _09614_/X vssd1 vssd1 vccd1 vccd1
+ _10760_/X sky130_fd_sc_hd__a311o_4
XFILLER_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12281__A2 _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10911__S0 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10292__A1 _10394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ _09419_/A vssd1 vssd1 vccd1 vccd1 _09671_/A sky130_fd_sc_hd__buf_4
XFILLER_160_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_clock clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
X_10691_ _10691_/A vssd1 vssd1 vccd1 vccd1 _10691_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16952__C1 _16933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _12430_/A _12430_/B _12430_/C vssd1 vssd1 vccd1 vccd1 _12432_/A sky130_fd_sc_hd__nand3_4
XFILLER_166_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10044__A1 _10046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12361_ _12388_/A _12361_/B vssd1 vssd1 vccd1 vccd1 _12363_/C sky130_fd_sc_hd__nand2_1
XFILLER_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14100_ _14100_/A vssd1 vssd1 vccd1 vccd1 _18565_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10595__A2 _10583_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ _18462_/Q _19053_/Q _19215_/Q _18430_/Q _10660_/X _10655_/X vssd1 vssd1 vccd1
+ vccd1 _11313_/B sky130_fd_sc_hd__mux4_1
XFILLER_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_6_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19373_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_153_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09737__A _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16180__A0 _13528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15080_ _15080_/A vssd1 vssd1 vccd1 vccd1 _15093_/S sky130_fd_sc_hd__buf_4
XFILLER_4_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _19417_/Q _12293_/B vssd1 vssd1 vccd1 vccd1 _12294_/A sky130_fd_sc_hd__nor2_1
XFILLER_154_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14031_ _18538_/Q _14029_/X _14043_/S vssd1 vssd1 vccd1 vccd1 _14032_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09198__C1 _19701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11243_ _18609_/Q _18944_/Q _11243_/S vssd1 vssd1 vccd1 vccd1 _11243_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11174_ _11174_/A _11174_/B vssd1 vssd1 vccd1 vccd1 _11174_/X sky130_fd_sc_hd__and2_1
XFILLER_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10125_ _11390_/A _10125_/B vssd1 vssd1 vccd1 vccd1 _10125_/Y sky130_fd_sc_hd__nor2_1
X_18770_ _19256_/CLK _18770_/D vssd1 vssd1 vccd1 vccd1 _18770_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14494__A0 _13909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15982_ _15982_/A vssd1 vssd1 vccd1 vccd1 _19322_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_122_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13297__A1 input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17721_ _17648_/S _17360_/X _17402_/A vssd1 vssd1 vccd1 vccd1 _17721_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14933_ _14933_/A vssd1 vssd1 vccd1 vccd1 _18912_/D sky130_fd_sc_hd__clkbuf_1
X_10056_ _10056_/A _10056_/B vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_94_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17652_ _17795_/A vssd1 vssd1 vccd1 vccd1 _17652_/X sky130_fd_sc_hd__clkbuf_4
X_14864_ _14864_/A vssd1 vssd1 vccd1 vccd1 _18880_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16603_ _19514_/Q _16604_/C _19515_/Q vssd1 vssd1 vccd1 vccd1 _16605_/B sky130_fd_sc_hd__a21oi_1
X_13815_ _13815_/A vssd1 vssd1 vccd1 vccd1 _18470_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17583_ _17587_/A _17587_/B vssd1 vssd1 vccd1 vccd1 _17583_/Y sky130_fd_sc_hd__nand2_1
X_14795_ _18850_/Q _13956_/X _14799_/S vssd1 vssd1 vccd1 vccd1 _14796_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19322_ _19610_/CLK _19322_/D vssd1 vssd1 vccd1 vccd1 _19322_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16534_ _16542_/D vssd1 vssd1 vccd1 vccd1 _16540_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13746_ _13746_/A vssd1 vssd1 vccd1 vccd1 _18440_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ _09432_/A _10951_/X _10953_/X _10957_/X _09614_/A vssd1 vssd1 vccd1 vccd1
+ _10958_/X sky130_fd_sc_hd__a311o_2
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17735__A1 _17734_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10283__A1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19253_ _19379_/CLK _19253_/D vssd1 vssd1 vccd1 vccd1 _19253_/Q sky130_fd_sc_hd__dfxtp_1
X_16465_ _16466_/B _16466_/C _16464_/Y vssd1 vssd1 vccd1 vccd1 _19472_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13677_ _13677_/A vssd1 vssd1 vccd1 vccd1 _13686_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_32_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _10889_/A _10889_/B vssd1 vssd1 vccd1 vccd1 _10889_/X sky130_fd_sc_hd__or2_1
XFILLER_148_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18204_ _18233_/A vssd1 vssd1 vccd1 vccd1 _18213_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_12628_ _16929_/B _12598_/X _12623_/X _12627_/X vssd1 vssd1 vccd1 vccd1 _19620_/D
+ sky130_fd_sc_hd__a22o_1
X_15416_ _19115_/Q _15035_/X _15422_/S vssd1 vssd1 vccd1 vccd1 _15417_/A sky130_fd_sc_hd__mux2_1
X_16396_ _19448_/Q _19447_/Q _16396_/C vssd1 vssd1 vccd1 vccd1 _16399_/B sky130_fd_sc_hd__and3_1
X_19184_ _19184_/CLK _19184_/D vssd1 vssd1 vccd1 vccd1 _19184_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12024__A2 _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16752__B _16752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13868__S _13871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18135_ _18135_/A _18135_/B vssd1 vssd1 vccd1 vccd1 _18135_/X sky130_fd_sc_hd__or2_1
X_15347_ _15347_/A vssd1 vssd1 vccd1 vccd1 _19084_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10035__B2 _10042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12559_ _16689_/C _12507_/X _12511_/X _19505_/Q vssd1 vssd1 vccd1 vccd1 _13132_/B
+ sky130_fd_sc_hd__a22o_2
XFILLER_145_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18066_ _19802_/Q _19423_/Q _18066_/S vssd1 vssd1 vccd1 vccd1 _18067_/A sky130_fd_sc_hd__mux2_1
X_15278_ _14566_/X _19054_/Q _15278_/S vssd1 vssd1 vccd1 vccd1 _15279_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17017_ _15620_/X _17010_/X _17016_/X _17008_/X vssd1 vssd1 vccd1 vccd1 _19659_/D
+ sky130_fd_sc_hd__o211a_1
X_14229_ _18622_/Q _13991_/X _14231_/S vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__mux2_1
XFILLER_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12732__A0 _18114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _10270_/A vssd1 vssd1 vccd1 vccd1 _10382_/A sky130_fd_sc_hd__buf_2
XFILLER_101_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17671__B1 _17670_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18968_ _19290_/CLK _18968_/D vssd1 vssd1 vccd1 vccd1 _18968_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09382__A _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17919_ _17920_/A _17744_/S _17626_/A _17918_/X vssd1 vssd1 vccd1 vccd1 _17919_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11814__A2_N _12450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18899_ _19285_/CLK _18899_/D vssd1 vssd1 vccd1 vccd1 _18899_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17423__B1 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16927__B _16929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14728__A _14785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12799__B1 _12795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16934__C1 _16933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16943__A _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ _18109_/A _19811_/Q _09200_/X _09201_/Y _09203_/Y vssd1 vssd1 vccd1 vccd1
+ _09204_/X sky130_fd_sc_hd__o2111a_1
XFILLER_33_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10026__A1 _09485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09135_ _11575_/A vssd1 vssd1 vccd1 vccd1 _11567_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_147_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16162__A0 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09557__A _09557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09276__B _13356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10329__A2 _10319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_144_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17331__C_N _17190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ _09968_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _09968_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14402__S _14406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09292__A _12621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09899_ _18634_/Q _18969_/Q _10168_/S vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11930_ _11903_/A _11903_/B _11900_/A vssd1 vssd1 vccd1 vccd1 _11931_/B sky130_fd_sc_hd__a21boi_1
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _11794_/A _11858_/X _11860_/Y vssd1 vssd1 vccd1 vccd1 _11861_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11137__S0 _11173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15233__S _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13600_ _18379_/Q _13599_/X _13609_/S vssd1 vssd1 vccd1 vccd1 _13601_/A sky130_fd_sc_hd__mux2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ _11252_/A vssd1 vssd1 vccd1 vccd1 _11184_/A sky130_fd_sc_hd__clkbuf_8
X_14580_ _14579_/X _18765_/Q _14583_/S vssd1 vssd1 vccd1 vccd1 _14581_/A sky130_fd_sc_hd__mux2_1
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11792_ _19398_/Q vssd1 vssd1 vccd1 vccd1 _11826_/A sky130_fd_sc_hd__buf_4
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15728__A0 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ _15015_/A vssd1 vssd1 vccd1 vccd1 _13531_/X sky130_fd_sc_hd__buf_2
X_10743_ _10743_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10360__S1 _10229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16250_ _16250_/A vssd1 vssd1 vccd1 vccd1 _19395_/D sky130_fd_sc_hd__clkbuf_1
X_13462_ _13025_/X _18331_/Q _13470_/S vssd1 vssd1 vccd1 vccd1 _13463_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10674_ _10669_/X _10671_/X _10672_/X _11309_/A _09995_/A vssd1 vssd1 vccd1 vccd1
+ _10674_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09407__B1 _10046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _15201_/A vssd1 vssd1 vccd1 vccd1 _19019_/D sky130_fd_sc_hd__clkbuf_1
X_12413_ _19358_/Q _12069_/X _12412_/X _12075_/X vssd1 vssd1 vccd1 vccd1 _12413_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11214__B1 _09469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13688__S _13690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16181_ _16181_/A vssd1 vssd1 vccd1 vccd1 _19364_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13393_ _12230_/A _13390_/X _15463_/A vssd1 vssd1 vccd1 vccd1 _13431_/S sky130_fd_sc_hd__a21o_1
XFILLER_138_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_154_clock clkbuf_opt_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19237_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_15132_ _18989_/Q _15041_/X _15134_/S vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__mux2_1
X_12344_ _19658_/Q _12326_/X _16086_/A vssd1 vssd1 vccd1 vccd1 _12344_/Y sky130_fd_sc_hd__o21ai_1
X_15063_ _15063_/A vssd1 vssd1 vccd1 vccd1 _15063_/X sky130_fd_sc_hd__clkbuf_2
X_12275_ _19655_/Q vssd1 vssd1 vccd1 vccd1 _17005_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14014_ _14030_/A vssd1 vssd1 vccd1 vccd1 _14027_/S sky130_fd_sc_hd__clkbuf_4
X_11226_ _11042_/A _11216_/Y _11221_/X _11225_/Y _09552_/A vssd1 vssd1 vccd1 vccd1
+ _11226_/X sky130_fd_sc_hd__o311a_1
XFILLER_141_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_169_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19071_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18822_ _19272_/CLK _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11157_ _11164_/A _11156_/X _11042_/X vssd1 vssd1 vccd1 vccd1 _11157_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10108_ _10108_/A _10108_/B vssd1 vssd1 vccd1 vccd1 _10108_/X sky130_fd_sc_hd__or2_1
X_18753_ _19306_/CLK _18753_/D vssd1 vssd1 vccd1 vccd1 _18753_/Q sky130_fd_sc_hd__dfxtp_1
X_15965_ _15965_/A vssd1 vssd1 vccd1 vccd1 _19314_/D sky130_fd_sc_hd__clkbuf_1
X_11088_ _19270_/Q _19108_/Q _18517_/Q _18287_/Q _10964_/S _11033_/X vssd1 vssd1 vccd1
+ vccd1 _11089_/B sky130_fd_sc_hd__mux4_1
X_17704_ _17477_/X _17699_/X _17703_/X _17518_/X _11968_/B vssd1 vssd1 vccd1 vccd1
+ _17704_/X sky130_fd_sc_hd__a32o_1
X_14916_ _14916_/A vssd1 vssd1 vccd1 vccd1 _18904_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10039_ _10046_/A _10036_/X _10038_/X _09989_/X vssd1 vssd1 vccd1 vccd1 _10040_/C
+ sky130_fd_sc_hd__o211a_1
X_18684_ _19367_/CLK _18684_/D vssd1 vssd1 vccd1 vccd1 _18684_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15896_ _19284_/Q _14579_/A _15898_/S vssd1 vssd1 vccd1 vccd1 _15897_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11150__C1 _11020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17635_ _17571_/X _17624_/X _17634_/X _17592_/X vssd1 vssd1 vccd1 vccd1 _17635_/X
+ sky130_fd_sc_hd__o211a_1
X_14847_ _14847_/A vssd1 vssd1 vccd1 vccd1 _18873_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16239__S _16239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15143__S _15145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17566_ _17390_/X _17871_/B _17565_/X _17333_/X vssd1 vssd1 vccd1 vccd1 _17566_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_107_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19828_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17708__A1 _17709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14778_ _14778_/A vssd1 vssd1 vccd1 vccd1 _18843_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10256__A1 _10323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19305_ _19305_/CLK _19305_/D vssd1 vssd1 vccd1 vccd1 _19305_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15719__A0 _13525_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16517_ _19617_/Q _19616_/Q _19618_/Q _16907_/A vssd1 vssd1 vccd1 vccd1 _16522_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_143_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13729_ _13729_/A vssd1 vssd1 vccd1 vccd1 _18432_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17497_ _17353_/X _17356_/X _17497_/S vssd1 vssd1 vccd1 vccd1 _17613_/B sky130_fd_sc_hd__mux2_1
XFILLER_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09661__A3 _09659_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19236_ _19300_/CLK _19236_/D vssd1 vssd1 vccd1 vccd1 _19236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16448_ _16450_/B _16450_/C _16447_/Y vssd1 vssd1 vccd1 vccd1 _19466_/D sky130_fd_sc_hd__o21a_1
XFILLER_104_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19167_ _19598_/CLK _19167_/D vssd1 vssd1 vccd1 vccd1 _19167_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09949__B2 _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16379_ _19442_/Q _19441_/Q _16379_/C vssd1 vssd1 vccd1 vccd1 _16381_/B sky130_fd_sc_hd__and3_1
XFILLER_158_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__B2 _18132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11700__A _12974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18118_ _18118_/A _18142_/B vssd1 vssd1 vccd1 vccd1 _18118_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09377__A _10990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19098_ _19098_/CLK _19098_/D vssd1 vssd1 vccd1 vccd1 _19098_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18049_ _18049_/A vssd1 vssd1 vccd1 vccd1 _19794_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12705__B1 _12704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_174_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09822_/A vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__buf_2
XFILLER_101_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _09753_/A vssd1 vssd1 vccd1 vccd1 _09754_/A sky130_fd_sc_hd__buf_4
XFILLER_39_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09684_ _10185_/S vssd1 vssd1 vccd1 vccd1 _10093_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14458__A _14515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15988__S _15992_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_99_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11995__A1 _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_71_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19290_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_149_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18124__A1 _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _18104_/A _09325_/A vssd1 vssd1 vccd1 vccd1 _17120_/D sky130_fd_sc_hd__nor2_1
XFILLER_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10390_ _10390_/A _10390_/B vssd1 vssd1 vccd1 vccd1 _10390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12425__B _17232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_86_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19688_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_89_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12060_ _12060_/A vssd1 vssd1 vccd1 vccd1 _12063_/B sky130_fd_sc_hd__inv_2
XFILLER_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15228__S _15228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _11011_/A vssd1 vssd1 vccd1 vccd1 _11011_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_150_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09573__C1 _09829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14132__S _14136_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16848__A _16848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _12962_/A vssd1 vssd1 vccd1 vccd1 _12962_/X sky130_fd_sc_hd__clkbuf_2
X_15750_ _13570_/X _19219_/Q _15754_/S vssd1 vssd1 vccd1 vccd1 _15751_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input10_A io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ _16967_/A _11939_/C _13411_/A vssd1 vssd1 vccd1 vccd1 _11913_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14701_ _14601_/X _18809_/Q _14709_/S vssd1 vssd1 vccd1 vccd1 _14702_/A sky130_fd_sc_hd__mux2_1
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19264_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15681_ _15681_/A vssd1 vssd1 vccd1 vccd1 _19188_/D sky130_fd_sc_hd__clkbuf_1
X_12893_ _19493_/Q vssd1 vssd1 vccd1 vccd1 _16540_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17407_/A _17410_/B _17419_/X vssd1 vssd1 vccd1 vccd1 _17420_/X sky130_fd_sc_hd__o21a_1
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _17630_/A _11844_/B vssd1 vssd1 vccd1 vccd1 _11847_/A sky130_fd_sc_hd__xnor2_1
X_14632_ _14635_/A _18209_/B vssd1 vssd1 vccd1 vccd1 _14633_/A sky130_fd_sc_hd__and2_2
XFILLER_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15898__S _15898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14563_/A vssd1 vssd1 vccd1 vccd1 _14563_/X sky130_fd_sc_hd__clkbuf_1
X_17351_ _17461_/A _17341_/X _17350_/Y vssd1 vssd1 vccd1 vccd1 _17351_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _11750_/A _11749_/A _11774_/X vssd1 vssd1 vccd1 vccd1 _11778_/C sky130_fd_sc_hd__a21oi_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _18170_/A _16302_/B vssd1 vssd1 vccd1 vccd1 _16303_/A sky130_fd_sc_hd__and2_1
XFILLER_9_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13514_ _14860_/B _18091_/A _14860_/D _14642_/D vssd1 vssd1 vccd1 vccd1 _13596_/A
+ sky130_fd_sc_hd__and4b_4
X_10726_ _10703_/Y _09578_/A _09617_/X _10725_/X vssd1 vssd1 vccd1 vccd1 _12455_/B
+ sky130_fd_sc_hd__o22ai_4
Xclkbuf_leaf_39_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19389_/CLK sky130_fd_sc_hd__clkbuf_16
X_14494_ _13909_/X _18731_/Q _14500_/S vssd1 vssd1 vccd1 vccd1 _14495_/A sky130_fd_sc_hd__mux2_1
X_17282_ _17856_/B _17587_/B _17286_/S vssd1 vssd1 vccd1 vccd1 _17282_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_3_1_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_19021_ _19373_/CLK _19021_/D vssd1 vssd1 vccd1 vccd1 _19021_/Q sky130_fd_sc_hd__dfxtp_1
X_13445_ _13445_/A vssd1 vssd1 vccd1 vccd1 _18323_/D sky130_fd_sc_hd__clkbuf_1
X_16233_ _13605_/X _19388_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16234_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10657_ _11313_/A _10656_/X _09608_/A vssd1 vssd1 vccd1 vccd1 _10657_/X sky130_fd_sc_hd__o21a_1
XFILLER_139_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10097__S0 _10093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13376_ _19169_/Q _13179_/X _13374_/X _13375_/X vssd1 vssd1 vccd1 vccd1 _13376_/X
+ sky130_fd_sc_hd__a211o_1
X_16164_ _16164_/A vssd1 vssd1 vccd1 vccd1 _19358_/D sky130_fd_sc_hd__clkbuf_1
X_10588_ _10682_/A _10587_/X _09630_/X vssd1 vssd1 vccd1 vccd1 _10588_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12327_ _12075_/X _12325_/Y _12326_/X _16278_/A vssd1 vssd1 vccd1 vccd1 _12327_/Y
+ sky130_fd_sc_hd__o31ai_2
X_15115_ _18981_/Q _15015_/X _15123_/S vssd1 vssd1 vccd1 vccd1 _15116_/A sky130_fd_sc_hd__mux2_1
XFILLER_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16095_ _16094_/X _19346_/Q _16112_/S vssd1 vssd1 vccd1 vccd1 _16096_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15927__A _15983_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15046_ _15046_/A vssd1 vssd1 vccd1 vccd1 _18958_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ _12298_/C _12257_/Y _11665_/X vssd1 vssd1 vccd1 vccd1 _12258_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_123_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13360__A0 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11209_ _19267_/Q _19105_/Q _18514_/Q _18284_/Q _11128_/S _10801_/A vssd1 vssd1 vccd1
+ vccd1 _11209_/X sky130_fd_sc_hd__mux4_1
X_19854_ _19854_/CLK _19854_/D vssd1 vssd1 vccd1 vccd1 _19854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12189_ _12208_/A _12470_/B _12188_/Y vssd1 vssd1 vccd1 vccd1 _17810_/A sky130_fd_sc_hd__o21ai_4
XFILLER_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11371__C1 _09754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11910__A1 _19338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18805_ _19502_/CLK _18805_/D vssd1 vssd1 vccd1 vccd1 _18805_/Q sky130_fd_sc_hd__dfxtp_1
X_19785_ _19786_/CLK _19785_/D vssd1 vssd1 vccd1 vccd1 _19785_/Q sky130_fd_sc_hd__dfxtp_1
X_16997_ _17010_/A vssd1 vssd1 vccd1 vccd1 _16997_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__16758__A _19561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15662__A _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18736_ _19324_/CLK _18736_/D vssd1 vssd1 vccd1 vccd1 _18736_/Q sky130_fd_sc_hd__dfxtp_1
X_15948_ _13544_/X _19307_/Q _15948_/S vssd1 vssd1 vccd1 vccd1 _15949_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10477__A1 _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09660__A _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10021__S0 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18667_ _19286_/CLK _18667_/D vssd1 vssd1 vccd1 vccd1 _18667_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15879_ _19276_/Q _14553_/A _15887_/S vssd1 vssd1 vccd1 vccd1 _15880_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17618_ _17612_/Y _17617_/Y _17717_/S vssd1 vssd1 vccd1 vccd1 _17618_/X sky130_fd_sc_hd__mux2_2
X_18598_ _19223_/CLK _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11414__B _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17549_ _17613_/A _17350_/B _17548_/Y vssd1 vssd1 vccd1 vccd1 _17549_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19219_ _19315_/CLK _19219_/D vssd1 vssd1 vccd1 vccd1 _19219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17314__C1 _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10046__A _10046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12154__A1 _19347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__C1 _09811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09805_ _10335_/A vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input2_A io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14887__S _14893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13103__A0 _19722_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09736_ _11380_/A _09736_/B vssd1 vssd1 vccd1 vccd1 _09736_/X sky130_fd_sc_hd__or2_1
XFILLER_74_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09570__A _10929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18042__A0 _19791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A1 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ _09667_/A vssd1 vssd1 vccd1 vccd1 _09667_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09598_ _09598_/A vssd1 vssd1 vccd1 vccd1 _10654_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11560_ _11560_/A _11560_/B vssd1 vssd1 vccd1 vccd1 _17175_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14635__B _18211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ _10511_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10511_/X sky130_fd_sc_hd__or2_1
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11491_ _17120_/A _11491_/B vssd1 vssd1 vccd1 vccd1 _11492_/B sky130_fd_sc_hd__nor2_1
XFILLER_137_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13230_ _13230_/A vssd1 vssd1 vccd1 vccd1 _18305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ _10471_/A _10441_/X _10297_/A vssd1 vssd1 vccd1 vccd1 _10442_/X sky130_fd_sc_hd__o21a_1
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13161_ _19539_/Q _12507_/X _12511_/X _19507_/Q _13160_/X vssd1 vssd1 vccd1 vccd1
+ _13161_/X sky130_fd_sc_hd__a221o_2
XFILLER_137_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10373_ _10461_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10373_/X sky130_fd_sc_hd__or2_1
XFILLER_3_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18123__A _18136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12112_ _17743_/A _12140_/B _12140_/D _12305_/A vssd1 vssd1 vccd1 vccd1 _12113_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_163_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input58_A io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _13092_/A vssd1 vssd1 vccd1 vccd1 _18297_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16920_ _19620_/Q _12230_/X _12653_/B _16932_/A vssd1 vssd1 vccd1 vccd1 _16920_/X
+ sky130_fd_sc_hd__o22a_1
X_12043_ _16978_/A _12044_/C _19646_/Q vssd1 vssd1 vccd1 vccd1 _12043_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_123_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10251__S0 _10247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16851_ _19594_/Q _16847_/B _16850_/Y vssd1 vssd1 vccd1 vccd1 _19594_/D sky130_fd_sc_hd__o21a_1
XFILLER_78_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14797__S _14799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15802_ _13541_/X _19242_/Q _15804_/S vssd1 vssd1 vccd1 vccd1 _15803_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19570_ _19668_/CLK _19570_/D vssd1 vssd1 vccd1 vccd1 _19570_/Q sky130_fd_sc_hd__dfxtp_1
X_16782_ _19568_/Q _19567_/Q _16782_/C _16782_/D vssd1 vssd1 vccd1 vccd1 _16790_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_19_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13994_ _14566_/A vssd1 vssd1 vccd1 vccd1 _13994_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10459__A1 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18521_ _19081_/CLK _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10003__S0 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09313__A2 _09309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09944__S0 _10137_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15733_ _15733_/A vssd1 vssd1 vccd1 vccd1 _19211_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _14544_/A vssd1 vssd1 vccd1 vccd1 _12945_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _19205_/CLK _18452_/D vssd1 vssd1 vccd1 vccd1 _18452_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_122_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15664_ _15664_/A vssd1 vssd1 vccd1 vccd1 _19180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12876_ _19142_/Q _12784_/X _12874_/X _12875_/X vssd1 vssd1 vccd1 vccd1 _12876_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17403_ _17392_/X _17400_/X _17402_/X vssd1 vssd1 vccd1 vccd1 _17403_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14615_ _14614_/X _18776_/Q _14615_/S vssd1 vssd1 vccd1 vccd1 _14616_/A sky130_fd_sc_hd__mux2_1
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _19264_/CLK _18383_/D vssd1 vssd1 vccd1 vccd1 _18383_/Q sky130_fd_sc_hd__dfxtp_1
X_11827_ _11827_/A _11879_/C vssd1 vssd1 vccd1 vccd1 _11827_/Y sky130_fd_sc_hd__nor2_1
XFILLER_159_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15595_ _19731_/Q _12715_/X _15595_/S vssd1 vssd1 vccd1 vccd1 _15595_/X sky130_fd_sc_hd__mux2_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__S1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09616__A3 _09615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17334_ _17575_/S vssd1 vssd1 vccd1 vccd1 _17524_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__17202__A _17202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11758_ _17563_/A _11758_/B vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__xnor2_1
X_14546_ _14546_/A vssd1 vssd1 vccd1 vccd1 _18754_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10709_ _10721_/A _10709_/B vssd1 vssd1 vccd1 vccd1 _10709_/Y sky130_fd_sc_hd__nor2_1
X_17265_ _17779_/B _17709_/B _17283_/S vssd1 vssd1 vccd1 vccd1 _17265_/X sky130_fd_sc_hd__mux2_1
X_11689_ _19331_/Q _11859_/A vssd1 vssd1 vccd1 vccd1 _11689_/X sky130_fd_sc_hd__or2_1
X_14477_ _14477_/A vssd1 vssd1 vccd1 vccd1 _18723_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14037__S _14043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19004_ _19326_/CLK _19004_/D vssd1 vssd1 vccd1 vccd1 _19004_/Q sky130_fd_sc_hd__dfxtp_1
X_16216_ _13579_/X _19380_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16217_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13428_ hold4/X _12549_/X _13427_/X vssd1 vssd1 vccd1 vccd1 _17023_/A sky130_fd_sc_hd__a21oi_4
X_17196_ _17240_/S vssd1 vssd1 vccd1 vccd1 _17251_/S sky130_fd_sc_hd__buf_2
XANTENNA__17856__B _17856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16760__B _16760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13359_ _19661_/Q _12565_/X _13353_/X _13355_/X _13358_/X vssd1 vssd1 vccd1 vccd1
+ _13359_/X sky130_fd_sc_hd__a2111o_4
X_16147_ _16145_/X _19355_/Q _16167_/S vssd1 vssd1 vccd1 vccd1 _16148_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15322__A1 _15003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16078_ _16078_/A vssd1 vssd1 vccd1 vccd1 _19343_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12136__A1 _12126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14280__B _18216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_47_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13177__A _13234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15029_ _18953_/Q _15028_/X _15029_/S vssd1 vssd1 vccd1 vccd1 _15030_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17075__A1 _15574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19837_ _19838_/CLK _19837_/D vssd1 vssd1 vccd1 vccd1 _19837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14500__S _14500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 io_dbus_rdata[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_19768_ _19799_/CLK _19768_/D vssd1 vssd1 vccd1 vccd1 _19768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09521_ _09521_/A vssd1 vssd1 vccd1 vccd1 _09521_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09390__A _09390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18719_ _19307_/CLK _18719_/D vssd1 vssd1 vccd1 vccd1 _18719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09935__S0 _10137_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19699_ _19699_/CLK _19699_/D vssd1 vssd1 vccd1 vccd1 _19699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16000__B _16000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09452_ _10040_/A _09452_/B _09452_/C vssd1 vssd1 vccd1 vccd1 _09452_/X sky130_fd_sc_hd__or3_4
XFILLER_25_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09383_ _11011_/A vssd1 vssd1 vccd1 vccd1 _11050_/S sky130_fd_sc_hd__buf_4
XFILLER_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17112__A _17112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12611__A2 _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11160__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12375__A1 _12233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10386__B1 _09764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09528__C1 _09557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17066__A1 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16398__A _16868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09719_ _10509_/A vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10991_ _11065_/A vssd1 vssd1 vccd1 vccd1 _11243_/S sky130_fd_sc_hd__buf_4
XFILLER_28_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11335__A _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _18112_/A _17994_/S _12730_/C vssd1 vssd1 vccd1 vccd1 _12730_/X sky130_fd_sc_hd__and3_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _19150_/Q _12895_/A _12640_/X _19340_/Q _12660_/X vssd1 vssd1 vccd1 vccd1
+ _12661_/X sky130_fd_sc_hd__a221o_1
XFILLER_31_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15241__S _15243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ _11612_/A _17317_/A vssd1 vssd1 vccd1 vccd1 _11612_/X sky130_fd_sc_hd__xor2_4
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14400_ _13877_/X _18689_/Q _14406_/S vssd1 vssd1 vccd1 vccd1 _14401_/A sky130_fd_sc_hd__mux2_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ _12557_/X _12590_/X _12591_/Y _12575_/X _18269_/Q vssd1 vssd1 vccd1 vccd1
+ _12593_/B sky130_fd_sc_hd__a32o_4
X_15380_ _15380_/A vssd1 vssd1 vccd1 vccd1 _19099_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11543_ _12450_/A vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14331_ _14331_/A vssd1 vssd1 vccd1 vccd1 _18659_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17050_ _19673_/Q _15515_/X _17050_/S vssd1 vssd1 vccd1 vccd1 _17051_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14262_ _18637_/Q _14039_/X _14264_/S vssd1 vssd1 vccd1 vccd1 _14263_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15552__A1 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11474_ _11444_/X _11446_/Y _11447_/X _11448_/Y _11473_/X vssd1 vssd1 vccd1 vccd1
+ _11474_/X sky130_fd_sc_hd__a221o_1
XFILLER_137_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_100_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17676__B _17680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16001_ _13392_/B _16000_/X _14623_/A vssd1 vssd1 vccd1 vccd1 _16146_/A sky130_fd_sc_hd__a21o_2
XANTENNA__17829__A0 _19729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13213_ _19760_/Q _19761_/Q _13213_/C vssd1 vssd1 vccd1 vccd1 _13233_/B sky130_fd_sc_hd__and3_1
X_10425_ _10429_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10425_/Y sky130_fd_sc_hd__nor2_1
XFILLER_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14193_ _18607_/Q _14045_/X _14195_/S vssd1 vssd1 vccd1 vccd1 _14194_/A sky130_fd_sc_hd__mux2_1
X_13144_ _13142_/X _13143_/X _13144_/S vssd1 vssd1 vccd1 vccd1 _13144_/X sky130_fd_sc_hd__mux2_1
X_10356_ _19188_/Q _18802_/Q _19252_/Q _18371_/Q _10315_/S _10229_/X vssd1 vssd1 vccd1
+ vccd1 _10357_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10472__S0 _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13075_ _19566_/Q vssd1 vssd1 vccd1 vccd1 _16782_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17952_ _17952_/A vssd1 vssd1 vccd1 vccd1 _19750_/D sky130_fd_sc_hd__clkbuf_1
X_10287_ _19190_/Q _18804_/Q _19254_/Q _18373_/Q _10286_/X _10275_/X vssd1 vssd1 vccd1
+ vccd1 _10288_/B sky130_fd_sc_hd__mux4_1
XFILLER_97_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17057__A1 _12669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16903_ _16904_/A _16904_/C _16902_/Y vssd1 vssd1 vccd1 vccd1 _19613_/D sky130_fd_sc_hd__o21a_1
X_12026_ _12111_/A _12140_/B vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__nand2_1
XFILLER_120_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17883_ _12337_/Y _17786_/X _17882_/X _17795_/X vssd1 vssd1 vccd1 vccd1 _17883_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19622_ _19669_/CLK _19622_/D vssd1 vssd1 vccd1 vccd1 _19622_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15416__S _15422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16834_ _16836_/A _16836_/B _16812_/X vssd1 vssd1 vccd1 vccd1 _16834_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19553_ _19828_/CLK _19553_/D vssd1 vssd1 vccd1 vccd1 _19553_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16765_ _16772_/C _16772_/D _16764_/X vssd1 vssd1 vccd1 vccd1 _16765_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13977_ _13977_/A vssd1 vssd1 vccd1 vccd1 _18521_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18504_ _18902_/CLK _18504_/D vssd1 vssd1 vccd1 vccd1 _18504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15716_ _15716_/A vssd1 vssd1 vccd1 vccd1 _19203_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19484_ _19491_/CLK _19484_/D vssd1 vssd1 vccd1 vccd1 _19484_/Q sky130_fd_sc_hd__dfxtp_1
X_12928_ _19745_/Q _19746_/Q _12928_/C vssd1 vssd1 vccd1 vccd1 _12971_/B sky130_fd_sc_hd__and3_1
X_16696_ _16696_/A _16696_/B _16704_/D vssd1 vssd1 vccd1 vccd1 _19541_/D sky130_fd_sc_hd__nor3_1
XFILLER_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18435_ _19058_/CLK _18435_/D vssd1 vssd1 vccd1 vccd1 _18435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15647_ _14531_/X _19173_/Q _15649_/S vssd1 vssd1 vccd1 vccd1 _15648_/A sky130_fd_sc_hd__mux2_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _13114_/A vssd1 vssd1 vccd1 vccd1 _13345_/S sky130_fd_sc_hd__buf_2
XFILLER_34_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18366_ _19247_/CLK _18366_/D vssd1 vssd1 vccd1 vccd1 _18366_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11899__B _17205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15578_ _15576_/X _19158_/Q _15596_/S vssd1 vssd1 vccd1 vccd1 _15579_/A sky130_fd_sc_hd__mux2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10065__C1 _09811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17317_ _17317_/A _17462_/A vssd1 vssd1 vccd1 vccd1 _17317_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10604__A1 _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14529_ _14528_/X _18749_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14530_/A sky130_fd_sc_hd__mux2_1
XFILLER_147_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18297_ _18894_/CLK _18297_/D vssd1 vssd1 vccd1 vccd1 _18297_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16771__A _16848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15543__A1 _15542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17248_ _17587_/B _12286_/A _17274_/A vssd1 vssd1 vccd1 vccd1 _17346_/B sky130_fd_sc_hd__mux2_1
XFILLER_128_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12357__A1 _11416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17179_ _17240_/S vssd1 vssd1 vccd1 vccd1 _17274_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14291__A _14291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12804__A _19701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09222__B2 _09331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_103_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17048__A1 _15509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15326__S _15328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09908__S0 _10112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13354__B _17028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11155__A _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09504_ _10965_/A vssd1 vssd1 vccd1 vccd1 _10640_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17220__A1 _17779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09435_ _09390_/X _09407_/X _09420_/X _10514_/A _09726_/A vssd1 vssd1 vccd1 vccd1
+ _09452_/B sky130_fd_sc_hd__o221a_1
XFILLER_169_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13370__A _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09366_ _09366_/A vssd1 vssd1 vccd1 vccd1 _09367_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15996__S _15996_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09297_ _19626_/Q _19621_/Q vssd1 vssd1 vccd1 vccd1 _09297_/X sky130_fd_sc_hd__and2_1
XFILLER_123_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10359__B1 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12714__A _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _19287_/Q _19125_/Q _18534_/Q _18304_/Q _10166_/S _09954_/A vssd1 vssd1 vccd1
+ vccd1 _10210_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11190_ _11184_/A _11189_/X _10883_/X vssd1 vssd1 vccd1 vccd1 _11190_/X sky130_fd_sc_hd__o21a_1
XFILLER_161_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10141_ _10148_/A _10136_/X _10138_/X _10140_/X vssd1 vssd1 vccd1 vccd1 _10141_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17716__S _17716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17039__A1 _15481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_clock clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_82_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10206__S0 _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _19293_/Q _19131_/Q _18540_/Q _18310_/Q _09500_/A _09507_/A vssd1 vssd1 vccd1
+ vccd1 _10072_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13900_ _13899_/X _18499_/Q _13903_/S vssd1 vssd1 vccd1 vccd1 _13901_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14880_ _18888_/Q _13975_/X _14882_/S vssd1 vssd1 vccd1 vccd1 _14881_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13831_ _13349_/X _18478_/Q _13831_/S vssd1 vssd1 vccd1 vccd1 _13832_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13076__A2 _12703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16550_ _16551_/B _16551_/C _19497_/Q vssd1 vssd1 vccd1 vccd1 _16552_/B sky130_fd_sc_hd__a21oi_1
X_10974_ _10981_/A _10967_/X _10973_/X vssd1 vssd1 vccd1 vccd1 _10974_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13762_ _13386_/X _18448_/Q _13762_/S vssd1 vssd1 vccd1 vccd1 _13763_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15501_ _12544_/X _15499_/X _15500_/Y _15549_/A _18258_/Q vssd1 vssd1 vccd1 vccd1
+ _16919_/A sky130_fd_sc_hd__a32o_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12713_ _12713_/A _18275_/Q vssd1 vssd1 vccd1 vccd1 _12713_/Y sky130_fd_sc_hd__nand2_1
X_16481_ _16483_/B _16483_/C _16446_/X vssd1 vssd1 vccd1 vccd1 _16481_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_44_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13693_ _13749_/A vssd1 vssd1 vccd1 vccd1 _13762_/S sky130_fd_sc_hd__buf_6
XFILLER_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18220_ _18224_/A _18220_/B vssd1 vssd1 vccd1 vccd1 _18221_/A sky130_fd_sc_hd__and2_1
XFILLER_102_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15432_ _15432_/A vssd1 vssd1 vccd1 vccd1 _19122_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12644_ _13265_/A vssd1 vssd1 vccd1 vccd1 _12644_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12587__B2 _19474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18151_ _18151_/A vssd1 vssd1 vccd1 vccd1 _19835_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11512__B _11512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12575_ _12714_/A vssd1 vssd1 vccd1 vccd1 _12575_/X sky130_fd_sc_hd__clkbuf_2
X_15363_ _15374_/A vssd1 vssd1 vccd1 vccd1 _15372_/S sky130_fd_sc_hd__buf_4
XFILLER_50_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17102_ _17102_/A _17102_/B vssd1 vssd1 vccd1 vccd1 _17163_/A sky130_fd_sc_hd__and2_2
XFILLER_50_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14314_ _14314_/A vssd1 vssd1 vccd1 vccd1 _18651_/D sky130_fd_sc_hd__clkbuf_1
X_18082_ _19808_/Q _12627_/X _18081_/X _17021_/X vssd1 vssd1 vccd1 vccd1 _19808_/D
+ sky130_fd_sc_hd__o211a_1
X_11526_ _11526_/A vssd1 vssd1 vccd1 vccd1 _12475_/A sky130_fd_sc_hd__clkbuf_2
X_15294_ _14589_/X _19061_/Q _15300_/S vssd1 vssd1 vccd1 vccd1 _15295_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17033_ _19665_/Q _13410_/X _17039_/S vssd1 vssd1 vccd1 vccd1 _17034_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14245_ _18629_/Q _14013_/X _14253_/S vssd1 vssd1 vccd1 vccd1 _14246_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09204__A1 _18109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _11460_/A _11462_/A _11459_/B _10751_/A vssd1 vssd1 vccd1 vccd1 _11457_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12624__A _17133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ _19283_/Q _19121_/Q _18530_/Q _18300_/Q _10451_/S _10311_/A vssd1 vssd1 vccd1
+ vccd1 _10409_/B sky130_fd_sc_hd__mux4_1
XANTENNA__15000__A _15099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14176_ _18599_/Q _14020_/X _14180_/S vssd1 vssd1 vccd1 vccd1 _14177_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11388_ _18640_/Q _18975_/Q _11388_/S vssd1 vssd1 vccd1 vccd1 _11389_/B sky130_fd_sc_hd__mux2_1
XANTENNA_output89_A _12317_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10339_ _18500_/Q _18995_/Q _10339_/S vssd1 vssd1 vccd1 vccd1 _10340_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10996__S1 _10990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13127_ _19756_/Q _13127_/B vssd1 vssd1 vccd1 vccd1 _13152_/C sky130_fd_sc_hd__and2_1
XFILLER_152_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _19367_/CLK _18984_/D vssd1 vssd1 vccd1 vccd1 _18984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_124_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _19565_/Q _13055_/X _13057_/X _13012_/X vssd1 vssd1 vccd1 vccd1 _13058_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _16011_/B _19775_/Q _17935_/S vssd1 vssd1 vccd1 vccd1 _17936_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12009_ _12392_/S _12009_/B vssd1 vssd1 vccd1 vccd1 _12009_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09912__C1 _09813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17866_ _17864_/X _17865_/Y _17898_/S vssd1 vssd1 vccd1 vccd1 _17866_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10798__B _12454_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16817_ _16838_/A _16817_/B _16821_/C vssd1 vssd1 vccd1 vccd1 _19578_/D sky130_fd_sc_hd__nor3_1
X_19605_ _19607_/CLK _19605_/D vssd1 vssd1 vccd1 vccd1 _19605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_94_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15461__A0 _09309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17797_ _19726_/Q _17570_/X _17796_/X vssd1 vssd1 vccd1 vccd1 _19726_/D sky130_fd_sc_hd__o21a_1
XFILLER_81_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19536_ _19540_/CLK _19536_/D vssd1 vssd1 vccd1 vccd1 _19536_/Q sky130_fd_sc_hd__dfxtp_1
X_16748_ _19559_/Q _19558_/Q _19555_/Q _19554_/Q vssd1 vssd1 vccd1 vccd1 _16750_/C
+ sky130_fd_sc_hd__and4_1
X_19467_ _19603_/CLK _19467_/D vssd1 vssd1 vccd1 vccd1 _19467_/Q sky130_fd_sc_hd__dfxtp_1
X_16679_ _19535_/Q _19534_/Q _19533_/Q _16679_/D vssd1 vssd1 vccd1 vccd1 _16687_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_62_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13190__A _15063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ _19858_/Q vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__buf_2
X_18418_ _19203_/CLK _18418_/D vssd1 vssd1 vccd1 vccd1 _18418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19398_ _19838_/CLK _19398_/D vssd1 vssd1 vccd1 vccd1 _19398_/Q sky130_fd_sc_hd__dfxtp_1
X_09151_ _09158_/B vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18349_ _19264_/CLK _18349_/D vssd1 vssd1 vccd1 vccd1 _18349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15516__A1 _15515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11250__A1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ _09146_/C _09180_/C vssd1 vssd1 vccd1 vccd1 _17121_/A sky130_fd_sc_hd__or2_4
XFILLER_174_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18205__B _18205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput60 io_ibus_inst[4] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__14225__S _14231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12750__A1 _18263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09984_ _09672_/A _09980_/X _09983_/X vssd1 vssd1 vccd1 vccd1 _09984_/X sky130_fd_sc_hd__a21o_1
XFILLER_107_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_169_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__A _14272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10911__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09418_ _09590_/A vssd1 vssd1 vccd1 vccd1 _09419_/A sky130_fd_sc_hd__buf_4
XFILLER_80_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10690_ _18492_/Q _18987_/Q _11320_/S vssd1 vssd1 vccd1 vccd1 _10691_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09349_ _19863_/Q vssd1 vssd1 vccd1 vccd1 _18140_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10229__A _10229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _12360_/A _17885_/B vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__or2_1
XFILLER_154_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_126_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ _09597_/X _11310_/X _09608_/A vssd1 vssd1 vccd1 vccd1 _11311_/X sky130_fd_sc_hd__o21a_1
XFILLER_138_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10595__A3 _10593_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ _12312_/B _12291_/B vssd1 vssd1 vccd1 vccd1 _12291_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14030_ _14030_/A vssd1 vssd1 vccd1 vccd1 _14043_/S sky130_fd_sc_hd__clkbuf_4
X_11242_ _11242_/A _11242_/B vssd1 vssd1 vccd1 vccd1 _11242_/X sky130_fd_sc_hd__and2_1
XANTENNA__12741__A1 hold19/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11173_ _18612_/Q _18947_/Q _11173_/S vssd1 vssd1 vccd1 vccd1 _11174_/B sky130_fd_sc_hd__mux2_1
XFILLER_164_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input40_A io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__A _09753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _19193_/Q _18807_/Q _19257_/Q _18376_/Q _09786_/A _10169_/A vssd1 vssd1 vccd1
+ vccd1 _10125_/B sky130_fd_sc_hd__mux4_1
XFILLER_164_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15981_ _13592_/X _19322_/Q _15981_/S vssd1 vssd1 vccd1 vccd1 _15982_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17720_ _11339_/Y _17652_/X _17719_/X vssd1 vssd1 vccd1 vccd1 _19720_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__13275__A _13275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14932_ _18912_/Q vssd1 vssd1 vccd1 vccd1 _14933_/A sky130_fd_sc_hd__clkbuf_1
X_10055_ _18636_/Q _18971_/Q _10055_/S vssd1 vssd1 vccd1 vccd1 _10056_/B sky130_fd_sc_hd__mux2_1
XFILLER_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17651_ _10795_/Y _12773_/X _17650_/X vssd1 vssd1 vccd1 vccd1 _19716_/D sky130_fd_sc_hd__a21oi_1
X_14863_ _18880_/Q _13943_/X _14871_/S vssd1 vssd1 vccd1 vccd1 _14864_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16602_ _19514_/Q _16604_/C _16601_/Y vssd1 vssd1 vccd1 vccd1 _19514_/D sky130_fd_sc_hd__o21a_1
XANTENNA__15490__A _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09899__S _10168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13814_ _13209_/X _18470_/Q _13820_/S vssd1 vssd1 vccd1 vccd1 _13815_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17582_ _17587_/A _17587_/B _17832_/S vssd1 vssd1 vccd1 vccd1 _17582_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14794_ _14794_/A vssd1 vssd1 vccd1 vccd1 _18849_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19321_ _19383_/CLK _19321_/D vssd1 vssd1 vccd1 vccd1 _19321_/Q sky130_fd_sc_hd__dfxtp_1
X_16533_ _19492_/Q _19491_/Q _19490_/Q _16533_/D vssd1 vssd1 vccd1 vccd1 _16542_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13745_ _13240_/X _18440_/Q _13747_/S vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ _10953_/A _10954_/X _10956_/X _09448_/A vssd1 vssd1 vccd1 vccd1 _10957_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12619__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11523__A _18087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19252_ _19378_/CLK _19252_/D vssd1 vssd1 vccd1 vccd1 _19252_/Q sky130_fd_sc_hd__dfxtp_1
X_16464_ _16466_/B _16466_/C _16446_/X vssd1 vssd1 vccd1 vccd1 _16464_/Y sky130_fd_sc_hd__a21oi_1
X_13676_ _13676_/A vssd1 vssd1 vccd1 vccd1 _18409_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10888_ _19305_/Q _18717_/Q _18754_/Q _18328_/Q _11172_/S _11174_/A vssd1 vssd1 vccd1
+ vccd1 _10889_/B sky130_fd_sc_hd__mux4_1
X_18203_ _18203_/A vssd1 vssd1 vccd1 vccd1 _19849_/D sky130_fd_sc_hd__clkbuf_1
X_15415_ _15415_/A vssd1 vssd1 vccd1 vccd1 _19114_/D sky130_fd_sc_hd__clkbuf_1
X_12627_ _18134_/A vssd1 vssd1 vccd1 vccd1 _12627_/X sky130_fd_sc_hd__clkbuf_2
X_19183_ _19247_/CLK _19183_/D vssd1 vssd1 vccd1 vccd1 _19183_/Q sky130_fd_sc_hd__dfxtp_1
X_16395_ _19447_/Q _16396_/C _19448_/Q vssd1 vssd1 vccd1 vccd1 _16397_/B sky130_fd_sc_hd__a21oi_1
XFILLER_169_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16752__C _19557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18134_ _18134_/A vssd1 vssd1 vccd1 vccd1 _18134_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10666__S0 _10650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ _19084_/Q _15038_/X _15350_/S vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__mux2_1
X_12558_ _19537_/Q vssd1 vssd1 vccd1 vccd1 _16689_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_18065_ _18065_/A vssd1 vssd1 vccd1 vccd1 _19801_/D sky130_fd_sc_hd__clkbuf_1
X_11509_ _11516_/A _12322_/B vssd1 vssd1 vccd1 vccd1 _11510_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15277_ _15277_/A vssd1 vssd1 vccd1 vccd1 _19053_/D sky130_fd_sc_hd__clkbuf_1
X_12489_ _12660_/B vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__buf_2
XFILLER_144_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17016_ _19659_/Q _17024_/B vssd1 vssd1 vccd1 vccd1 _17016_/X sky130_fd_sc_hd__or2_1
XFILLER_132_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14228_ _14228_/A vssd1 vssd1 vccd1 vccd1 _18621_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12732__A1 _11677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _14159_/A vssd1 vssd1 vccd1 vccd1 _18591_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18041__A _18188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18967_ _19127_/CLK _18967_/D vssd1 vssd1 vccd1 vccd1 _18967_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17918_ _17534_/A _17232_/A _17462_/A _17917_/X vssd1 vssd1 vccd1 vccd1 _17918_/X
+ sky130_fd_sc_hd__o211a_1
X_18898_ _19284_/CLK _18898_/D vssd1 vssd1 vccd1 vccd1 _18898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09361__B1 _09360_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17849_ _17434_/X _17599_/Y _17848_/X _17473_/X vssd1 vssd1 vccd1 vccd1 _17849_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12799__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19519_ _19550_/CLK _19519_/D vssd1 vssd1 vccd1 vccd1 _19519_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12799__B2 _12798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_170_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _19853_/Q _14197_/B vssd1 vssd1 vccd1 vccd1 _09203_/Y sky130_fd_sc_hd__xnor2_1
X_09134_ _09176_/A _11569_/A _09134_/C vssd1 vssd1 vccd1 vccd1 _11575_/A sky130_fd_sc_hd__and3_1
XFILLER_135_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10329__A3 _10328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13794__S _13798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15575__A _15601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_95_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09967_ _18473_/Q _19064_/Q _19226_/Q _18441_/Q _09782_/A _09773_/A vssd1 vssd1 vccd1
+ vccd1 _09968_/B sky130_fd_sc_hd__mux4_1
XFILLER_58_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17790__A _17790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09898_ _10217_/S vssd1 vssd1 vccd1 vccd1 _10168_/S sky130_fd_sc_hd__clkbuf_4
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11860_ _19336_/Q _11859_/X _15488_/A vssd1 vssd1 vccd1 vccd1 _11860_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11137__S1 _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10811_ _18781_/Q vssd1 vssd1 vccd1 vccd1 _11252_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11791_ _11791_/A _11791_/B vssd1 vssd1 vccd1 vccd1 _11796_/A sky130_fd_sc_hd__xor2_4
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13530_ _13530_/A vssd1 vssd1 vccd1 vccd1 _18357_/D sky130_fd_sc_hd__clkbuf_1
X_10742_ _18459_/Q _19050_/Q _19212_/Q _18427_/Q _11297_/S _09600_/A vssd1 vssd1 vccd1
+ vccd1 _10743_/B sky130_fd_sc_hd__mux4_1
XFILLER_40_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13739__A0 _13191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13461_ _13507_/S vssd1 vssd1 vccd1 vccd1 _13470_/S sky130_fd_sc_hd__buf_2
X_10673_ _11305_/A vssd1 vssd1 vccd1 vccd1 _11309_/A sky130_fd_sc_hd__buf_2
XANTENNA__09407__A1 _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _19019_/Q _15035_/X _15206_/S vssd1 vssd1 vccd1 vccd1 _15201_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12412_ _12435_/A _12408_/X _12411_/X vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__11214__A1 _09366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16180_ _13528_/X _19364_/Q _16180_/S vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11214__B2 _19708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13392_ _13392_/A _13392_/B vssd1 vssd1 vccd1 vccd1 _15463_/A sky130_fd_sc_hd__nand2_1
XFILLER_139_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10422__C1 _09669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15131_ _15131_/A vssd1 vssd1 vccd1 vccd1 _18988_/D sky130_fd_sc_hd__clkbuf_1
X_12343_ _19658_/Q _19657_/Q _12343_/C vssd1 vssd1 vccd1 vccd1 _12394_/C sky130_fd_sc_hd__and3_1
XANTENNA__10973__B1 _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15062_ _15062_/A vssd1 vssd1 vccd1 vccd1 _18963_/D sky130_fd_sc_hd__clkbuf_1
X_12274_ _19352_/Q _12274_/B vssd1 vssd1 vccd1 vccd1 _12274_/X sky130_fd_sc_hd__or2_1
XFILLER_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14013_ _14585_/A vssd1 vssd1 vccd1 vccd1 _14013_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15485__A hold19/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ _11228_/A _11222_/X _11224_/X vssd1 vssd1 vccd1 vccd1 _11225_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09483__A _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11156_ _18580_/Q _18851_/Q _19075_/Q _18819_/Q _09496_/A _11100_/A vssd1 vssd1 vccd1
+ vccd1 _11156_/X sky130_fd_sc_hd__mux4_1
X_18821_ _19271_/CLK _18821_/D vssd1 vssd1 vccd1 vccd1 _18821_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12621__B _12621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10107_ _19289_/Q _19127_/Q _18536_/Q _18306_/Q _10185_/S _09714_/A vssd1 vssd1 vccd1
+ vccd1 _10108_/B sky130_fd_sc_hd__mux4_1
XANTENNA__11518__A _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18752_ _19239_/CLK _18752_/D vssd1 vssd1 vccd1 vccd1 _18752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15964_ _13567_/X _19314_/Q _15970_/S vssd1 vssd1 vccd1 vccd1 _15965_/A sky130_fd_sc_hd__mux2_1
X_11087_ _11026_/A _11086_/X _11022_/X vssd1 vssd1 vccd1 vccd1 _11087_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_48_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17703_ _17871_/A _17703_/B vssd1 vssd1 vccd1 vccd1 _17703_/X sky130_fd_sc_hd__or2_1
X_14915_ _18904_/Q _14026_/X _14915_/S vssd1 vssd1 vccd1 vccd1 _14916_/A sky130_fd_sc_hd__mux2_1
X_10038_ _10667_/A _10038_/B vssd1 vssd1 vccd1 vccd1 _10038_/X sky130_fd_sc_hd__or2_1
XFILLER_64_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18683_ _19365_/CLK _18683_/D vssd1 vssd1 vccd1 vccd1 _18683_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15895_ _15895_/A vssd1 vssd1 vccd1 vccd1 _19283_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17634_ _17390_/A _17625_/X _17632_/X _17633_/X vssd1 vssd1 vccd1 vccd1 _17634_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17205__A _17205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14846_ _18873_/Q _14029_/X _14854_/S vssd1 vssd1 vccd1 vccd1 _14847_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _17413_/X _17562_/X _17564_/Y _17532_/X vssd1 vssd1 vccd1 vccd1 _17565_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14777_ _14608_/X _18843_/Q _14781_/S vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__mux2_1
X_11989_ _19405_/Q vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12349__A _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19304_ _19306_/CLK _19304_/D vssd1 vssd1 vccd1 vccd1 _19304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16516_ _19613_/Q _19615_/Q _19614_/Q _16899_/A vssd1 vssd1 vccd1 vccd1 _16907_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13728_ _13107_/X _18432_/Q _13736_/S vssd1 vssd1 vccd1 vccd1 _13729_/A sky130_fd_sc_hd__mux2_1
XFILLER_149_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _17478_/X _17484_/Y _17495_/X _17422_/A vssd1 vssd1 vccd1 vccd1 _17496_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_32_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19235_ _19235_/CLK _19235_/D vssd1 vssd1 vccd1 vccd1 _19235_/Q sky130_fd_sc_hd__dfxtp_1
X_16447_ _16450_/B _16450_/C _16446_/X vssd1 vssd1 vccd1 vccd1 _16447_/Y sky130_fd_sc_hd__a21oi_1
X_13659_ _13659_/A vssd1 vssd1 vccd1 vccd1 _18401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ _19598_/CLK _19166_/D vssd1 vssd1 vccd1 vccd1 _19166_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09658__A _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16378_ _19441_/Q _16379_/C _19442_/Q vssd1 vssd1 vccd1 vccd1 _16380_/B sky130_fd_sc_hd__a21oi_1
XFILLER_157_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18117_ _19822_/Q _18106_/X _18116_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _19822_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15329_ _15329_/A vssd1 vssd1 vccd1 vccd1 _19076_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12084__A _17768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19097_ _19385_/CLK _19097_/D vssd1 vssd1 vccd1 vccd1 _19097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18048_ _19794_/Q _19415_/Q _18050_/S vssd1 vssd1 vccd1 vccd1 _18049_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_117_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12812__A _13387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14503__S _14511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09821_ _09821_/A vssd1 vssd1 vccd1 vccd1 _09822_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09393__A _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10192__A1 _10195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09752_ _09752_/A vssd1 vssd1 vccd1 vccd1 _09753_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_100_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09683_ _10186_/S vssd1 vssd1 vccd1 vccd1 _10185_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__15407__A0 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14739__A _14785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11692__A1 _11686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19310_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11610__B _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09117_ _09328_/A vssd1 vssd1 vccd1 vccd1 _18104_/A sky130_fd_sc_hd__inv_2
XFILLER_164_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17883__A1 _12337_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14413__S _14417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11010_ _11064_/A _11010_/B vssd1 vssd1 vccd1 vccd1 _11010_/X sky130_fd_sc_hd__or2_1
XFILLER_132_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13121__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _16760_/B _12518_/A _12565_/A _16963_/A _13012_/A vssd1 vssd1 vccd1 vccd1
+ _12961_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14700_ _14700_/A vssd1 vssd1 vccd1 vccd1 _14709_/S sky130_fd_sc_hd__buf_6
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _19641_/Q vssd1 vssd1 vccd1 vccd1 _16967_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15680_ _14579_/X _19188_/Q _15682_/S vssd1 vssd1 vccd1 vccd1 _15681_/A sky130_fd_sc_hd__mux2_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12892_ _12892_/A _12928_/C vssd1 vssd1 vccd1 vccd1 _12892_/Y sky130_fd_sc_hd__nor2_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14631_ input42/X _18148_/A _14293_/X _14623_/X _18112_/A vssd1 vssd1 vccd1 vccd1
+ _18209_/B sky130_fd_sc_hd__a32o_2
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _11949_/A _11950_/A vssd1 vssd1 vccd1 vccd1 _11844_/B sky130_fd_sc_hd__nand2_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17350_ _17609_/A _17350_/B vssd1 vssd1 vccd1 vccd1 _17350_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12632__B1 _18234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ _14562_/A vssd1 vssd1 vccd1 vccd1 _18759_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _13419_/A _16951_/A vssd1 vssd1 vccd1 vccd1 _11774_/X sky130_fd_sc_hd__and2b_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16301_/A vssd1 vssd1 vccd1 vccd1 _18170_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _19701_/Q _16000_/B _14998_/A vssd1 vssd1 vccd1 vccd1 _14860_/D sky130_fd_sc_hd__and3_1
XFILLER_14_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13699__S _13703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17281_ _17269_/X _17279_/X _17613_/A vssd1 vssd1 vccd1 vccd1 _17281_/X sky130_fd_sc_hd__mux2_1
X_10725_ _10710_/X _10715_/X _10724_/X _09571_/A vssd1 vssd1 vccd1 vccd1 _10725_/X
+ sky130_fd_sc_hd__a22o_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14493_ _14493_/A vssd1 vssd1 vccd1 vccd1 _18730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19020_ _19086_/CLK _19020_/D vssd1 vssd1 vccd1 vccd1 _19020_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13188__A1 input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16232_ _16232_/A vssd1 vssd1 vccd1 vccd1 _19387_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13444_ _12851_/X _18323_/Q _13448_/S vssd1 vssd1 vccd1 vccd1 _13445_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10656_ _19309_/Q _18721_/Q _18758_/Q _18332_/Q _10729_/S _10655_/X vssd1 vssd1 vccd1
+ vccd1 _10656_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ _16162_/X _19358_/Q _16167_/S vssd1 vssd1 vccd1 vccd1 _16164_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11520__B _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13375_ _19695_/Q _13008_/X _13009_/X _19662_/Q vssd1 vssd1 vccd1 vccd1 _13375_/X
+ sky130_fd_sc_hd__a22o_1
X_10587_ _19312_/Q _18724_/Q _18761_/Q _18335_/Q _10566_/X _10586_/X vssd1 vssd1 vccd1
+ vccd1 _10587_/X sky130_fd_sc_hd__mux4_1
XFILLER_154_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15114_ _15171_/S vssd1 vssd1 vccd1 vccd1 _15123_/S sky130_fd_sc_hd__buf_2
X_12326_ _19657_/Q _12343_/C vssd1 vssd1 vccd1 vccd1 _12326_/X sky130_fd_sc_hd__and2_1
XFILLER_86_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16094_ _12233_/X _12593_/B _16093_/Y vssd1 vssd1 vccd1 vccd1 _16094_/X sky130_fd_sc_hd__a21o_1
XFILLER_114_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15045_ _18958_/Q _15044_/X _15045_/S vssd1 vssd1 vccd1 vccd1 _15046_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ _19654_/Q _12235_/X _11773_/X vssd1 vssd1 vccd1 vccd1 _12257_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output71_A _12488_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13360__A1 _13359_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__B1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _11208_/A _11208_/B vssd1 vssd1 vccd1 vccd1 _11208_/X sky130_fd_sc_hd__or2_1
X_19853_ _19854_/CLK _19853_/D vssd1 vssd1 vccd1 vccd1 _19853_/Q sky130_fd_sc_hd__dfxtp_1
X_12188_ _09331_/A _11507_/A _12209_/A vssd1 vssd1 vccd1 vccd1 _12188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_69_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10713__A3 _18826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18804_ _19319_/CLK _18804_/D vssd1 vssd1 vccd1 vccd1 _18804_/Q sky130_fd_sc_hd__dfxtp_1
X_11139_ _19300_/Q _18712_/Q _18749_/Q _18323_/Q _11173_/S _11124_/X vssd1 vssd1 vccd1
+ vccd1 _11140_/B sky130_fd_sc_hd__mux4_1
X_16996_ _15574_/X _16983_/X _16993_/X _16995_/X vssd1 vssd1 vccd1 vccd1 _19651_/D
+ sky130_fd_sc_hd__o211a_1
X_19784_ _19786_/CLK _19784_/D vssd1 vssd1 vccd1 vccd1 _19784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15947_ _15947_/A vssd1 vssd1 vccd1 vccd1 _19306_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18735_ _19291_/CLK _18735_/D vssd1 vssd1 vccd1 vccd1 _18735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15154__S _15156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18666_ _19089_/CLK _18666_/D vssd1 vssd1 vccd1 vccd1 _18666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10021__S1 _10056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15878_ _15924_/S vssd1 vssd1 vccd1 vccd1 _15887_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_63_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14829_ _14829_/A vssd1 vssd1 vccd1 vccd1 _18865_/D sky130_fd_sc_hd__clkbuf_1
X_17617_ _17654_/A _17614_/Y _17616_/X vssd1 vssd1 vccd1 vccd1 _17617_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18597_ _19286_/CLK _18597_/D vssd1 vssd1 vccd1 vccd1 _18597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17548_ _17613_/A _17548_/B vssd1 vssd1 vccd1 vccd1 _17548_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_43_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11977__A2 _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17479_ _17732_/S vssd1 vssd1 vccd1 vccd1 _17479_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14376__A0 _13837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19218_ _19314_/CLK _19218_/D vssd1 vssd1 vccd1 vccd1 _19218_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09388__A _10030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19149_ _19687_/CLK _19149_/D vssd1 vssd1 vccd1 vccd1 _19149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09804_ _10471_/A vssd1 vssd1 vccd1 vccd1 _10335_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09307__B1 _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13103__A1 _15546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15572__B _15572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _18413_/Q _18674_/Q _18573_/Q _18908_/Q _09743_/A _09733_/A vssd1 vssd1 vccd1
+ vccd1 _09736_/B sky130_fd_sc_hd__mux4_1
XFILLER_86_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11114__B1 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14469__A _14515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18042__A1 _19412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_153_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19205_/CLK sky130_fd_sc_hd__clkbuf_16
X_09666_ _09666_/A vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15800__A0 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09597_ _10547_/A vssd1 vssd1 vccd1 vccd1 _09597_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_168_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19297_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10936__S _11196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11621__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13312__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ _19313_/Q _18725_/Q _18762_/Q _18336_/Q _10496_/X _09710_/A vssd1 vssd1 vccd1
+ vccd1 _10511_/B sky130_fd_sc_hd__mux4_1
XFILLER_11_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11490_ _11491_/B _17121_/B vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__or2_1
XFILLER_168_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _18594_/Q _18865_/Q _19089_/Q _18833_/Q _10435_/S _10348_/A vssd1 vssd1 vccd1
+ vccd1 _10441_/X sky130_fd_sc_hd__mux4_1
XFILLER_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13160_ _19443_/Q _12515_/X _13159_/X vssd1 vssd1 vccd1 vccd1 _13160_/X sky130_fd_sc_hd__o21a_1
X_10372_ _18403_/Q _18664_/Q _18563_/Q _18898_/Q _10413_/S _10229_/A vssd1 vssd1 vccd1
+ vccd1 _10373_/B sky130_fd_sc_hd__mux4_1
XFILLER_40_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12111_ _12111_/A vssd1 vssd1 vccd1 vccd1 _12305_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15239__S _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13091_ _13090_/X _18297_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13092_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13548__A _13615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12042_ _19343_/Q _11859_/X _12037_/X _12041_/X _12230_/A vssd1 vssd1 vccd1 vccd1
+ _12042_/X sky130_fd_sc_hd__o221a_1
XFILLER_46_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_106_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19564_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_172_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10156__A1 _09667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10156__B2 _19729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15619__A0 _13325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16850_ _16883_/A _16854_/C vssd1 vssd1 vccd1 vccd1 _16850_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10251__S1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15801_ _15801_/A vssd1 vssd1 vccd1 vccd1 _19241_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16781_ _16777_/Y _16778_/Y _16788_/D _16293_/X vssd1 vssd1 vccd1 vccd1 _19567_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13993_ _13993_/A vssd1 vssd1 vccd1 vccd1 _18526_/D sky130_fd_sc_hd__clkbuf_1
X_18520_ _19367_/CLK _18520_/D vssd1 vssd1 vccd1 vccd1 _18520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15732_ _13544_/X _19211_/Q _15732_/S vssd1 vssd1 vccd1 vccd1 _15733_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11200__S0 _11128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ _15022_/A vssd1 vssd1 vccd1 vccd1 _14544_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10003__S1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09944__S1 _09714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18451_ _19300_/CLK _18451_/D vssd1 vssd1 vccd1 vccd1 _18451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15663_ _14553_/X _19180_/Q _15671_/S vssd1 vssd1 vccd1 vccd1 _15664_/A sky130_fd_sc_hd__mux2_1
X_12875_ _19668_/Q _12703_/X _12521_/A _16951_/A vssd1 vssd1 vccd1 vccd1 _12875_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16594__A _16806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17402_/A vssd1 vssd1 vccd1 vccd1 _17402_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15702__S _15704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__A1 _09831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14614_ _14614_/A vssd1 vssd1 vccd1 vccd1 _14614_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _11826_/A _19399_/Q _12098_/C vssd1 vssd1 vccd1 vccd1 _11879_/C sky130_fd_sc_hd__and3_1
X_18382_ _19389_/CLK _18382_/D vssd1 vssd1 vccd1 vccd1 _18382_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15594_ _15594_/A vssd1 vssd1 vccd1 vccd1 _19161_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17333_ _17646_/A vssd1 vssd1 vccd1 vccd1 _17333_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14545_ _14544_/X _18754_/Q _14551_/S vssd1 vssd1 vccd1 vccd1 _14546_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12081__A1 _18112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _11717_/A _11782_/B _12050_/A vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__a21o_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17264_ _17790_/B _17696_/B _17283_/S vssd1 vssd1 vccd1 vccd1 _17264_/X sky130_fd_sc_hd__mux2_1
X_10708_ _18922_/Q _18688_/Q _19370_/Q _19018_/Q _10704_/S _10623_/A vssd1 vssd1 vccd1
+ vccd1 _10709_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14476_ _13883_/X _18723_/Q _14478_/S vssd1 vssd1 vccd1 vccd1 _14477_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11688_ _11687_/X _11683_/X _12179_/B vssd1 vssd1 vccd1 vccd1 _11688_/X sky130_fd_sc_hd__mux2_1
X_19003_ _19035_/CLK _19003_/D vssd1 vssd1 vccd1 vccd1 _19003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16215_ _16226_/A vssd1 vssd1 vccd1 vccd1 _16224_/S sky130_fd_sc_hd__buf_6
XFILLER_146_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ hold4/A _13380_/X _13426_/Y _15565_/A vssd1 vssd1 vccd1 vccd1 _13427_/X sky130_fd_sc_hd__o211a_1
XFILLER_174_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17195_ _17195_/A vssd1 vssd1 vccd1 vccd1 _17642_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_10639_ _10719_/A vssd1 vssd1 vccd1 vccd1 _10639_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16146_ _16146_/A vssd1 vssd1 vccd1 vccd1 _16167_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13358_ _19618_/Q _12697_/X _12507_/X _19550_/Q _13357_/X vssd1 vssd1 vccd1 vccd1
+ _13358_/X sky130_fd_sc_hd__a221o_1
XFILLER_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12309_ _12309_/A vssd1 vssd1 vccd1 vccd1 _17867_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_170_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ _16076_/X _19343_/Q _16083_/S vssd1 vssd1 vccd1 vccd1 _16078_/A sky130_fd_sc_hd__mux2_1
X_13289_ _19614_/Q _13260_/X _13261_/X _19482_/Q _13288_/X vssd1 vssd1 vccd1 vccd1
+ _15606_/B sky130_fd_sc_hd__a221o_4
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13333__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15028_ _15028_/A vssd1 vssd1 vccd1 vccd1 _15028_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16769__A _16778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15673__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19836_ _19838_/CLK _19836_/D vssd1 vssd1 vccd1 vccd1 _19836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_70_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19096_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold11_A hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09671__A _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15625__A3 _09234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19767_ _19793_/CLK _19767_/D vssd1 vssd1 vccd1 vccd1 _19767_/Q sky130_fd_sc_hd__dfxtp_1
X_16979_ _15542_/X _16970_/X _16978_/X _16968_/X vssd1 vssd1 vccd1 vccd1 _19645_/D
+ sky130_fd_sc_hd__o211a_1
Xinput3 io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_110_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09520_ _18510_/Q _19005_/Q _10017_/S vssd1 vssd1 vccd1 vccd1 _09521_/A sky130_fd_sc_hd__mux2_1
X_18718_ _19307_/CLK _18718_/D vssd1 vssd1 vccd1 vccd1 _18718_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12844__A0 _19709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19698_ _19866_/CLK _19698_/D vssd1 vssd1 vccd1 vccd1 _19698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09451_ _09998_/A _09439_/X _09445_/X _09737_/A vssd1 vssd1 vccd1 vccd1 _09452_/C
+ sky130_fd_sc_hd__o211a_1
X_18649_ _19300_/CLK _18649_/D vssd1 vssd1 vccd1 vccd1 _18649_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_85_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19687_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_80_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09382_ _18779_/Q vssd1 vssd1 vccd1 vccd1 _11011_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12072__A1 _19344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19328_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_145_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_161_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14898__S _14904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_38_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19375_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11616__A _16000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _09993_/A vssd1 vssd1 vccd1 vccd1 _10509_/A sky130_fd_sc_hd__buf_2
X_10990_ _10990_/A _10990_/B vssd1 vssd1 vccd1 vccd1 _10990_/X sky130_fd_sc_hd__and2_1
XFILLER_56_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09649_ _10579_/A vssd1 vssd1 vccd1 vccd1 _10785_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_76_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12660_ _19587_/Q _12660_/B vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__and2_1
XFILLER_150_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18118__B _18142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09520__S _10017_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11611_ _11611_/A vssd1 vssd1 vccd1 vccd1 _17317_/A sky130_fd_sc_hd__buf_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12591_ _15599_/A _18269_/Q vssd1 vssd1 vccd1 vccd1 _12591_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11351__A _11351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14330_ _13883_/X _18659_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14331_/A sky130_fd_sc_hd__mux2_1
X_11542_ _11542_/A vssd1 vssd1 vccd1 vccd1 _12450_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15001__A1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12166__B _17202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14261_ _14261_/A vssd1 vssd1 vccd1 vccd1 _18636_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11473_ _11449_/X _11451_/Y _11452_/Y _11454_/Y _11472_/X vssd1 vssd1 vccd1 vccd1
+ _11473_/X sky130_fd_sc_hd__a2111o_1
XFILLER_13_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16000_ _18746_/Q _16000_/B vssd1 vssd1 vccd1 vccd1 _16000_/X sky130_fd_sc_hd__or2_1
XFILLER_7_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13212_ _13195_/X _13213_/C _19761_/Q vssd1 vssd1 vccd1 vccd1 _13214_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_input70_A reset vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17829__A1 _17828_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _19187_/Q _18801_/Q _19251_/Q _18370_/Q _10381_/S _09886_/A vssd1 vssd1 vccd1
+ vccd1 _10425_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09756__A _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14192_ _14192_/A vssd1 vssd1 vccd1 vccd1 _18606_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09862__S0 _09846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13143_ _19725_/Q _12590_/B _13143_/S vssd1 vssd1 vccd1 vccd1 _13143_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10355_ _11351_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _11441_/A sky130_fd_sc_hd__or2_1
XFILLER_98_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13074_ _19534_/Q vssd1 vssd1 vccd1 vccd1 _16681_/C sky130_fd_sc_hd__clkbuf_2
X_10286_ _10435_/S vssd1 vssd1 vccd1 vccd1 _10286_/X sky130_fd_sc_hd__buf_4
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17951_ _16055_/A _19782_/Q _17957_/S vssd1 vssd1 vccd1 vccd1 _17952_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output157_A _16295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16902_ _16904_/A _16904_/C _16868_/X vssd1 vssd1 vccd1 vccd1 _16902_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__15493__A hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12025_ _12025_/A _12025_/B _12025_/C _17722_/A vssd1 vssd1 vccd1 vccd1 _12140_/B
+ sky130_fd_sc_hd__or4_2
X_17882_ _17852_/X _17529_/Y _17881_/X _17860_/X vssd1 vssd1 vccd1 vccd1 _17882_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19621_ _19669_/CLK _19621_/D vssd1 vssd1 vccd1 vccd1 _19621_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16833_ _16833_/A _16836_/A vssd1 vssd1 vccd1 vccd1 _19588_/D sky130_fd_sc_hd__nor2_1
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19552_ _19564_/CLK _19552_/D vssd1 vssd1 vccd1 vccd1 _19552_/Q sky130_fd_sc_hd__dfxtp_1
X_16764_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16764_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12826__B1 _12825_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13976_ _18521_/Q _13975_/X _13979_/S vssd1 vssd1 vccd1 vccd1 _13977_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18503_ _19088_/CLK _18503_/D vssd1 vssd1 vccd1 vccd1 _18503_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15715_ _13519_/X _19203_/Q _15721_/S vssd1 vssd1 vccd1 vccd1 _15716_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12927_ _16021_/B _12928_/C _19746_/Q vssd1 vssd1 vccd1 vccd1 _12929_/A sky130_fd_sc_hd__a21oi_1
XFILLER_80_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16695_ _19541_/Q _19540_/Q _19539_/Q _16695_/D vssd1 vssd1 vccd1 vccd1 _16704_/D
+ sky130_fd_sc_hd__and4_1
X_19483_ _19491_/CLK _19483_/D vssd1 vssd1 vccd1 vccd1 _19483_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18434_ _19284_/CLK _18434_/D vssd1 vssd1 vccd1 vccd1 _18434_/Q sky130_fd_sc_hd__dfxtp_1
X_15646_ _15646_/A vssd1 vssd1 vccd1 vccd1 _19172_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12858_ _15998_/A _16011_/A _12861_/A vssd1 vssd1 vccd1 vccd1 _12858_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11809_ _11809_/A _11830_/B vssd1 vssd1 vccd1 vccd1 _11809_/Y sky130_fd_sc_hd__xnor2_1
X_18365_ _19248_/CLK _18365_/D vssd1 vssd1 vccd1 vccd1 _18365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15577_ _15603_/A vssd1 vssd1 vccd1 vccd1 _15596_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_15_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12789_ _19520_/Q _12782_/X _12635_/X _19488_/Q _12788_/X vssd1 vssd1 vccd1 vccd1
+ _12789_/X sky130_fd_sc_hd__a221o_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17316_ _17864_/S _12487_/B _17294_/S vssd1 vssd1 vccd1 vccd1 _17316_/X sky130_fd_sc_hd__a21o_1
X_14528_ _14528_/A vssd1 vssd1 vccd1 vccd1 _14528_/X sky130_fd_sc_hd__clkbuf_1
X_18296_ _19311_/CLK _18296_/D vssd1 vssd1 vccd1 vccd1 _18296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17247_ _17247_/A vssd1 vssd1 vccd1 vccd1 _17587_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14459_ _13857_/X _18715_/Q _14467_/S vssd1 vssd1 vccd1 vccd1 _14460_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16740__A1 _16752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17178_ _17203_/A vssd1 vssd1 vccd1 vccd1 _17240_/S sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09222__A2 _13619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12804__B _16000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16129_ _16114_/X _12715_/X _16128_/Y vssd1 vssd1 vccd1 vccd1 _16129_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12109__A2 _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09605__S0 _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11868__B2 _19864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14511__S _14511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19819_ _19845_/CLK _19819_/D vssd1 vssd1 vccd1 vccd1 _19819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09908__S1 _09905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16008__B1 _13423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09503_ _11100_/A vssd1 vssd1 vccd1 vccd1 _10965_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13490__A0 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15342__S _15350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _09434_/A vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__clkbuf_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12045__A1 _16114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ _09341_/A _11522_/A _09468_/A vssd1 vssd1 vccd1 vccd1 _09366_/A sky130_fd_sc_hd__o21ba_4
XFILLER_21_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11171__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09296_ _19627_/Q _19622_/Q _19623_/Q _19628_/Q vssd1 vssd1 vccd1 vccd1 _09296_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10151__S0 _09930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13545__A1 _13544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09576__A _09576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10140_ _09715_/A _10139_/X _09941_/A vssd1 vssd1 vccd1 vccd1 _10140_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_165_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput170 _16255_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[6] sky130_fd_sc_hd__buf_2
XFILLER_88_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10071_ _10289_/A _10071_/B vssd1 vssd1 vccd1 vccd1 _10071_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12730__A _18112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13830_ _13830_/A vssd1 vssd1 vccd1 vccd1 _18477_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ _13761_/A vssd1 vssd1 vccd1 vccd1 _18447_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12284__A1 _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10973_ _11085_/A _10972_/X _09481_/A vssd1 vssd1 vccd1 vccd1 _10973_/X sky130_fd_sc_hd__o21a_1
XFILLER_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15500_ _15629_/A _18258_/Q vssd1 vssd1 vccd1 vccd1 _15500_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15252__S _15256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12712_ _18275_/Q _12712_/B vssd1 vssd1 vccd1 vccd1 _12712_/X sky130_fd_sc_hd__or2_1
X_16480_ _19477_/Q _16476_/B _16479_/Y vssd1 vssd1 vccd1 vccd1 _19477_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13692_ _18091_/A _15173_/A _13947_/B vssd1 vssd1 vccd1 vccd1 _13749_/A sky130_fd_sc_hd__or3_4
XFILLER_70_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15431_ _19122_/Q _15057_/X _15433_/S vssd1 vssd1 vccd1 vccd1 _15432_/A sky130_fd_sc_hd__mux2_1
XFILLER_102_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12643_ _19675_/Q _12601_/A _12565_/A _19642_/Q _12642_/X vssd1 vssd1 vccd1 vccd1
+ _12643_/X sky130_fd_sc_hd__a221o_1
XFILLER_169_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12587__A2 _12584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18150_ _18150_/A _18150_/B vssd1 vssd1 vccd1 vccd1 _18151_/A sky130_fd_sc_hd__or2_1
X_15362_ _15362_/A vssd1 vssd1 vccd1 vccd1 _19091_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _15599_/A _18268_/Q vssd1 vssd1 vccd1 vccd1 _12574_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11512__C _11918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10142__S0 _09930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17101_ _18146_/B vssd1 vssd1 vccd1 vccd1 _18091_/B sky130_fd_sc_hd__buf_2
X_14313_ _13857_/X _18651_/Q _14321_/S vssd1 vssd1 vccd1 vccd1 _14314_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18081_ _18081_/A _18087_/B vssd1 vssd1 vccd1 vccd1 _18081_/X sky130_fd_sc_hd__or2_1
XFILLER_7_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11525_ _11525_/A _17114_/C vssd1 vssd1 vccd1 vccd1 _11574_/B sky130_fd_sc_hd__nand2_1
XFILLER_156_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15293_ _15293_/A vssd1 vssd1 vccd1 vccd1 _19060_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17032_ _17032_/A vssd1 vssd1 vccd1 vccd1 _19664_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13536__A1 _13535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14244_ _14255_/A vssd1 vssd1 vccd1 vccd1 _14253_/S sky130_fd_sc_hd__buf_2
X_11456_ _11456_/A _12457_/B vssd1 vssd1 vccd1 vccd1 _11456_/X sky130_fd_sc_hd__and2_1
XANTENNA__09204__A2 _19811_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10407_ _18466_/Q _19057_/Q _19219_/Q _18434_/Q _09681_/A _10312_/A vssd1 vssd1 vccd1
+ vccd1 _10407_/X sky130_fd_sc_hd__mux4_2
X_14175_ _14175_/A vssd1 vssd1 vccd1 vccd1 _18598_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11387_ _11387_/A vssd1 vssd1 vccd1 vccd1 _11388_/S sky130_fd_sc_hd__buf_2
XFILLER_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13126_ _13126_/A vssd1 vssd1 vccd1 vccd1 _18299_/D sky130_fd_sc_hd__clkbuf_1
X_10338_ _10331_/Y _10333_/Y _10335_/Y _10337_/Y _09831_/A vssd1 vssd1 vccd1 vccd1
+ _10338_/X sky130_fd_sc_hd__o221a_4
XFILLER_124_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18983_ _19109_/CLK _18983_/D vssd1 vssd1 vccd1 vccd1 _18983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10770__A1 _09597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15427__S _15433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _19151_/Q _13007_/X _12566_/X _19341_/Q _13056_/X vssd1 vssd1 vccd1 vccd1
+ _13057_/X sky130_fd_sc_hd__a221o_2
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _17934_/A vssd1 vssd1 vccd1 vccd1 _19742_/D sky130_fd_sc_hd__clkbuf_1
X_10269_ _10269_/A vssd1 vssd1 vccd1 vccd1 _10269_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12008_ _12008_/A _12008_/B vssd1 vssd1 vccd1 vccd1 _12009_/B sky130_fd_sc_hd__xor2_4
XFILLER_120_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17865_ _17867_/A _17867_/B vssd1 vssd1 vccd1 vccd1 _17865_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19604_ _19607_/CLK _19604_/D vssd1 vssd1 vccd1 vccd1 _19604_/Q sky130_fd_sc_hd__dfxtp_1
X_16816_ _19578_/Q _16816_/B _19576_/Q _16816_/D vssd1 vssd1 vccd1 vccd1 _16821_/C
+ sky130_fd_sc_hd__and4_1
X_17796_ _12149_/Y _17786_/X _17794_/X _17795_/X vssd1 vssd1 vccd1 vccd1 _17796_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15461__A1 _13404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19535_ _19541_/CLK _19535_/D vssd1 vssd1 vccd1 vccd1 _19535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16747_ _16752_/B _16742_/B _19559_/Q vssd1 vssd1 vccd1 vccd1 _16751_/B sky130_fd_sc_hd__a21oi_1
X_13959_ _14531_/A vssd1 vssd1 vccd1 vccd1 _13959_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16678_ _16681_/C _16681_/D _19535_/Q vssd1 vssd1 vccd1 vccd1 _16680_/B sky130_fd_sc_hd__a21oi_1
X_19466_ _19603_/CLK _19466_/D vssd1 vssd1 vccd1 vccd1 _19466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11703__B _11703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18417_ _19202_/CLK _18417_/D vssd1 vssd1 vccd1 vccd1 _18417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15629_ _15629_/A hold7/A vssd1 vssd1 vccd1 vccd1 _15629_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17878__A _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19397_ _19699_/CLK _19397_/D vssd1 vssd1 vccd1 vccd1 _19397_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_166_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12578__A2 _12556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11235__C1 _10929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09150_ _09338_/C _09175_/C vssd1 vssd1 vccd1 vccd1 _09158_/B sky130_fd_sc_hd__nor2_1
X_18348_ _19325_/CLK _18348_/D vssd1 vssd1 vccd1 vccd1 _18348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18279_ _18282_/CLK _18279_/D vssd1 vssd1 vccd1 vccd1 _18279_/Q sky130_fd_sc_hd__dfxtp_1
X_09081_ _19841_/Q _19839_/Q _19840_/Q vssd1 vssd1 vccd1 vccd1 _09180_/C sky130_fd_sc_hd__or3b_1
XFILLER_174_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__clkbuf_2
Xinput61 io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
XFILLER_128_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10335__A _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09983_ _09688_/A _09981_/X _10559_/A vssd1 vssd1 vccd1 vccd1 _09983_/X sky130_fd_sc_hd__a21o_1
XFILLER_103_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15580__B _15580_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ _09705_/A vssd1 vssd1 vccd1 vccd1 _09590_/A sky130_fd_sc_hd__buf_2
XFILLER_53_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17788__A _17790_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16952__A1 _15481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ _19864_/Q vssd1 vssd1 vccd1 vccd1 _17125_/A sky130_fd_sc_hd__buf_4
XANTENNA__10124__S0 _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09279_ _09274_/C _09270_/A _12584_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _09280_/D
+ sky130_fd_sc_hd__a31o_1
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ _19311_/Q _18723_/Q _18760_/Q _18334_/Q _10660_/X _09707_/A vssd1 vssd1 vccd1
+ vccd1 _11310_/X sky130_fd_sc_hd__mux4_1
XFILLER_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12290_ _12312_/A _12268_/B _12265_/A _17845_/B vssd1 vssd1 vccd1 vccd1 _12291_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_147_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12444__B _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09198__A1 _09194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11241_ _18481_/Q _18976_/Q _11241_/S vssd1 vssd1 vccd1 vccd1 _11242_/B sky130_fd_sc_hd__mux2_1
XFILLER_10_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12741__A2 _12739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ _18484_/Q _18979_/Q _11172_/S vssd1 vssd1 vccd1 vccd1 _11172_/X sky130_fd_sc_hd__mux2_1
XFILLER_164_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17028__A _17028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ _10116_/X _10118_/Y _10120_/Y _10122_/Y _09813_/X vssd1 vssd1 vccd1 vccd1
+ _10123_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15980_ _15980_/A vssd1 vssd1 vccd1 vccd1 _19321_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12460__A _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input33_A io_dbus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _10054_/A vssd1 vssd1 vccd1 vccd1 _10054_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14931_ _14931_/A vssd1 vssd1 vccd1 vccd1 _18911_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14862_ _14930_/S vssd1 vssd1 vccd1 vccd1 _14871_/S sky130_fd_sc_hd__clkbuf_4
X_17650_ _11877_/A _17737_/A _17645_/Y _17649_/X _11539_/S vssd1 vssd1 vccd1 vccd1
+ _17650_/X sky130_fd_sc_hd__o221a_2
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16601_ _19514_/Q _16604_/C _16590_/X vssd1 vssd1 vccd1 vccd1 _16601_/Y sky130_fd_sc_hd__a21oi_1
X_13813_ _13813_/A vssd1 vssd1 vccd1 vccd1 _18469_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17581_ _17864_/S vssd1 vssd1 vccd1 vccd1 _17832_/S sky130_fd_sc_hd__buf_2
XFILLER_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14793_ _18849_/Q _13953_/X _14799_/S vssd1 vssd1 vccd1 vccd1 _14794_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16532_ _16714_/A vssd1 vssd1 vccd1 vccd1 _16570_/A sky130_fd_sc_hd__clkbuf_2
X_19320_ _19320_/CLK _19320_/D vssd1 vssd1 vccd1 vccd1 _19320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ _13744_/A vssd1 vssd1 vccd1 vccd1 _18439_/D sky130_fd_sc_hd__clkbuf_1
X_10956_ _11048_/A _10956_/B vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__or2_1
XFILLER_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19251_ _19315_/CLK _19251_/D vssd1 vssd1 vccd1 vccd1 _19251_/Q sky130_fd_sc_hd__dfxtp_1
X_16463_ _19471_/Q _16460_/B _16462_/Y vssd1 vssd1 vccd1 vccd1 _19471_/D sky130_fd_sc_hd__o21a_1
X_13675_ _13251_/X _18409_/Q _13675_/S vssd1 vssd1 vccd1 vccd1 _13676_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10887_ _11184_/A _10887_/B vssd1 vssd1 vccd1 vccd1 _10887_/X sky130_fd_sc_hd__or2_1
XFILLER_31_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18202_ _18231_/A _18202_/B vssd1 vssd1 vccd1 vccd1 _18203_/A sky130_fd_sc_hd__and2_1
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _19114_/Q _15031_/X _15422_/S vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__mux2_1
X_12626_ _18099_/A vssd1 vssd1 vccd1 vccd1 _18134_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19182_ _19184_/CLK _19182_/D vssd1 vssd1 vccd1 vccd1 _19182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16394_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16442_/A sky130_fd_sc_hd__buf_2
XFILLER_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18133_ _19828_/Q _18120_/X _18132_/X _18123_/X vssd1 vssd1 vccd1 vccd1 _19828_/D
+ sky130_fd_sc_hd__o211a_1
X_15345_ _15345_/A vssd1 vssd1 vccd1 vccd1 _19083_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16752__D _16752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12557_ _13397_/A vssd1 vssd1 vccd1 vccd1 _12557_/X sky130_fd_sc_hd__buf_2
XANTENNA__10854__S _10854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14326__S _14332_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__S1 _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18064_ _19801_/Q _19422_/Q _18066_/S vssd1 vssd1 vccd1 vccd1 _18065_/A sky130_fd_sc_hd__mux2_1
X_11508_ _11508_/A _11943_/A vssd1 vssd1 vccd1 vccd1 _12322_/B sky130_fd_sc_hd__and2_2
XFILLER_157_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15276_ _14563_/X _19053_/Q _15278_/S vssd1 vssd1 vccd1 vccd1 _15277_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12488_ _17317_/A _12488_/B vssd1 vssd1 vccd1 vccd1 _12488_/Y sky130_fd_sc_hd__nor2_4
X_17015_ _15615_/X _17010_/X _17014_/X _17008_/X vssd1 vssd1 vccd1 vccd1 _19658_/D
+ sky130_fd_sc_hd__o211a_1
X_14227_ _18621_/Q _13988_/X _14231_/S vssd1 vssd1 vccd1 vccd1 _14228_/A sky130_fd_sc_hd__mux2_1
XFILLER_160_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10418__S1 _09674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11439_ _11439_/A _11441_/A _11439_/C vssd1 vssd1 vccd1 vccd1 _11439_/Y sky130_fd_sc_hd__nand3_1
XFILLER_171_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14158_ _18591_/Q _13994_/X _14158_/S vssd1 vssd1 vccd1 vccd1 _14159_/A sky130_fd_sc_hd__mux2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13109_ _13107_/X _18298_/Q _13172_/S vssd1 vssd1 vccd1 vccd1 _13110_/A sky130_fd_sc_hd__mux2_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14061__S _14063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _19127_/CLK _18966_/D vssd1 vssd1 vccd1 vccd1 _18966_/Q sky130_fd_sc_hd__dfxtp_1
X_14089_ _14089_/A vssd1 vssd1 vccd1 vccd1 _18560_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_101_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12370__A _19420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17671__A2 _17652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17917_ _17917_/A _17917_/B vssd1 vssd1 vccd1 vccd1 _17917_/X sky130_fd_sc_hd__or2_1
X_18897_ _19376_/CLK _18897_/D vssd1 vssd1 vccd1 vccd1 _18897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09361__A1 _13132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17848_ _17597_/X _17618_/X _17847_/X _17542_/X vssd1 vssd1 vccd1 vccd1 _17848_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_39_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14297__A _18089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17779_ _17779_/A _17779_/B vssd1 vssd1 vccd1 vccd1 _17779_/X sky130_fd_sc_hd__or2_1
XFILLER_47_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19518_ _19550_/CLK _19518_/D vssd1 vssd1 vccd1 vccd1 _19518_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12799__A2 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19449_ _19550_/CLK _19449_/D vssd1 vssd1 vccd1 vccd1 _19449_/Q sky130_fd_sc_hd__dfxtp_1
X_09202_ _19813_/Q vssd1 vssd1 vccd1 vccd1 _14197_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_10_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10106__S0 _10093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18216__B _18216_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09133_ _09174_/A _09174_/B vssd1 vssd1 vccd1 vccd1 _09134_/C sky130_fd_sc_hd__or2b_1
XANTENNA__10764__S _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14236__S _14242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12545__A _13400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10431__B1 _09764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15856__A _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09854__A _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _09968_/A _09965_/X _09823_/A vssd1 vssd1 vccd1 vccd1 _09966_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_104_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17790__B _17790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09897_ _09905_/A vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__clkbuf_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _18457_/Q _19048_/Q _19210_/Q _18425_/Q _09598_/A _10802_/X vssd1 vssd1 vccd1
+ vccd1 _10810_/X sky130_fd_sc_hd__mux4_2
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11790_/A _11790_/B vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__or2_2
XFILLER_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10741_ _10547_/A _10740_/X _09432_/A vssd1 vssd1 vccd1 vccd1 _10741_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_14_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17311__A _17317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _13460_/A vssd1 vssd1 vccd1 vccd1 _18330_/D sky130_fd_sc_hd__clkbuf_1
X_10672_ _18923_/Q _18689_/Q _19371_/Q _19019_/Q _10729_/S _10655_/X vssd1 vssd1 vccd1
+ vccd1 _10672_/X sky130_fd_sc_hd__mux4_1
X_12411_ _12175_/A _12409_/Y _12434_/B _11653_/X vssd1 vssd1 vccd1 vccd1 _12411_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ _13391_/A _13391_/B _13391_/C _13391_/D vssd1 vssd1 vccd1 vccd1 _13392_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15130_ _18988_/Q _15038_/X _15134_/S vssd1 vssd1 vccd1 vccd1 _15131_/A sky130_fd_sc_hd__mux2_1
XFILLER_166_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12342_ _19355_/Q _11733_/X _11734_/X _12341_/X _11691_/X vssd1 vssd1 vccd1 vccd1
+ _12342_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10973__A1 _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15061_ _18963_/Q _15060_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15062_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12273_ _12435_/A _12269_/Y _12272_/X vssd1 vssd1 vccd1 vccd1 _12273_/X sky130_fd_sc_hd__a21bo_1
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_3_0_clock_A clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ _14012_/A vssd1 vssd1 vccd1 vccd1 _18532_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09764__A _09764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _10920_/A _11223_/X _10914_/A vssd1 vssd1 vccd1 vccd1 _11224_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15485__B _15485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18820_ _19302_/CLK _18820_/D vssd1 vssd1 vccd1 vccd1 _18820_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11155_ _11160_/A _11155_/B vssd1 vssd1 vccd1 vccd1 _11155_/Y sky130_fd_sc_hd__nor2_1
XFILLER_150_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10703__A _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10106_ _18472_/Q _19063_/Q _19225_/Q _18440_/Q _10093_/S _09715_/A vssd1 vssd1 vccd1
+ vccd1 _10106_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_122_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18751_ _19302_/CLK _18751_/D vssd1 vssd1 vccd1 vccd1 _18751_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15963_ _15963_/A vssd1 vssd1 vccd1 vccd1 _19313_/D sky130_fd_sc_hd__clkbuf_1
X_11086_ _19302_/Q _18714_/Q _18751_/Q _18325_/Q _10969_/X _11266_/A vssd1 vssd1 vccd1
+ vccd1 _11086_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17702_ _17700_/Y _17701_/X _17739_/S vssd1 vssd1 vccd1 vccd1 _17703_/B sky130_fd_sc_hd__mux2_1
XFILLER_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14914_ _14914_/A vssd1 vssd1 vccd1 vccd1 _18903_/D sky130_fd_sc_hd__clkbuf_1
X_10037_ _18412_/Q _18673_/Q _18572_/Q _18907_/Q _10764_/S _09380_/A vssd1 vssd1 vccd1
+ vccd1 _10038_/B sky130_fd_sc_hd__mux4_1
X_15894_ _19283_/Q _14576_/A _15898_/S vssd1 vssd1 vccd1 vccd1 _15895_/A sky130_fd_sc_hd__mux2_1
X_18682_ _19012_/CLK _18682_/D vssd1 vssd1 vccd1 vccd1 _18682_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11150__A1 _10904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10584__S0 _10576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17633_ _17633_/A vssd1 vssd1 vccd1 vccd1 _17633_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14845_ _14845_/A vssd1 vssd1 vccd1 vccd1 _14854_/S sky130_fd_sc_hd__buf_4
XFILLER_84_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15006__A _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17564_ _17468_/A _17560_/Y _17563_/Y vssd1 vssd1 vccd1 vccd1 _17564_/Y sky130_fd_sc_hd__a21oi_1
X_14776_ _14776_/A vssd1 vssd1 vccd1 vccd1 _18842_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10336__S0 _10286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11988_ _11988_/A vssd1 vssd1 vccd1 vccd1 _11988_/Y sky130_fd_sc_hd__inv_2
X_19303_ _19305_/CLK _19303_/D vssd1 vssd1 vccd1 vccd1 _19303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16515_ _19611_/Q _19610_/Q _19612_/Q _16891_/A vssd1 vssd1 vccd1 vccd1 _16899_/A
+ sky130_fd_sc_hd__and4_1
X_13727_ _13749_/A vssd1 vssd1 vccd1 vccd1 _13736_/S sky130_fd_sc_hd__buf_6
X_10939_ _11241_/S vssd1 vssd1 vccd1 vccd1 _10940_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10110__C1 _09754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17495_ _17466_/X _17489_/X _17493_/Y _17494_/X vssd1 vssd1 vccd1 vccd1 _17495_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15440__S _15444_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19234_ _19298_/CLK _19234_/D vssd1 vssd1 vccd1 vccd1 _19234_/Q sky130_fd_sc_hd__dfxtp_1
X_16446_ _16546_/A vssd1 vssd1 vccd1 vccd1 _16446_/X sky130_fd_sc_hd__clkbuf_2
X_13658_ _13124_/X _18401_/Q _13664_/S vssd1 vssd1 vccd1 vccd1 _13659_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ _19141_/Q _12526_/X _12565_/X _19634_/Q _12608_/X vssd1 vssd1 vccd1 vccd1
+ _12609_/X sky130_fd_sc_hd__a221o_1
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16377_ _19441_/Q _16379_/C _16376_/Y vssd1 vssd1 vccd1 vccd1 _19441_/D sky130_fd_sc_hd__o21a_1
X_19165_ _19598_/CLK _19165_/D vssd1 vssd1 vccd1 vccd1 _19165_/Q sky130_fd_sc_hd__dfxtp_1
X_13589_ _15073_/A vssd1 vssd1 vccd1 vccd1 _13589_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18116_ _18116_/A _18116_/B vssd1 vssd1 vccd1 vccd1 _18116_/X sky130_fd_sc_hd__or2_1
X_15328_ _19076_/Q _15012_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15329_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19096_ _19096_/CLK _19096_/D vssd1 vssd1 vccd1 vccd1 _19096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15259_ _14537_/X _19045_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15260_/A sky130_fd_sc_hd__mux2_1
X_18047_ _18047_/A vssd1 vssd1 vccd1 vccd1 _19793_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18052__A _18188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12705__A2 _12703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__A _09674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10177__C1 _09813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _09820_/A vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__buf_2
XFILLER_87_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16852__B1 _16812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09751_ _11368_/A _09748_/X _09750_/X _09740_/X vssd1 vssd1 vccd1 vccd1 _09751_/X
+ sky130_fd_sc_hd__o211a_1
X_18949_ _19109_/CLK _18949_/D vssd1 vssd1 vccd1 vccd1 _18949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09682_ _09682_/A vssd1 vssd1 vccd1 vccd1 _10186_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10101__C1 _09859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15350__S _15350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17131__A _18142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09849__A _10546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_164_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09116_ _09116_/A vssd1 vssd1 vccd1 vccd1 _17122_/A sky130_fd_sc_hd__buf_4
XFILLER_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16135__A2 _15600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09584__A _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10707__A1 _11321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11619__A _11619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09949_ _09667_/A _09939_/X _09948_/X _09758_/A _19731_/Q vssd1 vssd1 vccd1 vccd1
+ _10087_/A sky130_fd_sc_hd__a32o_4
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12960_ _19560_/Q vssd1 vssd1 vccd1 vccd1 _16760_/B sky130_fd_sc_hd__buf_2
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09420__S1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11911_ _11794_/A _11909_/X _11910_/Y vssd1 vssd1 vccd1 vccd1 _11911_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_85_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _19743_/Q _19744_/Q _12891_/C vssd1 vssd1 vccd1 vccd1 _12928_/C sky130_fd_sc_hd__and3_1
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16071__A1 _19342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ _14630_/A vssd1 vssd1 vccd1 vccd1 _18780_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11354__A _11354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11842_/A _11842_/B _11842_/C _11842_/D vssd1 vssd1 vccd1 vccd1 _11950_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_33_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14560_/X _18759_/Q _14567_/S vssd1 vssd1 vccd1 vccd1 _14562_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12632__A1 _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ _15474_/A vssd1 vssd1 vccd1 vccd1 _11773_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16300_ _12321_/A _16278_/X _12324_/X _12327_/Y _16280_/X vssd1 vssd1 vccd1 vccd1
+ _19418_/D sky130_fd_sc_hd__o221a_1
X_13512_ _13619_/C vssd1 vssd1 vccd1 vccd1 _18091_/A sky130_fd_sc_hd__buf_4
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17280_ _17572_/S vssd1 vssd1 vccd1 vccd1 _17613_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10724_ _09563_/A _10717_/Y _10719_/Y _10721_/Y _10723_/Y vssd1 vssd1 vccd1 vccd1
+ _10724_/X sky130_fd_sc_hd__o32a_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _13905_/X _18730_/Q _14500_/S vssd1 vssd1 vccd1 vccd1 _14493_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16231_ _13602_/X _19387_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16232_/A sky130_fd_sc_hd__mux2_1
X_13443_ _13443_/A vssd1 vssd1 vccd1 vccd1 _18322_/D sky130_fd_sc_hd__clkbuf_1
X_10655_ _10655_/A vssd1 vssd1 vccd1 vccd1 _10655_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11199__A1 _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16162_ _15631_/X _16161_/Y _16162_/S vssd1 vssd1 vccd1 vccd1 _16162_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13374_ _18320_/Q _12603_/X _12958_/A _19359_/Q vssd1 vssd1 vccd1 vccd1 _13374_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_155_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10586_ _10586_/A vssd1 vssd1 vccd1 vccd1 _10586_/X sky130_fd_sc_hd__buf_2
XFILLER_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15113_ _15113_/A vssd1 vssd1 vccd1 vccd1 _18980_/D sky130_fd_sc_hd__clkbuf_1
X_12325_ _19657_/Q _12343_/C vssd1 vssd1 vccd1 vccd1 _12325_/Y sky130_fd_sc_hd__nor2_1
XFILLER_115_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16093_ _16098_/B _16092_/Y _13418_/A vssd1 vssd1 vccd1 vccd1 _16093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_127_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_170_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09494__A _11219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15044_ _15044_/A vssd1 vssd1 vccd1 vccd1 _15044_/X sky130_fd_sc_hd__clkbuf_2
X_12256_ _19654_/Q _19653_/Q _12256_/C vssd1 vssd1 vccd1 vccd1 _12298_/C sky130_fd_sc_hd__and3_1
XFILLER_107_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11207_ _19299_/Q _18711_/Q _18748_/Q _18322_/Q _11243_/S _11177_/A vssd1 vssd1 vccd1
+ vccd1 _11208_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09564__A1 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19852_ _19854_/CLK _19852_/D vssd1 vssd1 vccd1 vccd1 _19852_/Q sky130_fd_sc_hd__dfxtp_1
X_12187_ _12181_/X _12186_/Y _19412_/Q _12078_/A vssd1 vssd1 vccd1 vccd1 _16288_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_150_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18803_ _19379_/CLK _18803_/D vssd1 vssd1 vccd1 vccd1 _18803_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16834__B1 _16812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ _11138_/A _11138_/B vssd1 vssd1 vccd1 vccd1 _11138_/X sky130_fd_sc_hd__or2_1
X_19783_ _19786_/CLK _19783_/D vssd1 vssd1 vccd1 vccd1 _19783_/Q sky130_fd_sc_hd__dfxtp_2
X_16995_ _18097_/A vssd1 vssd1 vccd1 vccd1 _16995_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18734_ _19384_/CLK _18734_/D vssd1 vssd1 vccd1 vccd1 _18734_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11069_ _11059_/X _11062_/X _11064_/X _11068_/X _09465_/A vssd1 vssd1 vccd1 vccd1
+ _11069_/X sky130_fd_sc_hd__a221o_2
X_15946_ _13541_/X _19306_/Q _15948_/S vssd1 vssd1 vccd1 vccd1 _15947_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18665_ _19027_/CLK _18665_/D vssd1 vssd1 vccd1 vccd1 _18665_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15877_ _15877_/A vssd1 vssd1 vccd1 vccd1 _19275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17616_ _17615_/A _17508_/A _17615_/Y _17716_/S vssd1 vssd1 vccd1 vccd1 _17616_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14828_ _18865_/Q _14004_/X _14832_/S vssd1 vssd1 vccd1 vccd1 _14829_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18596_ _19091_/CLK _18596_/D vssd1 vssd1 vccd1 vccd1 _18596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17547_ _19711_/Q _17430_/X _17545_/X _17546_/X vssd1 vssd1 vccd1 vccd1 _19711_/D
+ sky130_fd_sc_hd__o22a_1
X_14759_ _14582_/X _18835_/Q _14759_/S vssd1 vssd1 vccd1 vccd1 _14760_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09669__A _09669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17478_ _17478_/A vssd1 vssd1 vccd1 vccd1 _17478_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19217_ _19249_/CLK _19217_/D vssd1 vssd1 vccd1 vccd1 _19217_/Q sky130_fd_sc_hd__dfxtp_1
X_16429_ _16431_/B _16431_/C _16402_/X vssd1 vssd1 vccd1 vccd1 _16429_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17886__A _17907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19148_ _19693_/CLK _19148_/D vssd1 vssd1 vccd1 vccd1 _19148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17314__A1 _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19079_ _19329_/CLK _19079_/D vssd1 vssd1 vccd1 vccd1 _19079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13887__A0 _13886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12542__B _12542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09803_ _09803_/A vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17126__A _18122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09734_ _18605_/Q _18876_/Q _19100_/Q _18844_/Q _09704_/X _09733_/X vssd1 vssd1 vccd1
+ vccd1 _09734_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16030__A _16086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__A1 _11116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ _09665_/A vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__buf_2
XFILLER_83_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16053__A1 _19339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__A _11174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ _09596_/A vssd1 vssd1 vccd1 vccd1 _10547_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16176__S _16180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12090__A2 _12089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10720__S0 _10631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11621__B _18125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10440_ _18402_/Q _18663_/Q _18562_/Q _18897_/Q _10341_/S _09886_/A vssd1 vssd1 vccd1
+ vccd1 _10440_/X sky130_fd_sc_hd__mux4_1
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10371_ _18595_/Q _18866_/Q _19090_/Q _18834_/Q _09700_/A _10229_/X vssd1 vssd1 vccd1
+ vccd1 _10371_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14424__S _14428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12110_ _12110_/A _17768_/B vssd1 vssd1 vccd1 vccd1 _12140_/D sky130_fd_sc_hd__nand2_1
X_13090_ _14566_/A vssd1 vssd1 vccd1 vccd1 _13090_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_152_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ _12040_/Y _12035_/Y _12179_/B vssd1 vssd1 vccd1 vccd1 _12041_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11349__A _11445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15800_ _13538_/X _19241_/Q _15804_/S vssd1 vssd1 vccd1 vccd1 _15801_/A sky130_fd_sc_hd__mux2_1
X_16780_ _19565_/Q _19564_/Q _16780_/C _16780_/D vssd1 vssd1 vccd1 vccd1 _16788_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13992_ _18526_/Q _13991_/X _13995_/S vssd1 vssd1 vccd1 vccd1 _13993_/A sky130_fd_sc_hd__mux2_1
XFILLER_120_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15731_ _15731_/A vssd1 vssd1 vccd1 vccd1 _19210_/D sky130_fd_sc_hd__clkbuf_1
X_12943_ input30/X _12781_/A _12942_/X _12831_/X vssd1 vssd1 vccd1 vccd1 _15022_/A
+ sky130_fd_sc_hd__a22o_2
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14055__A0 _13837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18450_ _19235_/CLK _18450_/D vssd1 vssd1 vccd1 vccd1 _18450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12874_ _18315_/Q _12603_/X _12640_/X _19332_/Q vssd1 vssd1 vccd1 vccd1 _12874_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15662_ _15708_/S vssd1 vssd1 vccd1 vccd1 _15671_/S sky130_fd_sc_hd__buf_2
XFILLER_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17483_/A vssd1 vssd1 vccd1 vccd1 _17402_/A sky130_fd_sc_hd__clkbuf_2
X_14613_ _14613_/A vssd1 vssd1 vccd1 vccd1 _18775_/D sky130_fd_sc_hd__clkbuf_1
X_11825_ _11826_/A _12098_/C _19399_/Q vssd1 vssd1 vccd1 vccd1 _11827_/A sky130_fd_sc_hd__a21oi_1
X_15593_ _15592_/X _19161_/Q _15596_/S vssd1 vssd1 vccd1 vccd1 _15594_/A sky130_fd_sc_hd__mux2_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output102_A _11877_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18381_ _19388_/CLK _18381_/D vssd1 vssd1 vccd1 vccd1 _18381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12908__A _13387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13503__S _13503_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14544_ _14544_/A vssd1 vssd1 vccd1 vccd1 _14544_/X sky130_fd_sc_hd__clkbuf_2
X_17332_ _17541_/A vssd1 vssd1 vccd1 vccd1 _17646_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _11670_/A _12448_/B _11813_/A _18132_/A vssd1 vssd1 vccd1 vccd1 _17563_/A
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10711__S0 _11318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _11321_/A _10706_/X _10719_/A vssd1 vssd1 vccd1 vccd1 _10707_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_81_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17263_ _17263_/A vssd1 vssd1 vccd1 vccd1 _17283_/S sky130_fd_sc_hd__clkbuf_2
X_14475_ _14475_/A vssd1 vssd1 vccd1 vccd1 _18722_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11687_ _19395_/Q _11736_/C vssd1 vssd1 vccd1 vccd1 _11687_/X sky130_fd_sc_hd__xor2_1
XFILLER_128_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19002_ _19098_/CLK _19002_/D vssd1 vssd1 vccd1 vccd1 _19002_/Q sky130_fd_sc_hd__dfxtp_1
X_16214_ _16214_/A vssd1 vssd1 vccd1 vccd1 _19379_/D sky130_fd_sc_hd__clkbuf_1
X_13426_ _15613_/A hold4/A vssd1 vssd1 vccd1 vccd1 _13426_/Y sky130_fd_sc_hd__nand2_1
X_10638_ _18397_/Q _18658_/Q _18557_/Q _18892_/Q _10576_/X _09651_/A vssd1 vssd1 vccd1
+ vccd1 _10638_/X sky130_fd_sc_hd__mux4_1
X_17194_ _17737_/A vssd1 vssd1 vccd1 vccd1 _17328_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_167_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_128_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16145_ _16114_/X _15615_/X _16144_/Y vssd1 vssd1 vccd1 vccd1 _16145_/X sky130_fd_sc_hd__a21o_1
X_13357_ _19454_/Q _12584_/Y _12586_/B _19518_/Q _13356_/X vssd1 vssd1 vccd1 vccd1
+ _13357_/X sky130_fd_sc_hd__a221o_1
XFILLER_127_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10569_ _10689_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__nor2_1
XFILLER_155_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19278_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_154_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12308_ _19797_/Q _10082_/A _12404_/S vssd1 vssd1 vccd1 vccd1 _12309_/A sky130_fd_sc_hd__mux2_4
XFILLER_143_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16076_ _15550_/X _16075_/Y _16082_/S vssd1 vssd1 vccd1 vccd1 _16076_/X sky130_fd_sc_hd__mux2_1
X_13288_ _16715_/C _13004_/X _13054_/X _19514_/Q _13287_/X vssd1 vssd1 vccd1 vccd1
+ _13288_/X sky130_fd_sc_hd__a221o_1
XFILLER_142_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15027_ _15027_/A vssd1 vssd1 vccd1 vccd1 _18952_/D sky130_fd_sc_hd__clkbuf_1
X_12239_ _12301_/A _12472_/B _12238_/Y vssd1 vssd1 vccd1 vccd1 _12240_/A sky130_fd_sc_hd__o21a_1
XFILLER_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13333__A2 _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__S0 _10633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16769__B _16772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19835_ _19838_/CLK _19835_/D vssd1 vssd1 vccd1 vccd1 _19835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15165__S _15167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19766_ _19799_/CLK _19766_/D vssd1 vssd1 vccd1 vccd1 _19766_/Q sky130_fd_sc_hd__dfxtp_1
X_16978_ _16978_/A _16984_/B vssd1 vssd1 vccd1 vccd1 _16978_/X sky130_fd_sc_hd__or2_1
XFILLER_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 io_dbus_rdata[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_65_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18717_ _19305_/CLK _18717_/D vssd1 vssd1 vccd1 vccd1 _18717_/Q sky130_fd_sc_hd__dfxtp_1
X_15929_ _13509_/X _19298_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15930_/A sky130_fd_sc_hd__mux2_1
X_19697_ _19845_/CLK _19697_/D vssd1 vssd1 vccd1 vccd1 _19697_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12844__A1 _13415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09450_ _09450_/A vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__buf_2
X_18648_ _19268_/CLK _18648_/D vssd1 vssd1 vccd1 vccd1 _18648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09381_ _10031_/A vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__clkbuf_4
X_18579_ _19074_/CLK _18579_/D vssd1 vssd1 vccd1 vccd1 _18579_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14509__S _14511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09399__A _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18224__B _18224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12780__B1 _18744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09528__A1 _10347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10073__A _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09717_ _09717_/A vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17223__A0 _17696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__S0 _11243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09648_ _10586_/A vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__buf_4
XFILLER_83_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17774__A1 _19724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15785__A0 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _09579_/A vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__clkbuf_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__A _12751_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_161_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ _17207_/A _12487_/B vssd1 vssd1 vccd1 vccd1 _11611_/A sky130_fd_sc_hd__and2_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12590_ _18269_/Q _12590_/B vssd1 vssd1 vccd1 vccd1 _12590_/X sky130_fd_sc_hd__or2_1
XFILLER_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12447__B _12447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15537__A0 _19720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09102__A _11528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11541_ _11541_/A vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__buf_2
XANTENNA__11351__B _12467_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14260_ _18636_/Q _14036_/X _14264_/S vssd1 vssd1 vccd1 vccd1 _14261_/A sky130_fd_sc_hd__mux2_1
X_11472_ _11453_/Y _11455_/X _11458_/X _11460_/Y _11471_/X vssd1 vssd1 vccd1 vccd1
+ _11472_/X sky130_fd_sc_hd__a2111o_1
XANTENNA__09216__B1 _19701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13211_ _13211_/A vssd1 vssd1 vccd1 vccd1 _18304_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10423_ _09666_/A _10411_/X _10422_/X _09757_/A _19724_/Q vssd1 vssd1 vccd1 vccd1
+ _11445_/A sky130_fd_sc_hd__a32o_4
XANTENNA__11023__B1 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14154__S _14158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14191_ _18606_/Q _14042_/X _14191_/S vssd1 vssd1 vccd1 vccd1 _14192_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12771__B1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13142_ _16091_/B _13152_/C vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__xor2_1
XANTENNA_input63_A io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10354_ _09762_/A _10338_/X _10352_/X _09835_/A _10353_/Y vssd1 vssd1 vccd1 vccd1
+ _12467_/B sky130_fd_sc_hd__o32a_4
XFILLER_151_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ input6/X _12974_/A _12977_/A vssd1 vssd1 vccd1 vccd1 _13088_/A sky130_fd_sc_hd__a21o_1
X_17950_ _17950_/A vssd1 vssd1 vccd1 vccd1 _19749_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10285_ _10429_/A vssd1 vssd1 vccd1 vccd1 _10390_/A sky130_fd_sc_hd__buf_2
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16901_ _19612_/Q _16898_/B _16900_/Y vssd1 vssd1 vccd1 vccd1 _19612_/D sky130_fd_sc_hd__o21a_1
X_12024_ _12020_/X _12462_/A _12023_/Y vssd1 vssd1 vccd1 vccd1 _12140_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__15493__B _15493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17881_ _17478_/X _17527_/X _17880_/X _17633_/X vssd1 vssd1 vccd1 vccd1 _17881_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19620_ _19834_/CLK _19620_/D vssd1 vssd1 vccd1 vccd1 _19620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16832_ _19588_/Q vssd1 vssd1 vccd1 vccd1 _16836_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19551_ _19564_/CLK _19551_/D vssd1 vssd1 vccd1 vccd1 _19551_/Q sky130_fd_sc_hd__dfxtp_2
X_16763_ _19562_/Q _16761_/B _16762_/Y vssd1 vssd1 vccd1 vccd1 _19562_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12826__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12826__B2 _12798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ _14547_/A vssd1 vssd1 vccd1 vccd1 _13975_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11185__S0 _10873_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18502_ _19286_/CLK _18502_/D vssd1 vssd1 vccd1 vccd1 _18502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15713__S _15721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15714_ _15714_/A vssd1 vssd1 vccd1 vccd1 _19202_/D sky130_fd_sc_hd__clkbuf_1
X_19482_ _19619_/CLK _19482_/D vssd1 vssd1 vccd1 vccd1 _19482_/Q sky130_fd_sc_hd__dfxtp_1
X_12926_ _12926_/A vssd1 vssd1 vccd1 vccd1 _18289_/D sky130_fd_sc_hd__clkbuf_1
X_16694_ _16697_/C _16697_/D _19541_/Q vssd1 vssd1 vccd1 vccd1 _16696_/B sky130_fd_sc_hd__a21oi_1
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10301__A2 _10284_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18433_ _19314_/CLK _18433_/D vssd1 vssd1 vccd1 vccd1 _18433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ _14528_/X _19172_/Q _15649_/S vssd1 vssd1 vccd1 vccd1 _15646_/A sky130_fd_sc_hd__mux2_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _19742_/Q vssd1 vssd1 vccd1 vccd1 _16011_/A sky130_fd_sc_hd__buf_2
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11542__A _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11808_ _11778_/C _11806_/Y _11807_/Y vssd1 vssd1 vccd1 vccd1 _11830_/B sky130_fd_sc_hd__a21oi_1
X_18364_ _19245_/CLK _18364_/D vssd1 vssd1 vccd1 vccd1 _18364_/Q sky130_fd_sc_hd__dfxtp_1
X_12788_ _19424_/Q _12636_/X _12787_/X vssd1 vssd1 vccd1 vccd1 _12788_/X sky130_fd_sc_hd__o21a_1
X_15576_ _19727_/Q _15574_/X _15595_/S vssd1 vssd1 vccd1 vccd1 _15576_/X sky130_fd_sc_hd__mux2_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10065__A1 _09485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15528__A0 _19718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17315_ _17485_/A vssd1 vssd1 vccd1 vccd1 _17864_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_147_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14527_ _14527_/A vssd1 vssd1 vccd1 vccd1 _18748_/D sky130_fd_sc_hd__clkbuf_1
X_11739_ _11737_/Y _11732_/X _14275_/B vssd1 vssd1 vccd1 vccd1 _11739_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10158__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18295_ _18894_/CLK _18295_/D vssd1 vssd1 vccd1 vccd1 _18295_/Q sky130_fd_sc_hd__dfxtp_1
X_17246_ _17605_/B _12289_/A _17274_/A vssd1 vssd1 vccd1 vccd1 _17246_/X sky130_fd_sc_hd__mux2_1
X_14458_ _14515_/S vssd1 vssd1 vccd1 vccd1 _14467_/S sky130_fd_sc_hd__buf_2
XFILLER_116_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13409_ _15494_/A _18252_/Q vssd1 vssd1 vccd1 vccd1 _13409_/Y sky130_fd_sc_hd__nand2_1
XFILLER_128_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14389_ _13861_/X _18684_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14390_/A sky130_fd_sc_hd__mux2_1
X_17177_ _17177_/A _17177_/B _17177_/C vssd1 vssd1 vccd1 vccd1 _17203_/A sky130_fd_sc_hd__nor3_4
XFILLER_116_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_152_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19300_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_155_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16128_ _16133_/B _16127_/Y _16109_/X vssd1 vssd1 vccd1 vccd1 _16128_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_115_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15684__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16059_ _12669_/X _16057_/Y _16082_/S vssd1 vssd1 vccd1 vccd1 _16059_/X sky130_fd_sc_hd__mux2_1
XFILLER_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11317__B2 _19720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__S1 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09682__A _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_167_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19201_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19818_ _19834_/CLK _19818_/D vssd1 vssd1 vccd1 vccd1 _19818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10540__A2 _10529_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12278__C1 _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19749_ _19779_/CLK _19749_/D vssd1 vssd1 vccd1 vccd1 _19749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ _11033_/A vssd1 vssd1 vccd1 vccd1 _11100_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09433_ _09608_/A vssd1 vssd1 vccd1 vccd1 _09434_/A sky130_fd_sc_hd__buf_4
XANTENNA__12548__A _12548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13143__S _13143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09341_/A _09193_/X _09198_/X _09204_/X _18742_/Q vssd1 vssd1 vccd1 vccd1
+ _09468_/A sky130_fd_sc_hd__o2111a_2
XFILLER_36_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_105_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19663_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09295_ _19629_/Q _19625_/Q _19663_/Q _19630_/Q vssd1 vssd1 vccd1 vccd1 _09295_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10151__S1 _10090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09857__A _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11598__S _12730_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14742__A1 _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12283__A _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12753__B1 _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_108_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput160 _12328_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[26] sky130_fd_sc_hd__buf_2
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput171 _16258_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[7] sky130_fd_sc_hd__buf_2
XFILLER_133_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10070_ _18476_/Q _19067_/Q _19229_/Q _18444_/Q _09500_/A _09543_/A vssd1 vssd1 vccd1
+ vccd1 _10071_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10516__C1 _09753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13842__A _13941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13760_ _13367_/X _18447_/Q _13762_/S vssd1 vssd1 vccd1 vccd1 _13761_/A sky130_fd_sc_hd__mux2_1
X_10972_ _18391_/Q _18652_/Q _18551_/Q _18886_/Q _10969_/X _11266_/A vssd1 vssd1 vccd1
+ vccd1 _10972_/X sky130_fd_sc_hd__mux4_1
X_12711_ _19612_/Q _12697_/X _12503_/A _19480_/Q _12710_/X vssd1 vssd1 vccd1 vccd1
+ _12712_/B sky130_fd_sc_hd__a221o_2
XFILLER_44_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13691_ _13691_/A vssd1 vssd1 vccd1 vccd1 _18416_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11362__A _11416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12642_ _19149_/Q _12895_/A _12640_/X _19339_/Q _12641_/X vssd1 vssd1 vccd1 vccd1
+ _12642_/X sky130_fd_sc_hd__a221o_1
X_15430_ _15430_/A vssd1 vssd1 vccd1 vccd1 _19121_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12177__B _19411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15361_ _19091_/Q _15060_/X _15361_/S vssd1 vssd1 vccd1 vccd1 _15362_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12573_ _15613_/A vssd1 vssd1 vccd1 vccd1 _15599_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_169_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17100_ _18071_/S vssd1 vssd1 vccd1 vccd1 _18146_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__10142__S1 _09871_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12992__A0 _19716_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14312_ _14369_/S vssd1 vssd1 vccd1 vccd1 _14321_/S sky130_fd_sc_hd__buf_2
XANTENNA__16183__A0 _13531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ _11647_/B _11521_/X _11523_/X vssd1 vssd1 vccd1 vccd1 _17110_/A sky130_fd_sc_hd__o21ai_2
X_15292_ _14585_/X _19060_/Q _15300_/S vssd1 vssd1 vccd1 vccd1 _15293_/A sky130_fd_sc_hd__mux2_1
X_18080_ _09172_/C _12739_/X _18079_/X vssd1 vssd1 vccd1 vccd1 _19807_/D sky130_fd_sc_hd__o21a_1
XFILLER_168_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17031_ _19664_/Q _13404_/X _17039_/S vssd1 vssd1 vccd1 vccd1 _17032_/A sky130_fd_sc_hd__mux2_1
X_14243_ _14243_/A vssd1 vssd1 vccd1 vccd1 _18628_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11455_ _11453_/B _11453_/C _11453_/A vssd1 vssd1 vccd1 vccd1 _11455_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10406_ _10406_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10406_/X sky130_fd_sc_hd__or2_1
XFILLER_171_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14174_ _18598_/Q _14017_/X _14180_/S vssd1 vssd1 vccd1 vccd1 _14175_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ _11386_/A vssd1 vssd1 vccd1 vccd1 _11386_/Y sky130_fd_sc_hd__inv_2
XFILLER_140_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13125_ _13124_/X _18299_/Q _13172_/S vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15708__S _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ _10390_/A _10336_/X _09765_/A vssd1 vssd1 vccd1 vccd1 _10337_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_84_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19693_/CLK sky130_fd_sc_hd__clkbuf_16
X_18982_ _19329_/CLK _18982_/D vssd1 vssd1 vccd1 vccd1 _18982_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14612__S _14615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _19677_/Q _13008_/X _13009_/X _19644_/Q vssd1 vssd1 vccd1 vccd1 _13056_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _16011_/A _19774_/Q _17935_/S vssd1 vssd1 vccd1 vccd1 _17934_/A sky130_fd_sc_hd__mux2_1
X_10268_ _18501_/Q _18996_/Q _10435_/S vssd1 vssd1 vccd1 vccd1 _10269_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10507__C1 _09669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12007_ _11959_/A _11959_/B _11987_/A _12006_/Y vssd1 vssd1 vccd1 vccd1 _12008_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_79_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15009__A _15009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11537__A _18744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17864_ _17867_/A _17867_/B _17864_/S vssd1 vssd1 vccd1 vccd1 _17864_/X sky130_fd_sc_hd__mux2_1
XFILLER_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10199_ _19287_/Q _19125_/Q _18534_/Q _18304_/Q _09868_/A _09927_/A vssd1 vssd1 vccd1
+ vccd1 _10200_/B sky130_fd_sc_hd__mux4_1
XFILLER_94_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_99_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19695_/CLK sky130_fd_sc_hd__clkbuf_16
X_19603_ _19603_/CLK _19603_/D vssd1 vssd1 vccd1 vccd1 _19603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16815_ _16816_/B _16810_/C _19578_/Q vssd1 vssd1 vccd1 vccd1 _16817_/B sky130_fd_sc_hd__a21oi_1
XFILLER_38_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17795_ _17795_/A vssd1 vssd1 vccd1 vccd1 _17795_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19534_ _19541_/CLK _19534_/D vssd1 vssd1 vccd1 vccd1 _19534_/Q sky130_fd_sc_hd__dfxtp_1
X_16746_ _16806_/A vssd1 vssd1 vccd1 vccd1 _16799_/A sky130_fd_sc_hd__clkbuf_2
X_13958_ _13958_/A vssd1 vssd1 vccd1 vccd1 _18515_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19465_ _19603_/CLK _19465_/D vssd1 vssd1 vccd1 vccd1 _19465_/Q sky130_fd_sc_hd__dfxtp_1
X_12909_ _12907_/X _18288_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12910_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_22_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19296_/CLK sky130_fd_sc_hd__clkbuf_16
X_16677_ _16681_/C _16681_/D _16676_/Y vssd1 vssd1 vccd1 vccd1 _19534_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14059__S _14063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13889_ _14569_/A vssd1 vssd1 vccd1 vccd1 _13889_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18416_ _19071_/CLK _18416_/D vssd1 vssd1 vccd1 vccd1 _18416_/Q sky130_fd_sc_hd__dfxtp_1
X_15628_ _15628_/A vssd1 vssd1 vccd1 vccd1 _19167_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19396_ _19699_/CLK _19396_/D vssd1 vssd1 vccd1 vccd1 _19396_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__12087__B _17215_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18347_ _19387_/CLK _18347_/D vssd1 vssd1 vccd1 vccd1 _18347_/Q sky130_fd_sc_hd__dfxtp_1
X_15559_ _19724_/Q _12577_/B _15569_/S vssd1 vssd1 vccd1 vccd1 _15559_/X sky130_fd_sc_hd__mux2_1
XFILLER_148_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11330__S0 _10692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__A1 _11288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19261_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16174__A0 _13519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ _09186_/B vssd1 vssd1 vccd1 vccd1 _09146_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18278_ _19725_/CLK _18278_/D vssd1 vssd1 vccd1 vccd1 _18278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 io_ibus_inst[15] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17229_ _17210_/X _17227_/X _17456_/S vssd1 vssd1 vccd1 vccd1 _17229_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput51 io_ibus_inst[25] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12735__A0 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput62 io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
XFILLER_116_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10746__C1 _11307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09982_ _09982_/A vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12831__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15353__S _15361_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10372__S1 _10229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _09416_/A vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__buf_2
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_34_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17788__B _17790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09347_ _11584_/B _09347_/B _17126_/C vssd1 vssd1 vccd1 vccd1 _11647_/B sky130_fd_sc_hd__or3_1
XFILLER_12_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10124__S1 _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09587__A _10660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09278_ _19829_/Q _12508_/B _12508_/C _19830_/Q vssd1 vssd1 vccd1 vccd1 _12606_/B
+ sky130_fd_sc_hd__or4b_4
XFILLER_138_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17901__A1 _17466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_3_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11240_ _18912_/Q _18678_/Q _19360_/Q _19008_/Q _11173_/S _11124_/X vssd1 vssd1 vccd1
+ vccd1 _11240_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10737__C1 _11307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10201__A1 _10195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11171_ _11171_/A _11171_/B vssd1 vssd1 vccd1 vccd1 _11171_/X sky130_fd_sc_hd__or2_1
XFILLER_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10122_ _10129_/A _10121_/X _09767_/A vssd1 vssd1 vccd1 vccd1 _10122_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09526__S _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17028__B _17133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11357__A _11357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ _18508_/Q _19003_/Q _10785_/S vssd1 vssd1 vccd1 vccd1 _10054_/A sky130_fd_sc_hd__mux2_1
X_14930_ _18911_/Q _14048_/X _14930_/S vssd1 vssd1 vccd1 vccd1 _14931_/A sky130_fd_sc_hd__mux2_1
XFILLER_88_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10261__A _10261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17968__A1 _19790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input26_A io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__S _12887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14861_ _14917_/A vssd1 vssd1 vccd1 vccd1 _14930_/S sky130_fd_sc_hd__buf_8
XFILLER_36_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16600_ _19513_/Q _16598_/B _16599_/Y vssd1 vssd1 vccd1 vccd1 _19513_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13812_ _13191_/X _18469_/Q _13820_/S vssd1 vssd1 vccd1 vccd1 _13813_/A sky130_fd_sc_hd__mux2_1
X_17580_ _17479_/X _17579_/X _17483_/X vssd1 vssd1 vccd1 vccd1 _17580_/Y sky130_fd_sc_hd__a21oi_1
X_14792_ _14792_/A vssd1 vssd1 vccd1 vccd1 _18848_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16531_ _16589_/A vssd1 vssd1 vccd1 vccd1 _16714_/A sky130_fd_sc_hd__clkbuf_2
X_13743_ _13228_/X _18439_/Q _13747_/S vssd1 vssd1 vccd1 vccd1 _13744_/A sky130_fd_sc_hd__mux2_1
X_10955_ _19272_/Q _19110_/Q _18519_/Q _18289_/Q _11196_/S _10934_/A vssd1 vssd1 vccd1
+ vccd1 _10956_/B sky130_fd_sc_hd__mux4_1
XFILLER_44_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16928__C1 _16269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19250_ _19250_/CLK _19250_/D vssd1 vssd1 vccd1 vccd1 _19250_/Q sky130_fd_sc_hd__dfxtp_1
X_16462_ _16470_/A _16466_/C vssd1 vssd1 vccd1 vccd1 _16462_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13206__A1 input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13674_ _13674_/A vssd1 vssd1 vccd1 vccd1 _18408_/D sky130_fd_sc_hd__clkbuf_1
X_10886_ _19177_/Q _18791_/Q _19241_/Q _18360_/Q _11172_/S _10817_/X vssd1 vssd1 vccd1
+ vccd1 _10887_/B sky130_fd_sc_hd__mux4_1
X_18201_ input39/X _18197_/X _18188_/X _18193_/X _11566_/A vssd1 vssd1 vccd1 vccd1
+ _18202_/B sky130_fd_sc_hd__a32o_1
X_15413_ _15459_/S vssd1 vssd1 vccd1 vccd1 _15422_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__15499__A _18258_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19181_ _19245_/CLK _19181_/D vssd1 vssd1 vccd1 vccd1 _19181_/Q sky130_fd_sc_hd__dfxtp_1
X_12625_ _17149_/A vssd1 vssd1 vccd1 vccd1 _18099_/A sky130_fd_sc_hd__clkbuf_4
X_16393_ _19447_/Q _16396_/C _16392_/Y vssd1 vssd1 vccd1 vccd1 _19447_/D sky130_fd_sc_hd__o21a_1
XANTENNA__11312__S0 _10660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ _18132_/A _18135_/B vssd1 vssd1 vccd1 vccd1 _18132_/X sky130_fd_sc_hd__or2_1
XFILLER_12_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09497__A _10854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12556_ _16301_/A vssd1 vssd1 vccd1 vccd1 _12556_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_106_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15344_ _19083_/Q _15035_/X _15350_/S vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _11507_/A vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18063_ _18229_/A vssd1 vssd1 vccd1 vccd1 _18066_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10436__A _10436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ _15275_/A vssd1 vssd1 vccd1 vccd1 _19052_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12487_ _17294_/S _12487_/B vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__nor2_1
XFILLER_172_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17014_ _19658_/Q _17024_/B vssd1 vssd1 vccd1 vccd1 _17014_/X sky130_fd_sc_hd__or2_1
XANTENNA_output94_A _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14226_ _14226_/A vssd1 vssd1 vccd1 vccd1 _18620_/D sky130_fd_sc_hd__clkbuf_1
X_11438_ _11441_/A _11439_/C _11439_/A vssd1 vssd1 vccd1 vccd1 _11438_/X sky130_fd_sc_hd__a21o_1
XFILLER_99_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12193__A1 _11354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15438__S _15444_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14157_ _14157_/A vssd1 vssd1 vccd1 vccd1 _18590_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17219__A _17219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11369_ _19297_/Q _19135_/Q _18544_/Q _18314_/Q _11374_/S _09733_/X vssd1 vssd1 vccd1
+ vccd1 _11369_/X sky130_fd_sc_hd__mux4_1
XFILLER_153_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11940__A1 _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13275_/A vssd1 vssd1 vccd1 vccd1 _13172_/S sky130_fd_sc_hd__buf_4
X_18965_ _19096_/CLK _18965_/D vssd1 vssd1 vccd1 vccd1 _18965_/Q sky130_fd_sc_hd__dfxtp_1
X_14088_ _13889_/X _18560_/Q _14096_/S vssd1 vssd1 vccd1 vccd1 _14089_/A sky130_fd_sc_hd__mux2_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13039_ _13038_/X _18294_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13040_/A sky130_fd_sc_hd__mux2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _19737_/Q _17430_/X _17915_/X vssd1 vssd1 vccd1 vccd1 _19737_/D sky130_fd_sc_hd__o21a_1
XFILLER_113_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18896_ _19282_/CLK _18896_/D vssd1 vssd1 vccd1 vccd1 _18896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10051__S0 _10017_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09361__A2 _09322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17847_ _17659_/X _17844_/X _17846_/Y _17673_/A vssd1 vssd1 vccd1 vccd1 _17847_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09992__S0 _09850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17778_ _17724_/A _17775_/X _17777_/Y _17413_/A vssd1 vssd1 vccd1 vccd1 _17778_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14297__B _14297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19517_ _19549_/CLK _19517_/D vssd1 vssd1 vccd1 vccd1 _19517_/Q sky130_fd_sc_hd__dfxtp_1
X_16729_ _16731_/B _16731_/C _16728_/Y vssd1 vssd1 vccd1 vccd1 _19552_/D sky130_fd_sc_hd__o21a_1
XFILLER_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15901__S _15909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19448_ _19448_/CLK _19448_/D vssd1 vssd1 vccd1 vccd1 _19448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09201_ _19854_/Q _19814_/Q vssd1 vssd1 vccd1 vccd1 _09201_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_23_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19379_ _19379_/CLK _19379_/D vssd1 vssd1 vccd1 vccd1 _19379_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11303__S0 _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09132_ _09113_/A _18081_/A _09182_/C vssd1 vssd1 vccd1 vccd1 _11569_/A sky130_fd_sc_hd__and3b_2
XFILLER_147_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10431__A1 _10394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13381__A0 _19738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15348__S _15350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12561__A _13356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09965_ _19322_/Q _18734_/Q _18771_/Q _18345_/Q _10112_/S _10218_/A vssd1 vssd1 vccd1
+ vccd1 _09965_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11177__A _11177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ _10342_/A vssd1 vssd1 vccd1 vccd1 _09905_/A sky130_fd_sc_hd__clkbuf_4
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11905__A _19402_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_10_0_clock_A clkbuf_3_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12239__A2 _12472_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15811__S _15815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _19308_/Q _18720_/Q _18757_/Q _18331_/Q _10660_/A _09442_/A vssd1 vssd1 vccd1
+ vccd1 _10740_/X sky130_fd_sc_hd__mux4_1
XFILLER_129_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ _09589_/A _10670_/X _10547_/A vssd1 vssd1 vccd1 vccd1 _10671_/X sky130_fd_sc_hd__a21o_1
XFILLER_167_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12410_ _19421_/Q _19422_/Q _12410_/C vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__and3_1
XFILLER_43_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13331__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_167_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13390_ _12606_/A _12600_/B _13391_/D _12602_/B vssd1 vssd1 vccd1 vccd1 _13390_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10958__C1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12455__B _12455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10422__A1 _09728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12341_ _12340_/Y _12337_/Y _12341_/S vssd1 vssd1 vccd1 vccd1 _12341_/X sky130_fd_sc_hd__mux2_1
XFILLER_154_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15060_ _15060_/A vssd1 vssd1 vccd1 vccd1 _15060_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12272_ _12372_/A _12270_/Y _12293_/B _11653_/X vssd1 vssd1 vccd1 vccd1 _12272_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_153_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18142__B _18142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011_ _18532_/Q _14010_/X _14011_/S vssd1 vssd1 vccd1 vccd1 _14012_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13567__A _15051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ _18578_/Q _18849_/Q _19073_/Q _18817_/Q _11219_/S _11020_/A vssd1 vssd1 vccd1
+ vccd1 _11223_/X sky130_fd_sc_hd__mux4_1
XFILLER_135_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10281__S0 _10339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ _18388_/Q _18649_/Q _18548_/Q _18883_/Q _10904_/X _11033_/X vssd1 vssd1 vccd1
+ vccd1 _11155_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10105_ _10105_/A _10105_/B vssd1 vssd1 vccd1 vccd1 _10105_/X sky130_fd_sc_hd__or2_1
X_18750_ _19237_/CLK _18750_/D vssd1 vssd1 vccd1 vccd1 _18750_/Q sky130_fd_sc_hd__dfxtp_1
X_15962_ _13563_/X _19313_/Q _15970_/S vssd1 vssd1 vccd1 vccd1 _15963_/A sky130_fd_sc_hd__mux2_1
X_11085_ _11085_/A _11085_/B vssd1 vssd1 vccd1 vccd1 _11085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09780__A _10215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17701_ _17524_/X _17522_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17701_/X sky130_fd_sc_hd__mux2_1
X_14913_ _18903_/Q _14023_/X _14915_/S vssd1 vssd1 vccd1 vccd1 _14914_/A sky130_fd_sc_hd__mux2_1
X_10036_ _18604_/Q _18875_/Q _19099_/Q _18843_/Q _09441_/X _10031_/A vssd1 vssd1 vccd1
+ vccd1 _10036_/X sky130_fd_sc_hd__mux4_1
X_18681_ _19012_/CLK _18681_/D vssd1 vssd1 vccd1 vccd1 _18681_/Q sky130_fd_sc_hd__dfxtp_1
X_15893_ _15893_/A vssd1 vssd1 vccd1 vccd1 _19282_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10584__S1 _10577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17632_ _17626_/X _17629_/X _17631_/Y _17589_/X vssd1 vssd1 vccd1 vccd1 _17632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_76_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14844_ _14844_/A vssd1 vssd1 vccd1 vccd1 _18872_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17563_ _17563_/A _17563_/B vssd1 vssd1 vccd1 vccd1 _17563_/Y sky130_fd_sc_hd__nor2_1
XFILLER_17_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14775_ _14605_/X _18842_/Q _14781_/S vssd1 vssd1 vccd1 vccd1 _14776_/A sky130_fd_sc_hd__mux2_1
X_11987_ _11987_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _11988_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10336__S1 _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15721__S _15721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19302_ _19302_/CLK _19302_/D vssd1 vssd1 vccd1 vccd1 _19302_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16514_ _19607_/Q _19609_/Q _19608_/Q _16882_/A vssd1 vssd1 vccd1 vccd1 _16891_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_72_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13726_ _13726_/A vssd1 vssd1 vccd1 vccd1 _18431_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17494_ _17530_/A vssd1 vssd1 vccd1 vccd1 _17494_/X sky130_fd_sc_hd__clkbuf_2
X_10938_ _18779_/Q vssd1 vssd1 vccd1 vccd1 _11241_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_44_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19233_ _19329_/CLK _19233_/D vssd1 vssd1 vccd1 vccd1 _19233_/Q sky130_fd_sc_hd__dfxtp_1
X_16445_ _19465_/Q _16442_/B _16444_/Y vssd1 vssd1 vccd1 vccd1 _19465_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14337__S _14343_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13657_ _13657_/A vssd1 vssd1 vccd1 vccd1 _18400_/D sky130_fd_sc_hd__clkbuf_1
X_10869_ _11291_/A _12453_/A vssd1 vssd1 vccd1 vccd1 _11461_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13241__S _13252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12938__B1 _12936_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15022__A _15022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _19620_/Q _12619_/A _12605_/Y _19663_/Q _12607_/X vssd1 vssd1 vccd1 vccd1
+ _12608_/X sky130_fd_sc_hd__a221o_1
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19164_ _19598_/CLK _19164_/D vssd1 vssd1 vccd1 vccd1 _19164_/Q sky130_fd_sc_hd__dfxtp_1
X_16376_ _19441_/Q _16379_/C _16359_/X vssd1 vssd1 vccd1 vccd1 _16376_/Y sky130_fd_sc_hd__a21oi_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13588_ _13588_/A vssd1 vssd1 vccd1 vccd1 _18375_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18115_ _19821_/Q _18106_/X _18114_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _19821_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_9_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15327_ _15327_/A vssd1 vssd1 vccd1 vccd1 _19075_/D sky130_fd_sc_hd__clkbuf_1
X_12539_ _19568_/Q _12518_/X _12535_/X _12538_/X vssd1 vssd1 vccd1 vccd1 _12539_/X
+ sky130_fd_sc_hd__a211o_1
X_19095_ _19127_/CLK _19095_/D vssd1 vssd1 vccd1 vccd1 _19095_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18046_ _19793_/Q _19414_/Q _18050_/S vssd1 vssd1 vccd1 vccd1 _18047_/A sky130_fd_sc_hd__mux2_1
X_15258_ _15315_/S vssd1 vssd1 vccd1 vccd1 _15267_/S sky130_fd_sc_hd__buf_2
XFILLER_126_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_173_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14209_ _18613_/Q _13962_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14210_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14072__S _14074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15189_ _19014_/Q _15019_/X _15195_/S vssd1 vssd1 vccd1 vccd1 _15190_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15104__A1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09750_ _11380_/A _09750_/B vssd1 vssd1 vccd1 vccd1 _09750_/X sky130_fd_sc_hd__or2_1
XFILLER_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18948_ _19076_/CLK _18948_/D vssd1 vssd1 vccd1 vccd1 _18948_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09690__A _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _09681_/A vssd1 vssd1 vccd1 vccd1 _09682_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09965__S0 _10112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__B1 _09756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18879_ _19297_/CLK _18879_/D vssd1 vssd1 vccd1 vccd1 _18879_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11429__B1 _12473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17565__C1 _17532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12556__A _16301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _17120_/B _09171_/B _17120_/C vssd1 vssd1 vccd1 vccd1 _09116_/A sky130_fd_sc_hd__and3_1
XFILLER_129_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15867__A _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__B1 _11600_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15586__B _15586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17096__A1 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09948_ _09844_/X _09941_/X _09943_/X _09947_/X _09754_/A vssd1 vssd1 vccd1 vccd1
+ _09948_/X sky130_fd_sc_hd__a311o_2
XFILLER_104_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10015__S _10572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _10520_/S vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__buf_2
XFILLER_46_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _19338_/Q _12068_/A _13411_/A vssd1 vssd1 vccd1 vccd1 _11910_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_58_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12890_ _16011_/B _12891_/C _16021_/A vssd1 vssd1 vccd1 vccd1 _12892_/A sky130_fd_sc_hd__a21oi_1
XFILLER_173_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10749__A_N _12455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10891__A1 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__B _12470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _17605_/A vssd1 vssd1 vccd1 vccd1 _11842_/D sky130_fd_sc_hd__inv_2
XFILLER_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _19333_/Q _11766_/X _11734_/X _11771_/X _11691_/X vssd1 vssd1 vccd1 vccd1
+ _11772_/X sky130_fd_sc_hd__o221a_1
X_14560_ _14560_/A vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _16619_/D vssd1 vssd1 vccd1 vccd1 _13619_/C sky130_fd_sc_hd__inv_2
X_10723_ _09632_/A _10722_/X _09630_/A vssd1 vssd1 vccd1 vccd1 _10723_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14491_ _14502_/A vssd1 vssd1 vccd1 vccd1 _14500_/S sky130_fd_sc_hd__buf_4
XFILLER_41_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16230_ _16230_/A vssd1 vssd1 vccd1 vccd1 _19386_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_110_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13442_ _12828_/X _18322_/Q _13448_/S vssd1 vssd1 vccd1 vccd1 _13443_/A sky130_fd_sc_hd__mux2_1
X_10654_ _10654_/A vssd1 vssd1 vccd1 vccd1 _10729_/S sky130_fd_sc_hd__buf_4
XFILLER_167_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13373_ _19487_/Q vssd1 vssd1 vccd1 vccd1 _16321_/B sky130_fd_sc_hd__clkbuf_2
X_16161_ _16165_/B _16161_/B vssd1 vssd1 vccd1 vccd1 _16161_/Y sky130_fd_sc_hd__nand2_1
XFILLER_103_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10585_ _10585_/A _10585_/B vssd1 vssd1 vccd1 vccd1 _10585_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18153__A _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15112_ _18980_/Q _15012_/X _15112_/S vssd1 vssd1 vccd1 vccd1 _15113_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12324_ _19354_/Q _12069_/X _12323_/X _12075_/X vssd1 vssd1 vccd1 vccd1 _12324_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_6_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16092_ _16091_/A _16091_/C _16091_/B vssd1 vssd1 vccd1 vccd1 _16092_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13345__A0 _19736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12255_ _19351_/Q _11733_/X _12037_/X _12254_/X _12102_/X vssd1 vssd1 vccd1 vccd1
+ _12255_/X sky130_fd_sc_hd__o221a_1
XFILLER_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15043_ _15043_/A vssd1 vssd1 vccd1 vccd1 _18957_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_3_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11206_ _11252_/A _11206_/B vssd1 vssd1 vccd1 vccd1 _11206_/X sky130_fd_sc_hd__or2_1
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19851_ _19854_/CLK _19851_/D vssd1 vssd1 vccd1 vccd1 _19851_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12186_ _12183_/X _12185_/Y _11623_/X vssd1 vssd1 vccd1 vccd1 _12186_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_156_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18802_ _19378_/CLK _18802_/D vssd1 vssd1 vccd1 vccd1 _18802_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11137_ _19172_/Q _18786_/Q _19236_/Q _18355_/Q _11173_/S _10817_/A vssd1 vssd1 vccd1
+ vccd1 _11138_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19782_ _19786_/CLK _19782_/D vssd1 vssd1 vccd1 vccd1 _19782_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_95_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16994_ _18172_/A vssd1 vssd1 vccd1 vccd1 _18097_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18733_ _19256_/CLK _18733_/D vssd1 vssd1 vccd1 vccd1 _18733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11068_ _11171_/A _11067_/X _09447_/A vssd1 vssd1 vccd1 vccd1 _11068_/X sky130_fd_sc_hd__o21a_1
X_15945_ _15945_/A vssd1 vssd1 vccd1 vccd1 _19305_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10019_ _10575_/A vssd1 vssd1 vccd1 vccd1 _10684_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18664_ _19284_/CLK _18664_/D vssd1 vssd1 vccd1 vccd1 _18664_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15876_ _19275_/Q _14550_/A _15876_/S vssd1 vssd1 vccd1 vccd1 _15877_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17615_ _17615_/A _17615_/B vssd1 vssd1 vccd1 vccd1 _17615_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14827_ _14827_/A vssd1 vssd1 vccd1 vccd1 _18864_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18595_ _19091_/CLK _18595_/D vssd1 vssd1 vccd1 vccd1 _18595_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15451__S _15455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17232__A _17232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17546_ _11732_/X _17427_/X _09359_/X vssd1 vssd1 vccd1 vccd1 _17546_/X sky130_fd_sc_hd__a21o_1
X_14758_ _14758_/A vssd1 vssd1 vccd1 vccd1 _18834_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _13709_/A vssd1 vssd1 vccd1 vccd1 _18423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17477_ _17860_/A vssd1 vssd1 vccd1 vccd1 _17477_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14689_ _14700_/A vssd1 vssd1 vccd1 vccd1 _14698_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_20_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19216_ _19248_/CLK _19216_/D vssd1 vssd1 vccd1 vccd1 _19216_/Q sky130_fd_sc_hd__dfxtp_1
X_16428_ _19459_/Q _16425_/B _16427_/Y vssd1 vssd1 vccd1 vccd1 _19459_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17886__B _17886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12095__B _19401_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19147_ _19796_/CLK _19147_/D vssd1 vssd1 vccd1 vccd1 _19147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16359_ _16546_/A vssd1 vssd1 vccd1 vccd1 _16359_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09685__A _10093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19078_ _19367_/CLK _19078_/D vssd1 vssd1 vccd1 vccd1 _19078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18029_ _18029_/A vssd1 vssd1 vccd1 vccd1 _18038_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__12542__C _12542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09802_ _18413_/Q _18674_/Q _18573_/Q _18908_/Q _11385_/S _09799_/X vssd1 vssd1 vccd1
+ vccd1 _09802_/X sky130_fd_sc_hd__mux4_1
XFILLER_140_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09733_ _09733_/A vssd1 vssd1 vccd1 vccd1 _09733_/X sky130_fd_sc_hd__buf_2
XFILLER_28_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09664_ _09664_/A vssd1 vssd1 vccd1 vccd1 _09664_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09595_ _09717_/A _09595_/B vssd1 vssd1 vccd1 vccd1 _09595_/X sky130_fd_sc_hd__or2_1
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15261__A0 _14541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15361__S _15361_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17002__A1 _15588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__A1 _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_126_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12286__A _12286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10720__S1 _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14705__S _14709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10370_ _09713_/A _10367_/X _10369_/X vssd1 vssd1 vccd1 vccd1 _10370_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10484__S0 _10274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13327__B1 _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11338__C1 _09572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12040_ _12040_/A _12065_/B vssd1 vssd1 vccd1 vccd1 _12040_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11349__B _12465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17317__A _17317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_93_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13991_ _14563_/A vssd1 vssd1 vccd1 vccd1 _13991_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ _13541_/X _19210_/Q _15732_/S vssd1 vssd1 vccd1 vccd1 _15731_/A sky130_fd_sc_hd__mux2_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _12929_/Y _12941_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12942_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _15661_/A vssd1 vssd1 vccd1 vccd1 _19179_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12873_ _19556_/Q vssd1 vssd1 vccd1 vccd1 _16752_/D sky130_fd_sc_hd__buf_2
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17577_/S _17398_/X _17399_/Y vssd1 vssd1 vccd1 vccd1 _17400_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14612_ _14611_/X _18775_/Q _14615_/S vssd1 vssd1 vccd1 vccd1 _14613_/A sky130_fd_sc_hd__mux2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ _11824_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11824_/Y sky130_fd_sc_hd__xnor2_4
X_18380_ _19197_/CLK _18380_/D vssd1 vssd1 vccd1 vccd1 _18380_/Q sky130_fd_sc_hd__dfxtp_1
X_15592_ _19730_/Q _12689_/X _15595_/S vssd1 vssd1 vccd1 vccd1 _15592_/X sky130_fd_sc_hd__mux2_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17331_ _17404_/B _17432_/B _17190_/A vssd1 vssd1 vccd1 vccd1 _17541_/A sky130_fd_sc_hd__nor3b_2
X_14543_ _14543_/A vssd1 vssd1 vccd1 vccd1 _18753_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11755_ _11755_/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11813_/A sky130_fd_sc_hd__and2_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_82_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17262_ _17260_/X _17261_/X _17266_/A vssd1 vssd1 vccd1 vccd1 _17262_/X sky130_fd_sc_hd__mux2_1
X_10706_ _18619_/Q _18954_/Q _11320_/S vssd1 vssd1 vccd1 vccd1 _10706_/X sky130_fd_sc_hd__mux2_1
XFILLER_159_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ _13880_/X _18722_/Q _14478_/S vssd1 vssd1 vccd1 vccd1 _14475_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11686_ _12037_/A vssd1 vssd1 vccd1 vccd1 _11686_/X sky130_fd_sc_hd__buf_2
XFILLER_174_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19001_ _19385_/CLK _19001_/D vssd1 vssd1 vccd1 vccd1 _19001_/Q sky130_fd_sc_hd__dfxtp_1
X_16213_ _13576_/X _19379_/Q _16213_/S vssd1 vssd1 vccd1 vccd1 _16214_/A sky130_fd_sc_hd__mux2_1
X_13425_ _13425_/A vssd1 vssd1 vccd1 vccd1 _18319_/D sky130_fd_sc_hd__clkbuf_1
X_17193_ _17471_/B vssd1 vssd1 vccd1 vccd1 _17737_/A sky130_fd_sc_hd__clkbuf_2
X_10637_ _10689_/A _10637_/B vssd1 vssd1 vccd1 vccd1 _10637_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14615__S _14615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16144_ _16150_/B _16143_/Y _16109_/X vssd1 vssd1 vccd1 vccd1 _16144_/Y sky130_fd_sc_hd__a21oi_1
X_13356_ _19486_/Q _13356_/B vssd1 vssd1 vccd1 vccd1 _13356_/X sky130_fd_sc_hd__and2_1
X_10568_ _18926_/Q _18692_/Q _19374_/Q _19022_/Q _10566_/X _10567_/X vssd1 vssd1 vccd1
+ vccd1 _10569_/B sky130_fd_sc_hd__mux4_1
XFILLER_128_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12307_ _17867_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__xnor2_1
XFILLER_170_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16075_ _16080_/B _16075_/B vssd1 vssd1 vccd1 vccd1 _16075_/Y sky130_fd_sc_hd__nand2_1
X_13287_ _19450_/Q _12962_/X _13286_/X vssd1 vssd1 vccd1 vccd1 _13287_/X sky130_fd_sc_hd__o21a_1
X_10499_ _18624_/Q _18959_/Q _10499_/S vssd1 vssd1 vccd1 vccd1 _10499_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11329__C1 _09658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15026_ _18952_/Q _15025_/X _15029_/S vssd1 vssd1 vccd1 vccd1 _15027_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12238_ _11618_/A _11507_/A _12302_/A vssd1 vssd1 vccd1 vccd1 _12238_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10001__C1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__S1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19834_ _19834_/CLK _19834_/D vssd1 vssd1 vccd1 vccd1 _19834_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14350__S _14354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _12169_/A vssd1 vssd1 vccd1 vccd1 _12173_/A sky130_fd_sc_hd__clkinv_2
XFILLER_122_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16977_ _15536_/X _16970_/X _16976_/X _16968_/X vssd1 vssd1 vccd1 vccd1 _19644_/D
+ sky130_fd_sc_hd__o211a_1
X_19765_ _19793_/CLK _19765_/D vssd1 vssd1 vccd1 vccd1 _19765_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13097__A2 _12817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14294__A1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14294__B2 _18130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput5 io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_18716_ _19305_/CLK _18716_/D vssd1 vssd1 vccd1 vccd1 _18716_/Q sky130_fd_sc_hd__dfxtp_1
X_15928_ _15996_/S vssd1 vssd1 vccd1 vccd1 _15937_/S sky130_fd_sc_hd__clkbuf_4
X_19696_ _19845_/CLK _19696_/D vssd1 vssd1 vccd1 vccd1 _19696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18647_ _19299_/CLK _18647_/D vssd1 vssd1 vccd1 vccd1 _18647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15859_ _19267_/Q _14525_/A _15865_/S vssd1 vssd1 vccd1 vccd1 _15860_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14586__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10950__S1 _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _09380_/A vssd1 vssd1 vccd1 vccd1 _10031_/A sky130_fd_sc_hd__clkbuf_4
X_18578_ _19712_/CLK _18578_/D vssd1 vssd1 vccd1 vccd1 _18578_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17529_ _17392_/X _17684_/A _17402_/X vssd1 vssd1 vccd1 vccd1 _17529_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_33_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09473__A1 _09665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__B2 _19736_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11280__A1 _11116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12553__B _18079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14260__S _14264_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15482__A0 _19711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09716_ _18940_/Q _18706_/Q _19388_/Q _19036_/Q _09704_/X _09715_/X vssd1 vssd1 vccd1
+ vccd1 _09716_/X sky130_fd_sc_hd__mux4_1
XFILLER_55_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17223__A1 _17790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11194__S1 _11177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ _10640_/A vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_104_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09578_ _09578_/A vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12728__B _12730_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15537__A1 _15536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11540_ _11540_/A vssd1 vssd1 vccd1 vccd1 _18744_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ _11461_/Y _11462_/Y _11463_/Y _11461_/B _11470_/X vssd1 vssd1 vccd1 vccd1
+ _11471_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14435__S _14439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09216__A1 _09331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12744__A _12744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13210_ _13209_/X _18304_/Q _13252_/S vssd1 vssd1 vccd1 vccd1 _13211_/A sky130_fd_sc_hd__mux2_1
X_10422_ _09728_/A _10417_/X _10419_/X _10421_/X _09669_/A vssd1 vssd1 vccd1 vccd1
+ _10422_/X sky130_fd_sc_hd__a221o_4
XANTENNA__11023__A1 _11116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14190_ _14190_/A vssd1 vssd1 vccd1 vccd1 _18605_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_100_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10353_ _19726_/Q vssd1 vssd1 vccd1 vccd1 _10353_/Y sky130_fd_sc_hd__inv_2
X_13141_ _19757_/Q vssd1 vssd1 vccd1 vccd1 _16091_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13072_ _13072_/A vssd1 vssd1 vccd1 vccd1 _18296_/D sky130_fd_sc_hd__clkbuf_1
X_10284_ _09765_/A _10265_/Y _10273_/X _10283_/Y _09813_/A vssd1 vssd1 vccd1 vccd1
+ _10284_/X sky130_fd_sc_hd__o311a_4
XANTENNA_input56_A io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16900_ _16915_/A _16904_/C vssd1 vssd1 vccd1 vccd1 _16900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12023_ _18107_/A _12021_/X _12022_/X vssd1 vssd1 vccd1 vccd1 _12023_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_2_0_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_17880_ _17626_/X _17877_/X _17879_/Y _17532_/A vssd1 vssd1 vccd1 vccd1 _17880_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_120_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16831_ _16833_/A _16831_/B vssd1 vssd1 vccd1 vccd1 _19583_/D sky130_fd_sc_hd__nor2_1
XFILLER_116_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19550_ _19550_/CLK _19550_/D vssd1 vssd1 vccd1 vccd1 _19550_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16762_ _16762_/A _16772_/D vssd1 vssd1 vccd1 vccd1 _16762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13974_ _13974_/A vssd1 vssd1 vccd1 vccd1 _18520_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12826__A2 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18501_ _18569_/CLK _18501_/D vssd1 vssd1 vccd1 vccd1 _18501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15713_ _13509_/X _19202_/Q _15721_/S vssd1 vssd1 vccd1 vccd1 _15714_/A sky130_fd_sc_hd__mux2_1
X_19481_ _19491_/CLK _19481_/D vssd1 vssd1 vccd1 vccd1 _19481_/Q sky130_fd_sc_hd__dfxtp_1
X_12925_ _12924_/X _18289_/Q _13000_/S vssd1 vssd1 vccd1 vccd1 _12926_/A sky130_fd_sc_hd__mux2_1
X_16693_ _16697_/C _16697_/D _16692_/Y vssd1 vssd1 vccd1 vccd1 _19540_/D sky130_fd_sc_hd__o21a_1
XFILLER_47_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10301__A3 _10299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18432_ _19314_/CLK _18432_/D vssd1 vssd1 vccd1 vccd1 _18432_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15644_ _15644_/A vssd1 vssd1 vccd1 vccd1 _19171_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12856_ _19741_/Q _19742_/Q vssd1 vssd1 vccd1 vccd1 _12891_/C sky130_fd_sc_hd__and2_2
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11807_ _19636_/Q _13423_/A vssd1 vssd1 vccd1 vccd1 _11807_/Y sky130_fd_sc_hd__nor2_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _19180_/CLK _18363_/D vssd1 vssd1 vccd1 vccd1 _18363_/Q sky130_fd_sc_hd__dfxtp_1
X_15575_ _15601_/A vssd1 vssd1 vccd1 vccd1 _15595_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12787_ _16731_/B _12638_/X _12786_/X _12644_/X vssd1 vssd1 vccd1 vccd1 _12787_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_15_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11034__S _11071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _12482_/A _17120_/A _17115_/A _18104_/A vssd1 vssd1 vccd1 vccd1 _17485_/A
+ sky130_fd_sc_hd__o211a_2
XANTENNA__15528__A1 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14526_ _14525_/X _18748_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14527_/A sky130_fd_sc_hd__mux2_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18294_ _19184_/CLK _18294_/D vssd1 vssd1 vccd1 vccd1 _18294_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10696__S0 _10579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11738_ _11738_/A vssd1 vssd1 vccd1 vccd1 _14275_/B sky130_fd_sc_hd__buf_2
X_17245_ _17245_/A vssd1 vssd1 vccd1 vccd1 _17605_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_14457_ _14457_/A vssd1 vssd1 vccd1 vccd1 _18714_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10873__S _10873_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ _11840_/A _11669_/B vssd1 vssd1 vccd1 vccd1 _11676_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11014__A1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13408_ _18252_/Q _13408_/B vssd1 vssd1 vccd1 vccd1 _13408_/X sky130_fd_sc_hd__or2_1
X_17176_ _17176_/A _17176_/B _17176_/C _17176_/D vssd1 vssd1 vccd1 vccd1 _17177_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_116_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14388_ _14388_/A vssd1 vssd1 vccd1 vccd1 _18683_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16127_ _16126_/A _16126_/C _13245_/A vssd1 vssd1 vccd1 vccd1 _16127_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_143_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13339_ _19693_/Q _12529_/A _12521_/A _19660_/Q vssd1 vssd1 vccd1 vccd1 _13339_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_142_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10174__A _10174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17150__B1 _17140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_142_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16058_ _16086_/A vssd1 vssd1 vccd1 vccd1 _16082_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11317__A2 _11307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ _15009_/A vssd1 vssd1 vccd1 vccd1 _15009_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15176__S _15184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19817_ _19834_/CLK _19817_/D vssd1 vssd1 vccd1 vccd1 _19817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10540__A3 _10538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19748_ _19779_/CLK _19748_/D vssd1 vssd1 vccd1 vccd1 _19748_/Q sky130_fd_sc_hd__dfxtp_1
X_09501_ _18642_/Q vssd1 vssd1 vccd1 vccd1 _11033_/A sky130_fd_sc_hd__buf_2
X_19679_ _19688_/CLK _19679_/D vssd1 vssd1 vccd1 vccd1 _19679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09432_ _09432_/A vssd1 vssd1 vccd1 vccd1 _09608_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09363_ _17117_/B vssd1 vssd1 vccd1 vccd1 _11491_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_80_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _16619_/B _12621_/B vssd1 vssd1 vccd1 vccd1 _11805_/C sky130_fd_sc_hd__nor2_1
XFILLER_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10783__S _11318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12753__A1 hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17141__B1 _17140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput150 _16282_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[17] sky130_fd_sc_hd__buf_2
Xoutput161 _16302_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[27] sky130_fd_sc_hd__buf_2
XFILLER_133_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput172 _16260_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_30_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12730__C _12730_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10611__S0 _10546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10971_ _10971_/A vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__buf_4
XFILLER_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12739__A _12744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12710_ _19544_/Q _12939_/S _12699_/X _19512_/Q _12709_/X vssd1 vssd1 vccd1 vccd1
+ _12710_/X sky130_fd_sc_hd__a221o_1
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_3_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19280_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_71_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13690_ _13386_/X _18416_/Q _13690_/S vssd1 vssd1 vccd1 vccd1 _13691_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12641_ _19586_/Q _12660_/B vssd1 vssd1 vccd1 vccd1 _12641_/X sky130_fd_sc_hd__and2_1
XANTENNA__11362__B _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11244__A1 _11005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12177__C _19412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15360_ _15360_/A vssd1 vssd1 vccd1 vccd1 _19090_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12572_ _18268_/Q _13132_/B _13132_/C _12571_/Y vssd1 vssd1 vccd1 vccd1 _12572_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17904__C1 _12744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14311_ _14311_/A vssd1 vssd1 vccd1 vccd1 _18650_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12992__A1 _15513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ _18087_/A _11620_/A _11523_/C _11523_/D vssd1 vssd1 vccd1 vccd1 _11523_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__14165__S _14169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15291_ _15302_/A vssd1 vssd1 vccd1 vccd1 _15300_/S sky130_fd_sc_hd__buf_4
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17030_ _17098_/S vssd1 vssd1 vccd1 vccd1 _17039_/S sky130_fd_sc_hd__buf_2
X_14242_ _18628_/Q _14010_/X _14242_/S vssd1 vssd1 vccd1 vccd1 _14243_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11454_ _10649_/A _11453_/Y _11344_/Y vssd1 vssd1 vccd1 vccd1 _11454_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_172_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10405_ _19187_/Q _18801_/Q _19251_/Q _18370_/Q _10450_/S _10238_/A vssd1 vssd1 vccd1
+ vccd1 _10406_/B sky130_fd_sc_hd__mux4_1
X_14173_ _14173_/A vssd1 vssd1 vccd1 vccd1 _18597_/D sky130_fd_sc_hd__clkbuf_1
X_11385_ _18512_/Q _19007_/Q _11385_/S vssd1 vssd1 vccd1 vccd1 _11386_/A sky130_fd_sc_hd__mux2_1
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13124_ _14573_/A vssd1 vssd1 vccd1 vccd1 _13124_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10336_ _19285_/Q _19123_/Q _18532_/Q _18302_/Q _10286_/X _10382_/A vssd1 vssd1 vccd1
+ vccd1 _10336_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output162_A _12376_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18981_ _19109_/CLK _18981_/D vssd1 vssd1 vccd1 vccd1 _18981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13055_/A vssd1 vssd1 vccd1 vccd1 _13055_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10267_ _10481_/S vssd1 vssd1 vccd1 vccd1 _10435_/S sky130_fd_sc_hd__buf_2
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _17932_/A vssd1 vssd1 vccd1 vccd1 _19741_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12006_ _11956_/A _11983_/A _11985_/B vssd1 vssd1 vccd1 vccd1 _12006_/Y sky130_fd_sc_hd__a21oi_1
X_17863_ _19732_/Q _17831_/X _17862_/X vssd1 vssd1 vccd1 vccd1 _19732_/D sky130_fd_sc_hd__o21a_1
XFILLER_79_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10198_ _18470_/Q _19061_/Q _19223_/Q _18438_/Q _09931_/S _09871_/A vssd1 vssd1 vccd1
+ vccd1 _10198_/X sky130_fd_sc_hd__mux4_1
XFILLER_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19602_ _19603_/CLK _19602_/D vssd1 vssd1 vccd1 vccd1 _19602_/Q sky130_fd_sc_hd__dfxtp_1
X_16814_ _16816_/B _16810_/C _16813_/Y vssd1 vssd1 vccd1 vccd1 _19577_/D sky130_fd_sc_hd__o21a_1
X_17794_ _17571_/X _17692_/Y _17793_/X _17592_/X vssd1 vssd1 vccd1 vccd1 _17794_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_81_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16745_ _16752_/B _16742_/B _16744_/Y vssd1 vssd1 vccd1 vccd1 _19558_/D sky130_fd_sc_hd__o21a_1
X_19533_ _19541_/CLK _19533_/D vssd1 vssd1 vccd1 vccd1 _19533_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17199__A0 _17630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13957_ _18515_/Q _13956_/X _13963_/S vssd1 vssd1 vccd1 vccd1 _13958_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12649__A _18262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19464_ _19607_/CLK _19464_/D vssd1 vssd1 vccd1 vccd1 _19464_/Q sky130_fd_sc_hd__dfxtp_1
X_12908_ _13387_/S vssd1 vssd1 vccd1 vccd1 _13000_/S sky130_fd_sc_hd__buf_2
XANTENNA__15025__A _15025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16676_ _16681_/C _16681_/D _16675_/X vssd1 vssd1 vccd1 vccd1 _16676_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13888_ _13888_/A vssd1 vssd1 vccd1 vccd1 _18495_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15627_ _15626_/X _19167_/Q _15627_/S vssd1 vssd1 vccd1 vccd1 _15628_/A sky130_fd_sc_hd__mux2_1
X_18415_ _19328_/CLK _18415_/D vssd1 vssd1 vccd1 vccd1 _18415_/Q sky130_fd_sc_hd__dfxtp_1
X_12839_ _16736_/B _12518_/A _12838_/X _13012_/A vssd1 vssd1 vccd1 vccd1 _12839_/X
+ sky130_fd_sc_hd__a211o_1
X_19395_ _19699_/CLK _19395_/D vssd1 vssd1 vccd1 vccd1 _19395_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10169__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18346_ _19197_/CLK _18346_/D vssd1 vssd1 vccd1 vccd1 _18346_/Q sky130_fd_sc_hd__dfxtp_1
X_15558_ _15558_/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__clkbuf_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_159_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11330__S1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14509_ _13931_/X _18738_/Q _14511_/S vssd1 vssd1 vccd1 vccd1 _14510_/A sky130_fd_sc_hd__mux2_1
X_18277_ _19725_/CLK _18277_/D vssd1 vssd1 vccd1 vccd1 _18277_/Q sky130_fd_sc_hd__dfxtp_1
X_15489_ _19712_/Q _15487_/X _15516_/S vssd1 vssd1 vccd1 vccd1 _15489_/X sky130_fd_sc_hd__mux2_1
X_17228_ _17256_/A vssd1 vssd1 vccd1 vccd1 _17456_/S sky130_fd_sc_hd__clkbuf_2
Xinput30 io_dbus_rdata[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_4
Xinput41 io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
Xinput52 io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_2
XFILLER_128_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput63 io_ibus_inst[7] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__12735__A1 _11070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15695__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17159_ _12482_/B _17149_/X _17140_/X _19705_/Q vssd1 vssd1 vccd1 vccd1 _17160_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_115_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09981_ _18507_/Q _19002_/Q _09981_/S vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__mux2_1
XFILLER_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ _09415_/A vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__buf_2
XANTENNA__10079__A _10080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09346_ _11618_/A _11619_/A _17127_/A vssd1 vssd1 vccd1 vccd1 _09352_/A sky130_fd_sc_hd__or3_1
XFILLER_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_166_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _19828_/Q _19827_/Q vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__or2_1
XFILLER_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__A _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15809__S _15815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14713__S _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _18915_/Q _18681_/Q _19363_/Q _19011_/Q _11011_/X _11012_/X vssd1 vssd1 vccd1
+ vccd1 _11171_/B sky130_fd_sc_hd__mux4_1
XFILLER_161_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_3_7_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10121_ _18600_/Q _18871_/Q _19095_/Q _18839_/Q _09918_/X _09900_/A vssd1 vssd1 vccd1
+ vccd1 _10121_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10542__A _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10052_ _10684_/A _10052_/B vssd1 vssd1 vccd1 vccd1 _10052_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11357__B _12472_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__B1 _09561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18090__A1 _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ _18096_/A _14860_/B _18091_/A _14860_/D vssd1 vssd1 vccd1 vccd1 _14917_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_29_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13811_ _13822_/A vssd1 vssd1 vccd1 vccd1 _13820_/S sky130_fd_sc_hd__buf_4
XFILLER_17_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14791_ _18848_/Q _13943_/X _14799_/S vssd1 vssd1 vccd1 vccd1 _14792_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input19_A io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16530_ _16541_/A _16530_/B _16530_/C vssd1 vssd1 vccd1 vccd1 _19491_/D sky130_fd_sc_hd__nor3_1
XFILLER_17_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13742_ _13742_/A vssd1 vssd1 vccd1 vccd1 _18438_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_151_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19202_/CLK sky130_fd_sc_hd__clkbuf_16
X_10954_ _18455_/Q _19046_/Q _19208_/Q _18423_/Q _09396_/A _09416_/A vssd1 vssd1 vccd1
+ vccd1 _10954_/X sky130_fd_sc_hd__mux4_2
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13999__S _14011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16461_ _16461_/A vssd1 vssd1 vccd1 vccd1 _16466_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13673_ _13240_/X _18408_/Q _13675_/S vssd1 vssd1 vccd1 vccd1 _13674_/A sky130_fd_sc_hd__mux2_1
X_10885_ _09431_/A _10871_/X _10877_/X _10884_/X _10949_/A vssd1 vssd1 vccd1 vccd1
+ _10885_/X sky130_fd_sc_hd__a311o_1
XFILLER_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18200_ _18200_/A vssd1 vssd1 vccd1 vccd1 _19848_/D sky130_fd_sc_hd__clkbuf_1
X_15412_ _15412_/A vssd1 vssd1 vccd1 vccd1 _19113_/D sky130_fd_sc_hd__clkbuf_1
X_12624_ _17133_/B vssd1 vssd1 vccd1 vccd1 _17149_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__09778__A _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19180_ _19180_/CLK _19180_/D vssd1 vssd1 vccd1 vccd1 _19180_/Q sky130_fd_sc_hd__dfxtp_1
X_16392_ _19447_/Q _16396_/C _16359_/X vssd1 vssd1 vccd1 vccd1 _16392_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__15499__B _15499_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18131_ _19827_/Q _18120_/X _18130_/X _18123_/X vssd1 vssd1 vccd1 vccd1 _19827_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11312__S1 _10655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_166_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19720_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11820__B _17245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15343_ _15343_/A vssd1 vssd1 vccd1 vccd1 _19082_/D sky130_fd_sc_hd__clkbuf_1
X_12555_ _17102_/A vssd1 vssd1 vccd1 vccd1 _16301_/A sky130_fd_sc_hd__buf_2
XFILLER_8_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11506_ _12159_/A vssd1 vssd1 vccd1 vccd1 _11507_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18062_ _18062_/A vssd1 vssd1 vccd1 vccd1 _19800_/D sky130_fd_sc_hd__clkbuf_1
X_15274_ _14560_/X _19052_/Q _15278_/S vssd1 vssd1 vccd1 vccd1 _15275_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12486_ _17356_/S vssd1 vssd1 vccd1 vccd1 _17294_/S sky130_fd_sc_hd__buf_2
X_17013_ _17013_/A vssd1 vssd1 vccd1 vccd1 _17024_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15719__S _15721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14225_ _18620_/Q _13985_/X _14231_/S vssd1 vssd1 vccd1 vccd1 _14226_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11076__S0 _11265_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11437_ _11437_/A _11437_/B vssd1 vssd1 vccd1 vccd1 _11437_/Y sky130_fd_sc_hd__nand2_1
XFILLER_172_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14156_ _18590_/Q _13991_/X _14158_/S vssd1 vssd1 vccd1 vccd1 _14157_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output87_A _12269_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11368_ _11368_/A _11368_/B vssd1 vssd1 vccd1 vccd1 _11368_/X sky130_fd_sc_hd__or2_1
XFILLER_98_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13107_ _14569_/A vssd1 vssd1 vccd1 vccd1 _13107_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _09857_/A _10307_/X _10309_/X _09670_/A _10318_/X vssd1 vssd1 vccd1 vccd1
+ _10319_/X sky130_fd_sc_hd__a311o_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ _18964_/CLK _18964_/D vssd1 vssd1 vccd1 vccd1 _18964_/Q sky130_fd_sc_hd__dfxtp_1
X_14087_ _14109_/A vssd1 vssd1 vccd1 vccd1 _14096_/S sky130_fd_sc_hd__buf_4
XFILLER_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _18494_/Q _18989_/Q _11299_/S vssd1 vssd1 vccd1 vccd1 _11299_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_104_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19667_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11379__S1 _09733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13038_ _14557_/A vssd1 vssd1 vccd1 vccd1 _13038_/X sky130_fd_sc_hd__clkbuf_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _12408_/X _17786_/A _17914_/X _12744_/A vssd1 vssd1 vccd1 vccd1 _17915_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_79_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18895_ _19282_/CLK _18895_/D vssd1 vssd1 vccd1 vccd1 _18895_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17846_ _17910_/A _17843_/Y _17845_/Y vssd1 vssd1 vccd1 vccd1 _17846_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10051__S1 _09507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17777_ _17800_/A _17777_/B vssd1 vssd1 vccd1 vccd1 _17777_/Y sky130_fd_sc_hd__nor2_1
X_14989_ _14989_/A vssd1 vssd1 vccd1 vccd1 _18940_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_119_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19866_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_75_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19516_ _19549_/CLK _19516_/D vssd1 vssd1 vccd1 vccd1 _19516_/Q sky130_fd_sc_hd__dfxtp_1
X_16728_ _16731_/B _16731_/C _16718_/X vssd1 vssd1 vccd1 vccd1 _16728_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12098__B _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19447_ _19448_/CLK _19447_/D vssd1 vssd1 vccd1 vccd1 _19447_/Q sky130_fd_sc_hd__dfxtp_1
X_16659_ _16659_/A _16659_/B _16659_/C _16659_/D vssd1 vssd1 vccd1 vccd1 _16669_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_35_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09200_ _19810_/Q _19850_/Q vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__or2b_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09688__A _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19378_ _19378_/CLK _19378_/D vssd1 vssd1 vccd1 vccd1 _19378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11303__S1 _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ _09235_/B _09130_/X input33/X vssd1 vssd1 vccd1 vccd1 _09241_/A sky130_fd_sc_hd__o21ba_2
XANTENNA__16147__A1 _19355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18329_ _19306_/CLK _18329_/D vssd1 vssd1 vccd1 vccd1 _18329_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11730__B _17237_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10627__A _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17895__A1 _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11067__S0 _11127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13381__A1 _13380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13149__S _13172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ _09964_/A _09964_/B vssd1 vssd1 vccd1 vccd1 _09964_/Y sky130_fd_sc_hd__nor2_1
XFILLER_98_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09895_ _09895_/A vssd1 vssd1 vccd1 vccd1 _09895_/Y sky130_fd_sc_hd__inv_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15364__S _15372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12289__A _12289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17799__B _17802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__S1 _09733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11998__A2 _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_14_0_clock_A clkbuf_3_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_83_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19349_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13612__S _13615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09598__A _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _18492_/Q _18987_/Q _10670_/S vssd1 vssd1 vccd1 vccd1 _10670_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _11565_/A _11487_/S _17115_/A _11559_/A vssd1 vssd1 vccd1 vccd1 _11918_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__16923__S _17026_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ _12340_/A _12371_/B vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__nor2_1
XFILLER_127_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_98_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19694_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11058__S0 _11011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14443__S _14443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ _19415_/Q _19416_/Q _12271_/C vssd1 vssd1 vccd1 vccd1 _12293_/B sky130_fd_sc_hd__and3_1
XANTENNA__12752__A _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14010_ _14582_/A vssd1 vssd1 vccd1 vccd1 _14010_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ _18386_/Q _18647_/Q _18546_/Q _18881_/Q _11074_/S _10971_/A vssd1 vssd1 vccd1
+ vccd1 _11222_/X sky130_fd_sc_hd__mux4_1
XFILLER_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _18974_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__12471__B _12471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11922__A2 _12457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _11262_/A _11147_/X _11150_/X _11152_/Y vssd1 vssd1 vccd1 vccd1 _11153_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10281__S1 _10270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ _19321_/Q _18733_/Q _18770_/Q _18344_/Q _10094_/S _10090_/X vssd1 vssd1 vccd1
+ vccd1 _10105_/B sky130_fd_sc_hd__mux4_1
XFILLER_49_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15961_ _15983_/A vssd1 vssd1 vccd1 vccd1 _15970_/S sky130_fd_sc_hd__buf_4
X_11084_ _19174_/Q _18788_/Q _19238_/Q _18357_/Q _10964_/S _11030_/X vssd1 vssd1 vccd1
+ vccd1 _11085_/B sky130_fd_sc_hd__mux4_1
XFILLER_88_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15274__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13583__A _15067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14912_ _14912_/A vssd1 vssd1 vccd1 vccd1 _18902_/D sky130_fd_sc_hd__clkbuf_1
X_17700_ _17700_/A vssd1 vssd1 vccd1 vccd1 _17700_/Y sky130_fd_sc_hd__clkinv_2
X_10035_ _10031_/X _10033_/X _10034_/X _10042_/A _09995_/A vssd1 vssd1 vccd1 vccd1
+ _10040_/B sky130_fd_sc_hd__o221a_1
X_15892_ _19282_/Q _14573_/A _15898_/S vssd1 vssd1 vccd1 vccd1 _15893_/A sky130_fd_sc_hd__mux2_1
X_18680_ _19736_/CLK _18680_/D vssd1 vssd1 vccd1 vccd1 _18680_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_36_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19197_/CLK sky130_fd_sc_hd__clkbuf_16
X_14843_ _18872_/Q _14026_/X _14843_/S vssd1 vssd1 vccd1 vccd1 _14844_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17631_ _17586_/X _17628_/Y _17630_/Y vssd1 vssd1 vccd1 vccd1 _17631_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10894__C1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14624__A1 input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13427__A2 _13380_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14624__B2 _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17562_ _17559_/X _17560_/Y _17744_/S vssd1 vssd1 vccd1 vccd1 _17562_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14774_ _14774_/A vssd1 vssd1 vccd1 vccd1 _18841_/D sky130_fd_sc_hd__clkbuf_1
X_11986_ _11959_/A _11959_/B _11956_/A vssd1 vssd1 vccd1 vccd1 _11987_/B sky130_fd_sc_hd__a21bo_1
X_16513_ _19605_/Q _19604_/Q _19606_/Q _16874_/A vssd1 vssd1 vccd1 vccd1 _16882_/A
+ sky130_fd_sc_hd__and4_1
X_19301_ _19301_/CLK _19301_/D vssd1 vssd1 vccd1 vccd1 _19301_/Q sky130_fd_sc_hd__dfxtp_1
X_13725_ _13090_/X _18431_/Q _13725_/S vssd1 vssd1 vccd1 vccd1 _13726_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17493_ _17490_/X _17487_/Y _17492_/Y vssd1 vssd1 vccd1 vccd1 _17493_/Y sky130_fd_sc_hd__a21oi_1
X_10937_ _10937_/A _10937_/B vssd1 vssd1 vccd1 vccd1 _10937_/X sky130_fd_sc_hd__and2_1
XFILLER_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14618__S _14621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_152_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16444_ _16470_/A _16450_/C vssd1 vssd1 vccd1 vccd1 _16444_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19232_ _19390_/CLK _19232_/D vssd1 vssd1 vccd1 vccd1 _19232_/Q sky130_fd_sc_hd__dfxtp_1
X_13656_ _13107_/X _18400_/Q _13664_/S vssd1 vssd1 vccd1 vccd1 _13657_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10868_ _09617_/A _10846_/X _10866_/X _09578_/A _10867_/Y vssd1 vssd1 vccd1 vccd1
+ _12453_/A sky130_fd_sc_hd__o32a_4
XFILLER_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12938__A1 _19495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ _19630_/Q _12490_/A _12606_/Y _19555_/Q _12584_/Y vssd1 vssd1 vccd1 vccd1
+ _12607_/X sky130_fd_sc_hd__a221o_1
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19163_ _19598_/CLK _19163_/D vssd1 vssd1 vccd1 vccd1 _19163_/Q sky130_fd_sc_hd__dfxtp_1
X_16375_ _19440_/Q _16373_/B _16374_/Y vssd1 vssd1 vccd1 vccd1 _19440_/D sky130_fd_sc_hd__o21a_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13587_ _18375_/Q _13586_/X _13593_/S vssd1 vssd1 vccd1 vccd1 _13588_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10447__A _11445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _18780_/Q vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18114_ _18114_/A _18116_/B vssd1 vssd1 vccd1 vccd1 _18114_/X sky130_fd_sc_hd__or2_1
XFILLER_9_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15326_ _19075_/Q _15009_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15327_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ _13012_/A vssd1 vssd1 vccd1 vccd1 _12538_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19094_ _19290_/CLK _19094_/D vssd1 vssd1 vccd1 vccd1 _19094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15449__S _15455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18045_ _18045_/A vssd1 vssd1 vccd1 vccd1 _19792_/D sky130_fd_sc_hd__clkbuf_1
X_15257_ _15257_/A vssd1 vssd1 vccd1 vccd1 _19044_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12469_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12474_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14208_ _14208_/A vssd1 vssd1 vccd1 vccd1 _18612_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15188_ _15188_/A vssd1 vssd1 vccd1 vccd1 _19013_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14139_ _18582_/Q _13965_/X _14147_/S vssd1 vssd1 vccd1 vccd1 _14140_/A sky130_fd_sc_hd__mux2_1
XFILLER_87_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18947_ _19012_/CLK _18947_/D vssd1 vssd1 vccd1 vccd1 _18947_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_77_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12323__C1 _11686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15184__S _15184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11677__A1 _09665_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09680_ _10451_/S vssd1 vssd1 vccd1 vccd1 _09681_/A sky130_fd_sc_hd__buf_2
XFILLER_39_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10910__A _10910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18878_ _19113_/CLK _18878_/D vssd1 vssd1 vccd1 vccd1 _18878_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11677__B2 _19710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10885__C1 _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17829_ _19729_/Q _17828_/X _17873_/S vssd1 vssd1 vccd1 vccd1 _17830_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15912__S _15920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__B2 _10087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_167_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09114_ _18083_/A _18081_/A _09172_/C vssd1 vssd1 vccd1 vccd1 _17120_/C sky130_fd_sc_hd__nor3_2
XFILLER_149_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_129_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15359__S _15361_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09881__A _10341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ _09941_/A _09944_/X _09946_/X _09740_/A vssd1 vssd1 vccd1 vccd1 _09947_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_77_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09878_ _10214_/A vssd1 vssd1 vccd1 vccd1 _09890_/A sky130_fd_sc_hd__clkbuf_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11127__S _11127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15822__S _15826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11840_/A vssd1 vssd1 vccd1 vccd1 _11949_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13290__A0 _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11770_/Y _11765_/Y _14275_/B vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__mux2_1
XFILLER_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13510_ _14371_/B vssd1 vssd1 vccd1 vccd1 _14860_/B sky130_fd_sc_hd__buf_6
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _19308_/Q _18720_/Q _18757_/Q _18331_/Q _10704_/S _10623_/A vssd1 vssd1 vccd1
+ vccd1 _10722_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14490_/A vssd1 vssd1 vccd1 vccd1 _18729_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12466__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ _13441_/A vssd1 vssd1 vccd1 vccd1 _18321_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11279__S0 _10962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10653_ _10667_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10653_/X sky130_fd_sc_hd__or2_1
XFILLER_70_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16160_ _16159_/A _16159_/C _19769_/Q vssd1 vssd1 vccd1 vccd1 _16161_/B sky130_fd_sc_hd__o21ai_1
XFILLER_155_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _19619_/Q vssd1 vssd1 vccd1 vccd1 _16520_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10584_ _19184_/Q _18798_/Q _19248_/Q _18367_/Q _10576_/X _10577_/X vssd1 vssd1 vccd1
+ vccd1 _10585_/B sky130_fd_sc_hd__mux4_2
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15111_ _15111_/A vssd1 vssd1 vccd1 vccd1 _18979_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_103_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12323_ _12369_/A _12317_/Y _12322_/X _11686_/X vssd1 vssd1 vccd1 vccd1 _12323_/X
+ sky130_fd_sc_hd__a211o_1
X_16091_ _16091_/A _16091_/B _16091_/C vssd1 vssd1 vccd1 vccd1 _16098_/B sky130_fd_sc_hd__or3_1
XANTENNA__12482__A _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14542__A0 _14541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09549__B1 _09485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13345__A1 _13344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15042_ _18957_/Q _15041_/X _15045_/S vssd1 vssd1 vccd1 vccd1 _15043_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12254_ _12253_/X _12252_/Y _12341_/S vssd1 vssd1 vccd1 vccd1 _12254_/X sky130_fd_sc_hd__mux2_1
XFILLER_108_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16889__A _16914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11205_ _19171_/Q _18785_/Q _19235_/Q _18354_/Q _11128_/S _11177_/A vssd1 vssd1 vccd1
+ vccd1 _11206_/B sky130_fd_sc_hd__mux4_2
XFILLER_122_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19850_ _19854_/CLK _19850_/D vssd1 vssd1 vccd1 vccd1 _19850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12185_ _16993_/A _12205_/C _15601_/A vssd1 vssd1 vccd1 vccd1 _12185_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18801_ _19315_/CLK _18801_/D vssd1 vssd1 vccd1 vccd1 _18801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11136_ _10943_/X _11126_/X _11130_/X _11135_/X _11001_/A vssd1 vssd1 vccd1 vccd1
+ _11136_/X sky130_fd_sc_hd__a311o_1
X_19781_ _19786_/CLK _19781_/D vssd1 vssd1 vccd1 vccd1 _19781_/Q sky130_fd_sc_hd__dfxtp_2
X_16993_ _16993_/A _16998_/B vssd1 vssd1 vccd1 vccd1 _16993_/X sky130_fd_sc_hd__or2_1
XFILLER_110_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13517__S _13529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18036__A1 _12126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11826__A _11826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18732_ _19320_/CLK _18732_/D vssd1 vssd1 vccd1 vccd1 _18732_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10006__S1 _09543_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11067_ _19270_/Q _19108_/Q _18517_/Q _18287_/Q _11127_/S _11012_/X vssd1 vssd1 vccd1
+ vccd1 _11067_/X sky130_fd_sc_hd__mux4_1
X_15944_ _13538_/X _19305_/Q _15948_/S vssd1 vssd1 vccd1 vccd1 _15945_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10018_ _10261_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10018_/Y sky130_fd_sc_hd__nand2_1
X_18663_ _19377_/CLK _18663_/D vssd1 vssd1 vccd1 vccd1 _18663_/Q sky130_fd_sc_hd__dfxtp_1
X_15875_ _15875_/A vssd1 vssd1 vccd1 vccd1 _19274_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14826_ _18864_/Q _14001_/X _14832_/S vssd1 vssd1 vccd1 vccd1 _14827_/A sky130_fd_sc_hd__mux2_1
X_17614_ _17461_/A _17512_/X _17613_/X vssd1 vssd1 vccd1 vccd1 _17614_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18594_ _19089_/CLK _18594_/D vssd1 vssd1 vccd1 vccd1 _18594_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10619__C1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14757_ _14579_/X _18834_/Q _14759_/S vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__mux2_1
X_17545_ _17434_/X _17527_/X _17544_/X _17473_/X vssd1 vssd1 vccd1 vccd1 _17545_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14348__S _14354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _19402_/Q _11969_/B _11969_/C _11969_/D vssd1 vssd1 vccd1 vccd1 _12011_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13252__S _13252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ _12924_/X _18423_/Q _13714_/S vssd1 vssd1 vccd1 vccd1 _13709_/A sky130_fd_sc_hd__mux2_1
X_17476_ _19709_/Q _17430_/X _17474_/X _17475_/Y vssd1 vssd1 vccd1 vccd1 _19709_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_60_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14688_ _14688_/A vssd1 vssd1 vccd1 vccd1 _18803_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19215_ _19245_/CLK _19215_/D vssd1 vssd1 vccd1 vccd1 _19215_/Q sky130_fd_sc_hd__dfxtp_1
X_16427_ _16427_/A _16431_/C vssd1 vssd1 vccd1 vccd1 _16427_/Y sky130_fd_sc_hd__nor2_1
X_13639_ _13639_/A vssd1 vssd1 vccd1 vccd1 _18392_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16358_ _16589_/A vssd1 vssd1 vccd1 vccd1 _16546_/A sky130_fd_sc_hd__clkbuf_4
X_19146_ _19356_/CLK _19146_/D vssd1 vssd1 vccd1 vccd1 _19146_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_158_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15309_ _14611_/X _19068_/Q _15311_/S vssd1 vssd1 vccd1 vccd1 _15310_/A sky130_fd_sc_hd__mux2_1
X_16289_ _16289_/A vssd1 vssd1 vccd1 vccd1 _19412_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14083__S _14085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19077_ _19109_/CLK _19077_/D vssd1 vssd1 vccd1 vccd1 _19077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18028_ _18028_/A vssd1 vssd1 vccd1 vccd1 _19785_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15907__S _15909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09801_ _09817_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _09801_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09960__B1 _09909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18027__A1 _19406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11736__A _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09732_ _09732_/A vssd1 vssd1 vccd1 vccd1 _11368_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09663_ _11418_/A _12479_/B _11468_/A vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__a21boi_1
XFILLER_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09594_ _18415_/Q _18676_/Q _18575_/Q _18910_/Q _10603_/S _10669_/A vssd1 vssd1 vccd1
+ vccd1 _09595_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14258__S _14264_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15878__A _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10087__A _10087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12378__A2 _12479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10815__A _18780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_100_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11889__A1 _19401_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11646__A _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13990_ _13990_/A vssd1 vssd1 vccd1 vccd1 _18525_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_105_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _19714_/Q _15499_/B _13103_/S vssd1 vssd1 vccd1 vccd1 _12941_/X sky130_fd_sc_hd__mux2_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _14550_/X _19179_/Q _15660_/S vssd1 vssd1 vccd1 vccd1 _15661_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12872_ _19524_/Q vssd1 vssd1 vccd1 vccd1 _16650_/B sky130_fd_sc_hd__clkbuf_1
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18148__B _18188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14611_ _14611_/A vssd1 vssd1 vccd1 vccd1 _14611_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _11791_/A _11791_/B _11822_/X vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__a21boi_2
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15591_ _15591_/A vssd1 vssd1 vccd1 vccd1 _19160_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09467__C1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17328_/X _17329_/Y _09309_/X _12739_/X vssd1 vssd1 vccd1 vccd1 _19707_/D
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _14541_/X _18753_/Q _14551_/S vssd1 vssd1 vccd1 vccd1 _14543_/A sky130_fd_sc_hd__mux2_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11754_ _19396_/Q _11640_/X _11740_/X _11753_/X vssd1 vssd1 vccd1 vccd1 _16251_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15004__A1 _15003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_25_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12196__B _17810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17261_ _12089_/X _17743_/B _17261_/S vssd1 vssd1 vccd1 vccd1 _17261_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10705_ _10705_/A _10704_/X vssd1 vssd1 vccd1 vccd1 _10705_/X sky130_fd_sc_hd__or2b_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14473_ _14473_/A vssd1 vssd1 vccd1 vccd1 _18721_/D sky130_fd_sc_hd__clkbuf_1
X_11685_ _11734_/A vssd1 vssd1 vccd1 vccd1 _12037_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16212_ _16212_/A vssd1 vssd1 vccd1 vccd1 _19378_/D sky130_fd_sc_hd__clkbuf_1
X_19000_ _19290_/CLK _19000_/D vssd1 vssd1 vccd1 vccd1 _19000_/Q sky130_fd_sc_hd__dfxtp_1
X_13424_ _13423_/X _18319_/Q _13424_/S vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09786__A _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17192_ _17404_/B _17726_/A vssd1 vssd1 vccd1 vccd1 _17471_/B sky130_fd_sc_hd__or2_1
X_10636_ _18924_/Q _18690_/Q _19372_/Q _19020_/Q _10022_/X _10567_/X vssd1 vssd1 vccd1
+ vccd1 _10637_/B sky130_fd_sc_hd__mux4_1
X_16143_ _16142_/A _16142_/C _16142_/B vssd1 vssd1 vccd1 vccd1 _16143_/Y sky130_fd_sc_hd__o21ai_1
X_13355_ _19582_/Q _12606_/Y _12600_/Y _19358_/Q _13354_/X vssd1 vssd1 vccd1 vccd1
+ _13355_/X sky130_fd_sc_hd__a221o_1
XFILLER_6_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10567_ _10586_/A vssd1 vssd1 vccd1 vccd1 _10567_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _17312_/A _17856_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__a21bo_1
XFILLER_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16074_ _16069_/A _16073_/C _13095_/A vssd1 vssd1 vccd1 vccd1 _16075_/B sky130_fd_sc_hd__o21ai_1
X_13286_ _19578_/Q _13055_/X _13285_/X _13265_/X vssd1 vssd1 vccd1 vccd1 _13286_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_142_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10498_ _10509_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10498_/X sky130_fd_sc_hd__or2_1
X_15025_ _15025_/A vssd1 vssd1 vccd1 vccd1 _15025_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12237_ _12232_/X _12236_/X _19414_/Q _11963_/X vssd1 vssd1 vccd1 vccd1 _12237_/X
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_151_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12541__A2 _12507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19833_ _19834_/CLK _19833_/D vssd1 vssd1 vccd1 vccd1 _19833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12168_ _12168_/A _12168_/B vssd1 vssd1 vccd1 vccd1 _12169_/A sky130_fd_sc_hd__or2_1
XFILLER_122_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11119_ _11111_/Y _11114_/Y _11116_/Y _11118_/Y _10929_/A vssd1 vssd1 vccd1 vccd1
+ _11119_/X sky130_fd_sc_hd__o221a_1
XANTENNA__15028__A _15028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19764_ _19793_/CLK _19764_/D vssd1 vssd1 vccd1 vccd1 _19764_/Q sky130_fd_sc_hd__dfxtp_1
X_16976_ _19644_/Q _16984_/B vssd1 vssd1 vccd1 vccd1 _16976_/X sky130_fd_sc_hd__or2_1
X_12099_ _12099_/A _12151_/C vssd1 vssd1 vccd1 vccd1 _12099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15491__A1 _19143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18715_ _19305_/CLK _18715_/D vssd1 vssd1 vccd1 vccd1 _18715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 io_dbus_rdata[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_15927_ _15983_/A vssd1 vssd1 vccd1 vccd1 _15996_/S sky130_fd_sc_hd__clkbuf_8
X_19695_ _19695_/CLK _19695_/D vssd1 vssd1 vccd1 vccd1 _19695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18646_ _19268_/CLK _18646_/D vssd1 vssd1 vccd1 vccd1 _18646_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15858_ _15858_/A vssd1 vssd1 vccd1 vccd1 _19266_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ _14809_/A vssd1 vssd1 vccd1 vccd1 _18856_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_52_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18577_ _19712_/CLK _18577_/D vssd1 vssd1 vccd1 vccd1 _18577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15789_ _13522_/X _19236_/Q _15793_/S vssd1 vssd1 vccd1 vccd1 _15790_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11291__A _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17528_ _17731_/S _17503_/X _17457_/X vssd1 vssd1 vccd1 vccd1 _17684_/A sky130_fd_sc_hd__o21ai_1
XFILLER_51_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09473__A2 _09452_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16743__A1 _19557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17459_ _17392_/X _17715_/A _17402_/X vssd1 vssd1 vccd1 vccd1 _17459_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19129_ _19385_/CLK _19129_/D vssd1 vssd1 vccd1 vccd1 _19129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13309__A1 _12798_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16322__A _16341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__A _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15482__A1 _15481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09715_ _09715_/A vssd1 vssd1 vccd1 vccd1 _09715_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__12296__A1 _19353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15372__S _15372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09646_ _09646_/A vssd1 vssd1 vccd1 vccd1 _09646_/Y sky130_fd_sc_hd__inv_2
XFILLER_83_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__buf_2
XFILLER_55_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16982__A1 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16734__A1 _16736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17931__A0 _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11470_ _11470_/A _11470_/B _11469_/X vssd1 vssd1 vccd1 vccd1 _11470_/X sky130_fd_sc_hd__or3b_1
XFILLER_137_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09847__S0 _09846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10421_ _10237_/X _10420_/X _10243_/X vssd1 vssd1 vccd1 vccd1 _10421_/X sky130_fd_sc_hd__o21a_1
XFILLER_51_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ _13140_/A vssd1 vssd1 vccd1 vccd1 _18300_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_124_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10352_ _09765_/A _10343_/X _10345_/Y _10351_/Y _09813_/A vssd1 vssd1 vccd1 vccd1
+ _10352_/X sky130_fd_sc_hd__o311a_4
XFILLER_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _13070_/X _18296_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__mux2_1
X_10283_ _10335_/A _10276_/X _10282_/X vssd1 vssd1 vccd1 vccd1 _10283_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12022_ _12022_/A vssd1 vssd1 vccd1 vccd1 _12022_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_104_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input49_A io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16830_ _19583_/Q _16830_/B vssd1 vssd1 vccd1 vccd1 _16831_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10280__A _10433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16761_ _19562_/Q _16761_/B vssd1 vssd1 vccd1 vccd1 _16772_/D sky130_fd_sc_hd__and2_1
XANTENNA__13484__A0 _13191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13973_ _18520_/Q _13972_/X _13979_/S vssd1 vssd1 vccd1 vccd1 _13974_/A sky130_fd_sc_hd__mux2_1
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10298__B1 _10297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18500_ _19286_/CLK _18500_/D vssd1 vssd1 vccd1 vccd1 _18500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17063__A _17085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ _14541_/A vssd1 vssd1 vccd1 vccd1 _12924_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_15712_ _15780_/S vssd1 vssd1 vccd1 vccd1 _15721_/S sky130_fd_sc_hd__clkbuf_4
X_16692_ _16697_/C _16697_/D _16675_/X vssd1 vssd1 vccd1 vccd1 _16692_/Y sky130_fd_sc_hd__a21oi_1
X_19480_ _19610_/CLK _19480_/D vssd1 vssd1 vccd1 vccd1 _19480_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10393__S0 _10274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18431_ _19248_/CLK _18431_/D vssd1 vssd1 vccd1 vccd1 _18431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15643_ _14525_/X _19171_/Q _15649_/S vssd1 vssd1 vccd1 vccd1 _15644_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12855_ _13164_/A vssd1 vssd1 vccd1 vccd1 _12855_/X sky130_fd_sc_hd__buf_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11806_ _19636_/Q _13423_/A vssd1 vssd1 vccd1 vccd1 _11806_/Y sky130_fd_sc_hd__nand2_1
X_15574_ _15519_/X _15572_/X _15573_/Y _15549_/X _18271_/Q vssd1 vssd1 vccd1 vccd1
+ _15574_/X sky130_fd_sc_hd__a32o_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _19243_/CLK _18362_/D vssd1 vssd1 vccd1 vccd1 _18362_/Q sky130_fd_sc_hd__dfxtp_1
X_12786_ _18316_/Q _12603_/X _12784_/X _19138_/Q _12785_/X vssd1 vssd1 vccd1 vccd1
+ _12786_/X sky130_fd_sc_hd__a221o_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12000__A _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14525_ _14525_/A vssd1 vssd1 vccd1 vccd1 _14525_/X sky130_fd_sc_hd__clkbuf_1
X_17313_ _17408_/A vssd1 vssd1 vccd1 vccd1 _17462_/A sky130_fd_sc_hd__clkbuf_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11737_/A _11768_/B vssd1 vssd1 vccd1 vccd1 _11737_/Y sky130_fd_sc_hd__nor2_1
X_18293_ _19307_/CLK _18293_/D vssd1 vssd1 vccd1 vccd1 _18293_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10696__S1 _10705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16407__A _16442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13539__A1 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ _13854_/X _18714_/Q _14456_/S vssd1 vssd1 vccd1 vccd1 _14457_/A sky130_fd_sc_hd__mux2_1
X_17244_ _17236_/X _17242_/X _17396_/A vssd1 vssd1 vccd1 vccd1 _17244_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11668_ _17225_/A _11668_/B _17575_/S vssd1 vssd1 vccd1 vccd1 _11669_/B sky130_fd_sc_hd__or3_1
XFILLER_168_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13407_ _13407_/A vssd1 vssd1 vccd1 vccd1 _18316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10619_ _09995_/X _10612_/X _10614_/X _10618_/X _09614_/X vssd1 vssd1 vccd1 vccd1
+ _10619_/X sky130_fd_sc_hd__a311o_4
X_17175_ _17175_/A _17175_/B _17175_/C _17175_/D vssd1 vssd1 vccd1 vccd1 _17176_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_128_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14387_ _13857_/X _18683_/Q _14395_/S vssd1 vssd1 vccd1 vccd1 _14388_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11599_ _19843_/Q _11721_/S _11596_/A _11755_/A vssd1 vssd1 vccd1 vccd1 _11599_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11050__S _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10222__B1 _09765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16126_ _16126_/A _19763_/Q _16126_/C vssd1 vssd1 vccd1 vccd1 _16133_/B sky130_fd_sc_hd__or3_1
X_13338_ _19549_/Q vssd1 vssd1 vccd1 vccd1 _16724_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17150__A1 _09096_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11970__B1 _11969_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15457__S _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13766__A _13822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ _16064_/B _16057_/B vssd1 vssd1 vccd1 vccd1 _16057_/Y sky130_fd_sc_hd__nand2_1
X_13269_ _16904_/A _13260_/X _13261_/X _16493_/A _13268_/X vssd1 vssd1 vccd1 vccd1
+ _15598_/B sky130_fd_sc_hd__a221o_4
XANTENNA__14361__S _14365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15008_ _15008_/A vssd1 vssd1 vccd1 vccd1 _18946_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11317__A3 _11316_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19816_ _19834_/CLK _19816_/D vssd1 vssd1 vccd1 vccd1 _19816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19747_ _19779_/CLK _19747_/D vssd1 vssd1 vccd1 vccd1 _19747_/Q sky130_fd_sc_hd__dfxtp_1
X_16959_ _16959_/A vssd1 vssd1 vccd1 vccd1 _17013_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09500_ _09500_/A vssd1 vssd1 vccd1 vccd1 _10518_/S sky130_fd_sc_hd__clkbuf_4
X_19678_ _19695_/CLK _19678_/D vssd1 vssd1 vccd1 vccd1 _19678_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10384__S0 _10274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09431_ _09431_/A vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__buf_2
X_18629_ _19286_/CLK _18629_/D vssd1 vssd1 vccd1 vccd1 _18629_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16964__A1 _15509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15920__S _15920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__B _14197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09362_ _17120_/B _11569_/A vssd1 vssd1 vccd1 vccd1 _17117_/B sky130_fd_sc_hd__nand2_1
XFILLER_162_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10136__S0 _09846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09293_ _19831_/Q vssd1 vssd1 vccd1 vccd1 _16619_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13440__S _13448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12202__A1 _12200_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_146_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12753__A2 _12752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17141__A1 _18099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput140 _12454_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[9] sky130_fd_sc_hd__buf_2
Xoutput151 _12136_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[18] sky130_fd_sc_hd__buf_2
XFILLER_121_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput162 _12376_/Y vssd1 vssd1 vccd1 vccd1 io_ibus_addr[28] sky130_fd_sc_hd__buf_2
XFILLER_115_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput173 _16262_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[9] sky130_fd_sc_hd__buf_2
XFILLER_115_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10516__A1 _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10611__S1 _09419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16198__S _16202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11924__A _19782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13615__S _13615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10970_ _18642_/Q vssd1 vssd1 vccd1 vccd1 _10971_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ _19328_/Q _18740_/Q _18777_/Q _18351_/Q _10692_/S _09628_/X vssd1 vssd1 vccd1
+ vccd1 _09629_/X sky130_fd_sc_hd__mux4_1
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16955__A1 _15487_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _12677_/A vssd1 vssd1 vccd1 vccd1 _12640_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _19441_/Q _12515_/X _12570_/X vssd1 vssd1 vccd1 vccd1 _12571_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__12755__A _12769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14310_ _13854_/X _18650_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _14311_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13350__S _13350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11522_ _11522_/A _11584_/B _11522_/C vssd1 vssd1 vccd1 vccd1 _11523_/D sky130_fd_sc_hd__or3_1
XFILLER_8_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15290_ _15290_/A vssd1 vssd1 vccd1 vccd1 _19059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12474__B _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14241_ _14241_/A vssd1 vssd1 vccd1 vccd1 _18627_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11453_ _11453_/A _11453_/B _11453_/C vssd1 vssd1 vccd1 vccd1 _11453_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__10275__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10404_ _10404_/A _10404_/B vssd1 vssd1 vccd1 vccd1 _10404_/X sky130_fd_sc_hd__or2_1
XFILLER_171_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14172_ _18597_/Q _14013_/X _14180_/S vssd1 vssd1 vccd1 vccd1 _14173_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11384_ _19738_/Q vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__inv_2
XFILLER_152_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ _15051_/A vssd1 vssd1 vccd1 vccd1 _14573_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13586__A _15070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10335_ _10335_/A _10335_/B vssd1 vssd1 vccd1 vccd1 _10335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18980_ _19012_/CLK _18980_/D vssd1 vssd1 vccd1 vccd1 _18980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13054_/A vssd1 vssd1 vccd1 vccd1 _13054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_97_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _15998_/A _19773_/Q _17935_/S vssd1 vssd1 vccd1 vccd1 _17932_/A sky130_fd_sc_hd__mux2_1
XFILLER_105_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10266_ _10518_/S vssd1 vssd1 vccd1 vccd1 _10481_/S sky130_fd_sc_hd__buf_2
XANTENNA__10507__A1 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output155_A _16290_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12005_ _12005_/A _12005_/B vssd1 vssd1 vccd1 vccd1 _12008_/A sky130_fd_sc_hd__and2_2
XFILLER_39_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17862_ _12291_/Y _17786_/X _17861_/X _17795_/X vssd1 vssd1 vccd1 vccd1 _17862_/X
+ sky130_fd_sc_hd__a211o_1
X_10197_ _10197_/A _10197_/B vssd1 vssd1 vccd1 vccd1 _10197_/X sky130_fd_sc_hd__or2_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19601_ _19603_/CLK _19601_/D vssd1 vssd1 vccd1 vccd1 _19601_/Q sky130_fd_sc_hd__dfxtp_1
X_16813_ _16816_/B _16810_/C _16812_/X vssd1 vssd1 vccd1 vccd1 _16813_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17793_ _17390_/A _17703_/B _17792_/X _17633_/X vssd1 vssd1 vccd1 vccd1 _17793_/X
+ sky130_fd_sc_hd__a211o_1
X_19532_ _19541_/CLK _19532_/D vssd1 vssd1 vccd1 vccd1 _19532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16744_ _16752_/B _16742_/B _16718_/X vssd1 vssd1 vccd1 vccd1 _16744_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13956_ _14528_/A vssd1 vssd1 vccd1 vccd1 _13956_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17199__A1 _12245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12649__B _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19463_ _19607_/CLK _19463_/D vssd1 vssd1 vccd1 vccd1 _19463_/Q sky130_fd_sc_hd__dfxtp_1
X_12907_ _14537_/A vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16675_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16675_/X sky130_fd_sc_hd__clkbuf_2
X_13887_ _13886_/X _18495_/Q _13887_/S vssd1 vssd1 vccd1 vccd1 _13888_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18414_ _19375_/CLK _18414_/D vssd1 vssd1 vccd1 vccd1 _18414_/Q sky130_fd_sc_hd__dfxtp_1
X_12838_ _19140_/Q _12784_/X _12836_/X _12837_/X vssd1 vssd1 vccd1 vccd1 _12838_/X
+ sky130_fd_sc_hd__a211o_1
X_15626_ _19736_/Q _15625_/X _15626_/S vssd1 vssd1 vccd1 vccd1 _15626_/X sky130_fd_sc_hd__mux2_1
XFILLER_62_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19394_ _19699_/CLK _19394_/D vssd1 vssd1 vccd1 vccd1 _19394_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_34_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18345_ _19384_/CLK _18345_/D vssd1 vssd1 vccd1 vccd1 _18345_/Q sky130_fd_sc_hd__dfxtp_1
X_15557_ _15556_/X _19154_/Q _15570_/S vssd1 vssd1 vccd1 vccd1 _15558_/A sky130_fd_sc_hd__mux2_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12769_/A vssd1 vssd1 vccd1 vccd1 _12769_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15041__A _15041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14508_ _14508_/A vssd1 vssd1 vccd1 vccd1 _18737_/D sky130_fd_sc_hd__clkbuf_1
X_15488_ _15488_/A vssd1 vssd1 vccd1 vccd1 _15516_/S sky130_fd_sc_hd__clkbuf_2
X_18276_ _19725_/CLK _18276_/D vssd1 vssd1 vccd1 vccd1 _18276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17227_ _17217_/X _17224_/X _17512_/S vssd1 vssd1 vccd1 vccd1 _17227_/X sky130_fd_sc_hd__mux2_1
Xinput20 io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
Xinput31 io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_2
X_14439_ _13934_/X _18707_/Q _14439_/S vssd1 vssd1 vccd1 vccd1 _14440_/A sky130_fd_sc_hd__mux2_1
Xinput42 io_ibus_inst[17] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 io_ibus_inst[27] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
Xinput64 io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09974__A _10087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17158_ _17158_/A vssd1 vssd1 vccd1 vccd1 _19704_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17123__A1 _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16109_ _16109_/A vssd1 vssd1 vccd1 vccd1 _16109_/X sky130_fd_sc_hd__clkbuf_2
X_17089_ _17089_/A vssd1 vssd1 vccd1 vccd1 _19690_/D sky130_fd_sc_hd__clkbuf_1
X_09980_ _18635_/Q _18970_/Q _09980_/S vssd1 vssd1 vccd1 vccd1 _09980_/X sky130_fd_sc_hd__mux2_1
XFILLER_171_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_143_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11728__B _17252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_147_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12671__A1 _16341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09414_ _10764_/S vssd1 vssd1 vccd1 vccd1 _09415_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_41_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10079__B _12477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09345_ _11620_/A _19842_/Q _17115_/A vssd1 vssd1 vccd1 vccd1 _17127_/A sky130_fd_sc_hd__or3b_1
XFILLER_80_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14266__S _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__A1 _12422_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__A _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09276_ _12697_/A _13356_/B vssd1 vssd1 vccd1 vccd1 _09280_/C sky130_fd_sc_hd__nor2_1
XFILLER_138_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14790__A _14858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12187__B1 _19412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09884__A _10347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10737__A1 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17665__A2 _17662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10823__A _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _11390_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _10120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10051_ _18939_/Q _18705_/Q _19387_/Q _19035_/Q _10017_/S _09507_/A vssd1 vssd1 vccd1
+ vccd1 _10052_/B sky130_fd_sc_hd__mux4_1
XFILLER_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__A1 _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17822__C1 _17466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18090__A2 _12694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17325__B _17432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13810_ _13810_/A vssd1 vssd1 vccd1 vccd1 _18468_/D sky130_fd_sc_hd__clkbuf_1
X_14790_ _14858_/S vssd1 vssd1 vccd1 vccd1 _14799_/S sky130_fd_sc_hd__buf_4
XFILLER_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13741_ _13209_/X _18438_/Q _13747_/S vssd1 vssd1 vccd1 vccd1 _13742_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10953_ _10953_/A _10953_/B vssd1 vssd1 vccd1 vccd1 _10953_/X sky130_fd_sc_hd__or2_1
XANTENNA__16928__A1 _19627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16460_ _16485_/A _16460_/B _16460_/C vssd1 vssd1 vccd1 vccd1 _19470_/D sky130_fd_sc_hd__nor3_1
X_13672_ _13672_/A vssd1 vssd1 vccd1 vccd1 _18407_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10884_ _10889_/A _10879_/X _10882_/X _10883_/X vssd1 vssd1 vccd1 vccd1 _10884_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12623_ _19624_/Q _12620_/X _14518_/B vssd1 vssd1 vccd1 vccd1 _12623_/X sky130_fd_sc_hd__mux2_1
X_15411_ _19113_/Q _15028_/X _15411_/S vssd1 vssd1 vccd1 vccd1 _15412_/A sky130_fd_sc_hd__mux2_1
X_16391_ _19446_/Q _16389_/B _16390_/Y vssd1 vssd1 vccd1 vccd1 _19446_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14176__S _14180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18130_ _18130_/A _18135_/B vssd1 vssd1 vccd1 vccd1 _18130_/X sky130_fd_sc_hd__or2_1
X_15342_ _19082_/Q _15031_/X _15350_/S vssd1 vssd1 vccd1 vccd1 _15343_/A sky130_fd_sc_hd__mux2_1
XFILLER_156_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12554_ _12498_/Y _12550_/X _12553_/X vssd1 vssd1 vccd1 vccd1 _19623_/D sky130_fd_sc_hd__o21a_1
XFILLER_40_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ _11567_/A _11541_/A vssd1 vssd1 vccd1 vccd1 _11721_/S sky130_fd_sc_hd__and2b_2
X_15273_ _15273_/A vssd1 vssd1 vccd1 vccd1 _19051_/D sky130_fd_sc_hd__clkbuf_1
X_18061_ _19800_/Q _12391_/A _18061_/S vssd1 vssd1 vccd1 vccd1 _18062_/A sky130_fd_sc_hd__mux2_1
X_12485_ _17336_/A vssd1 vssd1 vccd1 vccd1 _17356_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__14904__S _14904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18172__A _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17012_ _15608_/X _17010_/X _17011_/X _17008_/X vssd1 vssd1 vccd1 vccd1 _19657_/D
+ sky130_fd_sc_hd__o211a_1
X_14224_ _14224_/A vssd1 vssd1 vccd1 vccd1 _18619_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11436_ _11439_/A _11441_/A _11439_/C _10304_/A vssd1 vssd1 vccd1 vccd1 _11436_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_172_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11076__S1 _11033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13390__A2 _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14155_ _14155_/A vssd1 vssd1 vccd1 vccd1 _18589_/D sky130_fd_sc_hd__clkbuf_1
X_11367_ _18480_/Q _19071_/Q _19233_/Q _18448_/Q _09704_/X _09733_/X vssd1 vssd1 vccd1
+ vccd1 _11368_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13106_ _15047_/A vssd1 vssd1 vccd1 vccd1 _14569_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10318_ _10314_/X _10316_/X _10317_/X _10200_/A _09728_/A vssd1 vssd1 vccd1 vccd1
+ _10318_/X sky130_fd_sc_hd__o221a_1
XFILLER_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18963_ _18964_/CLK _18963_/D vssd1 vssd1 vccd1 vccd1 _18963_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14086_ _14086_/A vssd1 vssd1 vccd1 vccd1 _18559_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _11298_/A _11298_/B vssd1 vssd1 vccd1 vccd1 _11298_/X sky130_fd_sc_hd__and2_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15735__S _15743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _17852_/X _17403_/Y _17860_/X _17913_/Y vssd1 vssd1 vccd1 vccd1 _17914_/X
+ sky130_fd_sc_hd__o211a_1
X_13037_ _15035_/A vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__clkbuf_2
X_10249_ _10361_/A _10249_/B vssd1 vssd1 vccd1 vccd1 _10249_/X sky130_fd_sc_hd__or2_1
XFILLER_26_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18894_ _18894_/CLK _18894_/D vssd1 vssd1 vccd1 vccd1 _18894_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10587__S0 _10566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17845_ _17845_/A _17845_/B vssd1 vssd1 vccd1 vccd1 _17845_/Y sky130_fd_sc_hd__nor2_1
XFILLER_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17776_ _17779_/A _17779_/B vssd1 vssd1 vccd1 vccd1 _17777_/B sky130_fd_sc_hd__and2_1
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14988_ _18940_/Q vssd1 vssd1 vccd1 vccd1 _14989_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19515_ _19549_/CLK _19515_/D vssd1 vssd1 vccd1 vccd1 _19515_/Q sky130_fd_sc_hd__dfxtp_1
X_16727_ _19551_/Q _16750_/B _16726_/Y vssd1 vssd1 vccd1 vccd1 _19551_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13939_ _13939_/A vssd1 vssd1 vccd1 vccd1 _18511_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19446_ _19448_/CLK _19446_/D vssd1 vssd1 vccd1 vccd1 _19446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16658_ _19529_/Q _19528_/Q vssd1 vssd1 vccd1 vccd1 _16659_/D sky130_fd_sc_hd__and2_1
XFILLER_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15609_ _19733_/Q _15608_/X _15626_/S vssd1 vssd1 vccd1 vccd1 _15609_/X sky130_fd_sc_hd__mux2_1
X_19377_ _19377_/CLK _19377_/D vssd1 vssd1 vccd1 vccd1 _19377_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16589_ _16589_/A vssd1 vssd1 vccd1 vccd1 _16812_/A sky130_fd_sc_hd__buf_2
XFILLER_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11503__S _11539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09130_ _19706_/Q _19705_/Q vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__or2_1
X_18328_ _19241_/CLK _18328_/D vssd1 vssd1 vccd1 vccd1 _18328_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18259_ _19720_/CLK _18259_/D vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_2
XFILLER_129_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11067__S1 _11012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _18894_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_143_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09963_ _19194_/Q _18808_/Q _19258_/Q _18377_/Q _10168_/S _09773_/A vssd1 vssd1 vccd1
+ vccd1 _09964_/B sky130_fd_sc_hd__mux4_1
XFILLER_116_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15645__S _15649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__A2 _19724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09894_ _18506_/Q _19001_/Q _10166_/S vssd1 vssd1 vccd1 vccd1 _09895_/A sky130_fd_sc_hd__mux2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11144__A1 _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10578__S0 _10576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11695__A2 _19584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__C1 _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16083__A1 _19344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ _09328_/A vssd1 vssd1 vccd1 vccd1 _11559_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10958__A1 _09432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _12494_/A _12522_/A _11803_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _12605_/B
+ sky130_fd_sc_hd__or4b_1
XANTENNA__14724__S _14726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12270_ _19415_/Q _12271_/C _19416_/Q vssd1 vssd1 vccd1 vccd1 _12270_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11058__S1 _11005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11221_ _11075_/A _11218_/Y _11220_/Y _10968_/A vssd1 vssd1 vccd1 vccd1 _11221_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11649__A _19394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11383__B2 _19738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _11072_/A _11151_/X _09531_/A vssd1 vssd1 vccd1 vccd1 _11152_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_150_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10103_ _11380_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _10103_/X sky130_fd_sc_hd__or2_1
XFILLER_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15960_ _15960_/A vssd1 vssd1 vccd1 vccd1 _19312_/D sky130_fd_sc_hd__clkbuf_1
X_11083_ _10915_/X _11078_/X _11080_/Y _11082_/Y _09553_/A vssd1 vssd1 vccd1 vccd1
+ _11083_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11135__A1 _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input31_A io_dbus_rdata[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ _18902_/Q _14020_/X _14915_/S vssd1 vssd1 vccd1 vccd1 _14912_/A sky130_fd_sc_hd__mux2_1
X_10034_ _18939_/Q _18705_/Q _19387_/Q _19035_/Q _09415_/A _09443_/X vssd1 vssd1 vccd1
+ vccd1 _10034_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10343__C1 _10378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15891_ _15891_/A vssd1 vssd1 vccd1 vccd1 _19281_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17271__A0 _17819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11384__A _19738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17630_ _17630_/A _17630_/B vssd1 vssd1 vccd1 vccd1 _17630_/Y sky130_fd_sc_hd__nor2_1
X_14842_ _14842_/A vssd1 vssd1 vccd1 vccd1 _18871_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14085__A0 _13886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17561_ _17584_/A vssd1 vssd1 vccd1 vccd1 _17744_/S sky130_fd_sc_hd__buf_2
X_11985_ _11985_/A _11985_/B vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__nor2_1
X_14773_ _14601_/X _18841_/Q _14781_/S vssd1 vssd1 vccd1 vccd1 _14774_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13803__S _13809_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19300_ _19300_/CLK _19300_/D vssd1 vssd1 vccd1 vccd1 _19300_/Q sky130_fd_sc_hd__dfxtp_1
X_16512_ _19601_/Q _19603_/Q _19602_/Q _16865_/A vssd1 vssd1 vccd1 vccd1 _16874_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__09789__A _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13724_ _13724_/A vssd1 vssd1 vccd1 vccd1 _18430_/D sky130_fd_sc_hd__clkbuf_1
X_10936_ _18615_/Q _18950_/Q _11196_/S vssd1 vssd1 vccd1 vccd1 _10937_/B sky130_fd_sc_hd__mux2_1
XFILLER_72_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17492_ _17716_/S _17492_/B vssd1 vssd1 vccd1 vccd1 _17492_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19231_ _19375_/CLK _19231_/D vssd1 vssd1 vccd1 vccd1 _19231_/Q sky130_fd_sc_hd__dfxtp_1
X_16443_ _16443_/A vssd1 vssd1 vccd1 vccd1 _16450_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_13655_ _13677_/A vssd1 vssd1 vccd1 vccd1 _13664_/S sky130_fd_sc_hd__clkbuf_8
X_10867_ _19715_/Q vssd1 vssd1 vccd1 vccd1 _10867_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10728__A _10769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12606_ _12606_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _12606_/Y sky130_fd_sc_hd__nor2_2
X_19162_ _19162_/CLK _19162_/D vssd1 vssd1 vccd1 vccd1 _19162_/Q sky130_fd_sc_hd__dfxtp_2
X_16374_ _16390_/A _16379_/C vssd1 vssd1 vccd1 vccd1 _16374_/Y sky130_fd_sc_hd__nor2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ _15070_/A vssd1 vssd1 vccd1 vccd1 _13586_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16129__A2 _12715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ _10798_/A _12454_/A vssd1 vssd1 vccd1 vccd1 _11462_/B sky130_fd_sc_hd__nand2_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10447__B _12465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18113_ _19820_/Q _18106_/X _18112_/X _18110_/X vssd1 vssd1 vccd1 vccd1 _19820_/D
+ sky130_fd_sc_hd__o211a_1
X_12537_ _13265_/A vssd1 vssd1 vccd1 vccd1 _13012_/A sky130_fd_sc_hd__clkbuf_2
X_15325_ _15325_/A vssd1 vssd1 vccd1 vccd1 _19074_/D sky130_fd_sc_hd__clkbuf_1
X_19093_ _19223_/CLK _19093_/D vssd1 vssd1 vccd1 vccd1 _19093_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18044_ _19792_/Q _19413_/Q _18050_/S vssd1 vssd1 vccd1 vccd1 _18045_/A sky130_fd_sc_hd__mux2_1
X_15256_ _14534_/X _19044_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15257_/A sky130_fd_sc_hd__mux2_1
X_12468_ _12468_/A _12468_/B vssd1 vssd1 vccd1 vccd1 _12468_/Y sky130_fd_sc_hd__nor2_1
XFILLER_172_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14207_ _18612_/Q _13959_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14208_/A sky130_fd_sc_hd__mux2_1
X_11419_ _11417_/Y _11361_/A _11361_/B _11414_/Y _11418_/Y vssd1 vssd1 vccd1 vccd1
+ _11419_/X sky130_fd_sc_hd__a311o_1
X_15187_ _19013_/Q _15015_/X _15195_/S vssd1 vssd1 vccd1 vccd1 _15188_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12399_ _12301_/X _12480_/B _12398_/Y vssd1 vssd1 vccd1 vccd1 _17907_/B sky130_fd_sc_hd__o21ai_4
XFILLER_113_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14138_ _14195_/S vssd1 vssd1 vccd1 vccd1 _14147_/S sky130_fd_sc_hd__buf_2
XFILLER_99_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14069_ _14069_/A vssd1 vssd1 vccd1 vccd1 _18551_/D sky130_fd_sc_hd__clkbuf_1
X_18946_ _19734_/CLK _18946_/D vssd1 vssd1 vccd1 vccd1 _18946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18877_ _19389_/CLK _18877_/D vssd1 vssd1 vccd1 vccd1 _18877_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12874__B2 _19332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17828_ _17592_/A _17826_/Y _17827_/X _17518_/X _12225_/B vssd1 vssd1 vccd1 vccd1
+ _17828_/X sky130_fd_sc_hd__a32o_1
XFILLER_27_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10980__S0 _10862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17759_ _17532_/X _17739_/X _17758_/X vssd1 vssd1 vccd1 vccd1 _17759_/X sky130_fd_sc_hd__o21ba_1
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09699__A _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19429_ _19436_/CLK _19429_/D vssd1 vssd1 vccd1 vccd1 _19429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09113_ _09113_/A vssd1 vssd1 vccd1 vccd1 _09172_/C sky130_fd_sc_hd__buf_2
XANTENNA__11062__B1 _11007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11601__A2 _12443_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12572__B _13132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_150_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19203_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15375__S _15383_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09946_ _10184_/A _09946_/B vssd1 vssd1 vccd1 vccd1 _09946_/X sky130_fd_sc_hd__or2_1
XFILLER_58_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_165_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _18917_/CLK sky130_fd_sc_hd__clkbuf_16
X_09877_ _09667_/X _09859_/X _09876_/X _09758_/X _19732_/Q vssd1 vssd1 vccd1 vccd1
+ _09975_/A sky130_fd_sc_hd__a32o_4
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16995__A _18097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__B1 _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12617__A1 _18254_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13623__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _11770_/A _12098_/C vssd1 vssd1 vccd1 vccd1 _11770_/Y sky130_fd_sc_hd__nor2_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13290__A1 _15606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10721_/A _10721_/B vssd1 vssd1 vccd1 vccd1 _10721_/Y sky130_fd_sc_hd__nor2_1
XFILLER_53_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13440_ _12801_/X _18321_/Q _13448_/S vssd1 vssd1 vccd1 vccd1 _13441_/A sky130_fd_sc_hd__mux2_1
X_10652_ _19181_/Q _18795_/Q _19245_/Q _18364_/Q _10650_/X _11298_/A vssd1 vssd1 vccd1
+ vccd1 _10653_/B sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_103_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19668_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11279__S1 _11220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13371_ _19770_/Q _13370_/B _12942_/S vssd1 vssd1 vccd1 vccd1 _13371_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14454__S _14456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ _10074_/X _10569_/Y _10574_/X _10582_/Y _09811_/A vssd1 vssd1 vccd1 vccd1
+ _10583_/X sky130_fd_sc_hd__o311a_4
XFILLER_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15110_ _18979_/Q _15009_/X _15112_/S vssd1 vssd1 vccd1 vccd1 _15111_/A sky130_fd_sc_hd__mux2_1
X_12322_ _12322_/A _12322_/B _12322_/C _12322_/D vssd1 vssd1 vccd1 vccd1 _12322_/X
+ sky130_fd_sc_hd__and4_1
X_16090_ _16090_/A vssd1 vssd1 vccd1 vccd1 _19345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12482__B _12482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15041_ _15041_/A vssd1 vssd1 vccd1 vccd1 _15041_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09549__A1 _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12253_ _19415_/Q _12271_/C vssd1 vssd1 vccd1 vccd1 _12253_/X sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_118_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19846_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11204_ _11007_/X _11195_/X _11199_/X _11203_/X _11001_/A vssd1 vssd1 vccd1 vccd1
+ _11204_/X sky130_fd_sc_hd__a311o_1
XFILLER_123_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12184_ _12184_/A vssd1 vssd1 vccd1 vccd1 _15601_/A sky130_fd_sc_hd__buf_2
XFILLER_107_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10564__C1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15285__S _15289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18800_ _19250_/CLK _18800_/D vssd1 vssd1 vccd1 vccd1 _18800_/Q sky130_fd_sc_hd__dfxtp_1
X_11135_ _10807_/A _11131_/X _11133_/X _11134_/X vssd1 vssd1 vccd1 vccd1 _11135_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_21_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19780_ _19780_/CLK _19780_/D vssd1 vssd1 vccd1 vccd1 _19780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16992_ _15568_/X _16983_/X _16991_/X _16981_/X vssd1 vssd1 vccd1 vccd1 _19650_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11108__A1 _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18731_ _19319_/CLK _18731_/D vssd1 vssd1 vccd1 vccd1 _18731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15943_ _15943_/A vssd1 vssd1 vccd1 vccd1 _19304_/D sky130_fd_sc_hd__clkbuf_1
X_11066_ _11128_/S vssd1 vssd1 vccd1 vccd1 _11127_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__11826__B _19399_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11318__S _11318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _18635_/Q _18970_/Q _10017_/S vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__mux2_1
X_18662_ _19282_/CLK _18662_/D vssd1 vssd1 vccd1 vccd1 _18662_/Q sky130_fd_sc_hd__dfxtp_1
X_15874_ _19274_/Q _14547_/A _15876_/S vssd1 vssd1 vccd1 vccd1 _15875_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17613_ _17613_/A _17613_/B vssd1 vssd1 vccd1 vccd1 _17613_/X sky130_fd_sc_hd__or2_1
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14825_ _14825_/A vssd1 vssd1 vccd1 vccd1 _18863_/D sky130_fd_sc_hd__clkbuf_1
X_18593_ _19088_/CLK _18593_/D vssd1 vssd1 vccd1 vccd1 _18593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13533__S _13545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17544_ _17390_/X _17529_/Y _17543_/X vssd1 vssd1 vccd1 vccd1 _17544_/X sky130_fd_sc_hd__a21o_1
X_14756_ _14756_/A vssd1 vssd1 vccd1 vccd1 _18833_/D sky130_fd_sc_hd__clkbuf_1
X_11968_ _12392_/S _11968_/B vssd1 vssd1 vccd1 vccd1 _11968_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17547__A1 _19711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10095__A1 _10138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13707_ _13707_/A vssd1 vssd1 vccd1 vccd1 _18422_/D sky130_fd_sc_hd__clkbuf_1
X_17475_ _11639_/A _17328_/B _09322_/X vssd1 vssd1 vccd1 vccd1 _17475_/Y sky130_fd_sc_hd__o21ai_1
X_10919_ _10977_/A _10919_/B vssd1 vssd1 vccd1 vccd1 _10919_/Y sky130_fd_sc_hd__nor2_1
X_14687_ _14582_/X _18803_/Q _14687_/S vssd1 vssd1 vccd1 vccd1 _14688_/A sky130_fd_sc_hd__mux2_1
X_11899_ _11899_/A _17205_/A vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__or2_1
XFILLER_149_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19214_ _19248_/CLK _19214_/D vssd1 vssd1 vccd1 vccd1 _19214_/Q sky130_fd_sc_hd__dfxtp_1
X_16426_ _16426_/A vssd1 vssd1 vccd1 vccd1 _16431_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13638_ _12945_/X _18392_/Q _13642_/S vssd1 vssd1 vccd1 vccd1 _13639_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19145_ _19796_/CLK _19145_/D vssd1 vssd1 vccd1 vccd1 _19145_/Q sky130_fd_sc_hd__dfxtp_1
X_16357_ _19434_/Q _16352_/C _16356_/Y vssd1 vssd1 vccd1 vccd1 _19434_/D sky130_fd_sc_hd__o21a_1
XFILLER_146_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13569_ _13569_/A vssd1 vssd1 vccd1 vccd1 _18369_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12792__A0 _09309_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15308_ _15308_/A vssd1 vssd1 vccd1 vccd1 _19067_/D sky130_fd_sc_hd__clkbuf_1
X_19076_ _19076_/CLK _19076_/D vssd1 vssd1 vccd1 vccd1 _19076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16288_ _16298_/A _16288_/B vssd1 vssd1 vccd1 vccd1 _16289_/A sky130_fd_sc_hd__and2_1
XFILLER_161_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15730__A0 _13541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18027_ _19785_/Q _19406_/Q _18027_/S vssd1 vssd1 vccd1 vccd1 _18028_/A sky130_fd_sc_hd__mux2_1
X_15239_ _19037_/Q _15092_/X _15239_/S vssd1 vssd1 vccd1 vccd1 _15240_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09982__A _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10555__C1 _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09800_ _18940_/Q _18706_/Q _19388_/Q _19036_/Q _11385_/S _09799_/X vssd1 vssd1 vccd1
+ vccd1 _09801_/B sky130_fd_sc_hd__mux4_1
XFILLER_141_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_82_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19598_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10921__A _11024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18929_ _19315_/CLK _18929_/D vssd1 vssd1 vccd1 vccd1 _18929_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11736__B _19396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09731_ _09687_/X _09697_/X _09716_/X _11373_/A _09730_/X vssd1 vssd1 vccd1 vccd1
+ _09742_/B sky130_fd_sc_hd__o221a_1
XANTENNA__13009__A _13009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09662_ _11413_/A _12480_/B vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_97_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19436_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09593_ _09717_/A _09586_/X _09589_/X _09592_/X vssd1 vssd1 vccd1 vccd1 _09593_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_43_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12848__A _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_clock clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19006_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10087__B _12473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12583__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_35_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19119_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10794__C1 _09658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15721__A0 _13528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_195_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09929_ _10197_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _09929_/X sky130_fd_sc_hd__or2_1
XFILLER_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15833__S _15837_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12940_ _16854_/A _12560_/X _12562_/X _16440_/A _12939_/X vssd1 vssd1 vccd1 vccd1
+ _15499_/B sky130_fd_sc_hd__a221o_2
XFILLER_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _19460_/Q vssd1 vssd1 vccd1 vccd1 _16431_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14610_ _14610_/A vssd1 vssd1 vccd1 vccd1 _18774_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11822_ _11822_/A _17247_/A vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__or2b_1
X_15590_ _15589_/X _19160_/Q _15596_/S vssd1 vssd1 vccd1 vccd1 _15591_/A sky130_fd_sc_hd__mux2_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12477__B _12477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ _16162_/S _11752_/X _11623_/X vssd1 vssd1 vccd1 vccd1 _11753_/X sky130_fd_sc_hd__a21o_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14541_/A vssd1 vssd1 vccd1 vccd1 _14541_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10704_ _18491_/Q _18986_/Q _10704_/S vssd1 vssd1 vccd1 vccd1 _10704_/X sky130_fd_sc_hd__mux2_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ _17215_/X _17722_/B _17261_/S vssd1 vssd1 vccd1 vccd1 _17260_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11684_ _18127_/A _18125_/A _11684_/C _11684_/D vssd1 vssd1 vccd1 vccd1 _11734_/A
+ sky130_fd_sc_hd__nor4_2
X_14472_ _13877_/X _18721_/Q _14478_/S vssd1 vssd1 vccd1 vccd1 _14473_/A sky130_fd_sc_hd__mux2_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ _13573_/X _19378_/Q _16213_/S vssd1 vssd1 vccd1 vccd1 _16212_/A sky130_fd_sc_hd__mux2_1
X_13423_ _13423_/A _13423_/B vssd1 vssd1 vccd1 vccd1 _13423_/X sky130_fd_sc_hd__or2_1
XFILLER_139_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13589__A _15073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10635_ _09543_/A _10632_/Y _10634_/Y _11331_/A vssd1 vssd1 vccd1 vccd1 _10635_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_139_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17191_ _17415_/A vssd1 vssd1 vccd1 vccd1 _17726_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12774__B1 _11416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13354_ _19694_/Q _17028_/A vssd1 vssd1 vccd1 vccd1 _13354_/X sky130_fd_sc_hd__and2_1
X_16142_ _16142_/A _16142_/B _16142_/C vssd1 vssd1 vccd1 vccd1 _16150_/B sky130_fd_sc_hd__or3_1
XFILLER_139_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10566_ _10704_/S vssd1 vssd1 vccd1 vccd1 _10566_/X sky130_fd_sc_hd__buf_4
XFILLER_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _12305_/A vssd1 vssd1 vccd1 vccd1 _17312_/A sky130_fd_sc_hd__clkbuf_2
X_13285_ _19164_/Q _13007_/X _12532_/X _19354_/Q _13284_/X vssd1 vssd1 vccd1 vccd1
+ _13285_/X sky130_fd_sc_hd__a221o_2
XFILLER_115_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16073_ _19753_/Q _19754_/Q _16073_/C vssd1 vssd1 vccd1 vccd1 _16080_/B sky130_fd_sc_hd__or3_1
X_10497_ _18927_/Q _18693_/Q _19375_/Q _19023_/Q _10496_/X _09672_/A vssd1 vssd1 vccd1
+ vccd1 _10498_/B sky130_fd_sc_hd__mux4_1
X_12236_ _12233_/X _12234_/Y _12235_/X _16278_/A vssd1 vssd1 vccd1 vccd1 _12236_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15024_ _15024_/A vssd1 vssd1 vccd1 vccd1 _18951_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19832_ _19834_/CLK _19832_/D vssd1 vssd1 vccd1 vccd1 _19832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12167_ _12167_/A _17202_/A vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__nor2_1
XFILLER_110_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11118_ _11278_/A _11117_/X _09481_/A vssd1 vssd1 vccd1 vccd1 _11118_/Y sky130_fd_sc_hd__o21ai_1
X_19763_ _19793_/CLK _19763_/D vssd1 vssd1 vccd1 vccd1 _19763_/Q sky130_fd_sc_hd__dfxtp_1
X_16975_ _12669_/X _16970_/X _16974_/X _16968_/X vssd1 vssd1 vccd1 vccd1 _19643_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12098_ _19408_/Q _19409_/Q _12098_/C _12098_/D vssd1 vssd1 vccd1 vccd1 _12151_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_77_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18714_ _19302_/CLK _18714_/D vssd1 vssd1 vccd1 vccd1 _18714_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15743__S _15743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15926_ _15926_/A _15926_/B vssd1 vssd1 vccd1 vccd1 _15983_/A sky130_fd_sc_hd__nand2_4
X_11049_ _18613_/Q _18948_/Q _11049_/S vssd1 vssd1 vccd1 vccd1 _11049_/X sky130_fd_sc_hd__mux2_1
X_19694_ _19694_/CLK _19694_/D vssd1 vssd1 vccd1 vccd1 _19694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_2
XFILLER_76_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18645_ _19711_/CLK _18645_/D vssd1 vssd1 vccd1 vccd1 _18645_/Q sky130_fd_sc_hd__dfxtp_1
X_15857_ _19266_/Q _14519_/A _15865_/S vssd1 vssd1 vccd1 vccd1 _15858_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14359__S _14365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15044__A _15044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14808_ _18856_/Q _13975_/X _14810_/S vssd1 vssd1 vccd1 vccd1 _14809_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18576_ _19388_/CLK _18576_/D vssd1 vssd1 vccd1 vccd1 _18576_/Q sky130_fd_sc_hd__dfxtp_1
X_15788_ _15788_/A vssd1 vssd1 vccd1 vccd1 _19235_/D sky130_fd_sc_hd__clkbuf_1
X_17527_ _17674_/A _17526_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17527_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11291__B _12453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14739_ _14785_/S vssd1 vssd1 vccd1 vccd1 _14748_/S sky130_fd_sc_hd__buf_2
XFILLER_44_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09473__A3 _09467_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09977__A _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17458_ _17738_/S _17456_/X _17457_/X vssd1 vssd1 vccd1 vccd1 _17715_/A sky130_fd_sc_hd__o21ai_1
XFILLER_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16409_ _16427_/A _16409_/B vssd1 vssd1 vccd1 vccd1 _16409_/Y sky130_fd_sc_hd__nor2_1
XFILLER_119_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14094__S _14096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17389_ _17597_/A vssd1 vssd1 vccd1 vccd1 _17390_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12765__B1 _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19128_ _19290_/CLK _19128_/D vssd1 vssd1 vccd1 vccd1 _19128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_119_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15918__S _15920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19059_ _19379_/CLK _19059_/D vssd1 vssd1 vccd1 vccd1 _19059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09933__A1 _09733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11740__A1 _19332_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11179__S0 _11243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09714_ _09714_/A vssd1 vssd1 vccd1 vccd1 _09715_/A sky130_fd_sc_hd__buf_2
XFILLER_28_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17759__A1 _17532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09645_ _18511_/Q _19006_/Q _09645_/S vssd1 vssd1 vccd1 vccd1 _09646_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09576_/A vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12048__A2 _12464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__S0 _10479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15889__A _15911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09887__A _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11008__B1 _11007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15942__A0 _13535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11103__S0 _09624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ _18594_/Q _18865_/Q _19089_/Q _18833_/Q _10368_/S _09674_/A vssd1 vssd1 vccd1
+ vccd1 _10420_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12756__B1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10351_ _10345_/A _10346_/X _10350_/X vssd1 vssd1 vccd1 vccd1 _10351_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_100_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13070_ _14563_/A vssd1 vssd1 vccd1 vccd1 _13070_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_151_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10282_ _10429_/A _10281_/X _09764_/A vssd1 vssd1 vccd1 vccd1 _10282_/X sky130_fd_sc_hd__o21a_1
XFILLER_124_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17328__B _17328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12021_ _12021_/A vssd1 vssd1 vccd1 vccd1 _12021_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11657__A _19628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09127__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16760_ _19561_/Q _16760_/B _16760_/C vssd1 vssd1 vccd1 vccd1 _16761_/B sky130_fd_sc_hd__and3_1
XFILLER_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13972_ _14544_/A vssd1 vssd1 vccd1 vccd1 _13972_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_101_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10298__A1 _10378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15711_ _15767_/A vssd1 vssd1 vccd1 vccd1 _15780_/S sky130_fd_sc_hd__buf_6
X_12923_ _15019_/A vssd1 vssd1 vccd1 vccd1 _14541_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16691_ _19539_/Q _16695_/D _16690_/Y vssd1 vssd1 vccd1 vccd1 _19539_/D sky130_fd_sc_hd__o21a_1
XFILLER_100_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12488__A _17317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10393__S1 _10275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18430_ _19309_/CLK _18430_/D vssd1 vssd1 vccd1 vccd1 _18430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15642_ _15642_/A vssd1 vssd1 vccd1 vccd1 _19170_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12854_ _18744_/Q vssd1 vssd1 vccd1 vccd1 _13164_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11805_ _16937_/A _13430_/A _11805_/C _11805_/D vssd1 vssd1 vccd1 vccd1 _13423_/A
+ sky130_fd_sc_hd__and4bb_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18361_ _19243_/CLK _18361_/D vssd1 vssd1 vccd1 vccd1 _18361_/Q sky130_fd_sc_hd__dfxtp_1
X_15573_ _15607_/A _18271_/Q vssd1 vssd1 vccd1 vccd1 _15573_/Y sky130_fd_sc_hd__nand2_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output100_A _11824_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _19664_/Q _12703_/X _12704_/X _19631_/Q vssd1 vssd1 vccd1 vccd1 _12785_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18175__B2 _18087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11798__A1 _19334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17312_ _17312_/A _17319_/B _17404_/C vssd1 vssd1 vccd1 vccd1 _17408_/A sky130_fd_sc_hd__or3_1
XFILLER_25_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14524_ _14524_/A vssd1 vssd1 vccd1 vccd1 _18747_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18292_ _19308_/CLK _18292_/D vssd1 vssd1 vccd1 vccd1 _18292_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _19395_/Q _19396_/Q _11736_/C vssd1 vssd1 vccd1 vccd1 _11768_/B sky130_fd_sc_hd__and3_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15933__A0 _13522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17243_ _17438_/S vssd1 vssd1 vccd1 vccd1 _17396_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14455_ _14455_/A vssd1 vssd1 vccd1 vccd1 _18713_/D sky130_fd_sc_hd__clkbuf_1
X_11667_ _19394_/Q _11640_/X _11656_/Y _11666_/Y vssd1 vssd1 vccd1 vccd1 _16247_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_128_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13406_ _13405_/X _18316_/Q _13424_/S vssd1 vssd1 vccd1 vccd1 _13407_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10618_ _10559_/A _10615_/X _10617_/X _09450_/A vssd1 vssd1 vccd1 vccd1 _10618_/X
+ sky130_fd_sc_hd__o211a_1
X_17174_ _17174_/A _17174_/B vssd1 vssd1 vccd1 vccd1 _17176_/C sky130_fd_sc_hd__or2_1
X_14386_ _14443_/S vssd1 vssd1 vccd1 vccd1 _14395_/S sky130_fd_sc_hd__buf_2
XANTENNA__12211__A2 _12471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ _09331_/A _09194_/X _12730_/C vssd1 vssd1 vccd1 vccd1 _11598_/X sky130_fd_sc_hd__mux2_1
XFILLER_155_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16125_ _16125_/A vssd1 vssd1 vccd1 vccd1 _19351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10549_ _10310_/A _10545_/X _10548_/X vssd1 vssd1 vccd1 vccd1 _10549_/X sky130_fd_sc_hd__a21o_1
X_13337_ _13335_/Y _13362_/B _11499_/X vssd1 vssd1 vccd1 vccd1 _13337_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_115_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11970__A1 _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16056_ _16055_/A _16055_/C _16055_/B vssd1 vssd1 vccd1 vccd1 _16057_/B sky130_fd_sc_hd__o21ai_1
X_13268_ _19545_/Q _13004_/X _13054_/X _19513_/Q _13267_/X vssd1 vssd1 vccd1 vccd1
+ _13268_/X sky130_fd_sc_hd__a221o_1
XFILLER_170_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15007_ _18946_/Q _15006_/X _15013_/S vssd1 vssd1 vccd1 vccd1 _15008_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12219_ _12219_/A vssd1 vssd1 vccd1 vccd1 _17819_/B sky130_fd_sc_hd__buf_2
X_13199_ _19159_/Q _13179_/X _12958_/X _19349_/Q _13198_/X vssd1 vssd1 vccd1 vccd1
+ _13199_/X sky130_fd_sc_hd__a221o_2
XFILLER_97_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19815_ _19834_/CLK _19815_/D vssd1 vssd1 vccd1 vccd1 _19815_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_110_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16958_ _15495_/X _16956_/X _16957_/X _16954_/X vssd1 vssd1 vccd1 vccd1 _19637_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_56_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19746_ _19780_/CLK _19746_/D vssd1 vssd1 vccd1 vccd1 _19746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15909_ _19290_/Q _14598_/A _15909_/S vssd1 vssd1 vccd1 vccd1 _15910_/A sky130_fd_sc_hd__mux2_1
X_19677_ _19687_/CLK _19677_/D vssd1 vssd1 vccd1 vccd1 _19677_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16889_ _16914_/A _16889_/B _16889_/C vssd1 vssd1 vccd1 vccd1 _19608_/D sky130_fd_sc_hd__nor3_1
XFILLER_38_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10384__S1 _10263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09430_ _11007_/A vssd1 vssd1 vccd1 vccd1 _09431_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_65_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18628_ _18964_/CLK _18628_/D vssd1 vssd1 vccd1 vccd1 _18628_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14424__A0 _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09361_ _13132_/A _09322_/X _09360_/X vssd1 vssd1 vccd1 vccd1 _18745_/D sky130_fd_sc_hd__o21ai_1
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18559_ _18894_/CLK _18559_/D vssd1 vssd1 vccd1 vccd1 _18559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14817__S _14821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10136__S1 _09871_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13721__S _13725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_143_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09292_ _12621_/B vssd1 vssd1 vccd1 vccd1 _09292_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09500__A _09500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11241__S _11241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09603__B1 _09602_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput130 _12479_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[29] sky130_fd_sc_hd__buf_2
Xoutput141 _11544_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wr_en sky130_fd_sc_hd__buf_2
XANTENNA__13163__A0 _19726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput152 _16286_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[19] sky130_fd_sc_hd__buf_2
Xoutput163 _12397_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[29] sky130_fd_sc_hd__buf_2
XFILLER_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10072__S0 _09500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_68_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13692__A _18091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15383__S _15383_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09628_ _10640_/A vssd1 vssd1 vccd1 vccd1 _09628_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_44_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13218__B2 _19350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _18644_/Q vssd1 vssd1 vccd1 vccd1 _11022_/A sky130_fd_sc_hd__inv_2
XFILLER_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13631__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _16790_/B _12518_/X _12569_/X _12538_/X vssd1 vssd1 vccd1 vccd1 _12570_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_169_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_141_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09842__B1 _10195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17904__A1 _12389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09410__A _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11521_ _11646_/C _11521_/B _11521_/C _11523_/C vssd1 vssd1 vccd1 vccd1 _11521_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_168_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14240_ _18627_/Q _14007_/X _14242_/S vssd1 vssd1 vccd1 vccd1 _14241_/A sky130_fd_sc_hd__mux2_1
X_11452_ _11452_/A _11452_/B vssd1 vssd1 vccd1 vccd1 _11452_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_149_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10403_ _19315_/Q _18727_/Q _18764_/Q _18338_/Q _09681_/A _10238_/A vssd1 vssd1 vccd1
+ vccd1 _10404_/B sky130_fd_sc_hd__mux4_1
X_14171_ _14182_/A vssd1 vssd1 vccd1 vccd1 _14180_/S sky130_fd_sc_hd__clkbuf_4
X_11383_ _11371_/X _11382_/X _09667_/X _09758_/X _19738_/Q vssd1 vssd1 vccd1 vccd1
+ _12422_/A sky130_fd_sc_hd__a32oi_4
XFILLER_139_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17132__A2 _17131_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10334_ _18468_/Q _19059_/Q _19221_/Q _18436_/Q _10215_/S _10272_/A vssd1 vssd1 vccd1
+ vccd1 _10335_/B sky130_fd_sc_hd__mux4_1
XANTENNA_input61_A io_ibus_inst[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15143__A1 _15057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ _12855_/X _13113_/X _13116_/X _13121_/X vssd1 vssd1 vccd1 vccd1 _15051_/A
+ sky130_fd_sc_hd__o31a_4
XFILLER_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13053_ _19469_/Q vssd1 vssd1 vccd1 vccd1 _16458_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ _17930_/A vssd1 vssd1 vccd1 vccd1 _19740_/D sky130_fd_sc_hd__clkbuf_1
X_10265_ _10378_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10265_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12004_ _12004_/A _17214_/A vssd1 vssd1 vccd1 vccd1 _12005_/B sky130_fd_sc_hd__or2_1
X_17861_ _17852_/X _17580_/Y _17859_/X _17860_/X vssd1 vssd1 vccd1 vccd1 _17861_/X
+ sky130_fd_sc_hd__o211a_1
X_10196_ _19191_/Q _18805_/Q _19255_/Q _18374_/Q _09854_/X _09676_/A vssd1 vssd1 vccd1
+ vccd1 _10197_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output148_A _16276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ _16812_/A vssd1 vssd1 vccd1 vccd1 _16812_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__17074__A _17085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19600_ _19603_/CLK _19600_/D vssd1 vssd1 vccd1 vccd1 _19600_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_120_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17792_ _17626_/X _17789_/X _17791_/Y _17589_/X vssd1 vssd1 vccd1 vccd1 _17792_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_66_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19531_ _19543_/CLK _19531_/D vssd1 vssd1 vccd1 vccd1 _19531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16743_ _19557_/Q _16739_/B _16742_/Y vssd1 vssd1 vccd1 vccd1 _19557_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13955_ _13955_/A vssd1 vssd1 vccd1 vccd1 _18514_/D sky130_fd_sc_hd__clkbuf_1
X_19462_ _19607_/CLK _19462_/D vssd1 vssd1 vccd1 vccd1 _19462_/Q sky130_fd_sc_hd__dfxtp_1
X_12906_ _15015_/A vssd1 vssd1 vccd1 vccd1 _14537_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16674_ _19533_/Q _16679_/D _16673_/Y vssd1 vssd1 vccd1 vccd1 _19533_/D sky130_fd_sc_hd__o21a_1
XANTENNA__12011__A _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14406__A0 _13886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ _14566_/A vssd1 vssd1 vccd1 vccd1 _13886_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18413_ _19264_/CLK _18413_/D vssd1 vssd1 vccd1 vccd1 _18413_/Q sky130_fd_sc_hd__dfxtp_1
X_15625_ _15612_/X _18280_/Q _09234_/X _13398_/X _15624_/X vssd1 vssd1 vccd1 vccd1
+ _15625_/X sky130_fd_sc_hd__a32o_2
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09508__S0 _10518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _19666_/Q _12703_/X _12704_/X _19633_/Q vssd1 vssd1 vccd1 vccd1 _12837_/X
+ sky130_fd_sc_hd__a22o_1
X_19393_ _19854_/CLK _19393_/D vssd1 vssd1 vccd1 vccd1 _19393_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_61_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12968__A0 _19715_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18344_ _19256_/CLK _18344_/D vssd1 vssd1 vccd1 vccd1 _18344_/Q sky130_fd_sc_hd__dfxtp_1
X_15556_ _19723_/Q _12550_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15556_/X sky130_fd_sc_hd__mux2_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _18275_/Q _12766_/X _10087_/A _12762_/X vssd1 vssd1 vccd1 vccd1 _18275_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09320__A _16245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14507_ _13928_/X _18737_/Q _14511_/S vssd1 vssd1 vccd1 vccd1 _14508_/A sky130_fd_sc_hd__mux2_1
X_18275_ _19725_/CLK _18275_/D vssd1 vssd1 vccd1 vccd1 _18275_/Q sky130_fd_sc_hd__dfxtp_1
X_11719_ _19854_/Q vssd1 vssd1 vccd1 vccd1 _18116_/A sky130_fd_sc_hd__buf_4
XANTENNA__10466__A _10509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ _15478_/X _15485_/X _15486_/Y _13403_/X hold19/X vssd1 vssd1 vccd1 vccd1
+ _15487_/X sky130_fd_sc_hd__a32o_4
X_12699_ _13054_/A vssd1 vssd1 vccd1 vccd1 _12699_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_159_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17226_ _17446_/S vssd1 vssd1 vccd1 vccd1 _17512_/S sky130_fd_sc_hd__clkbuf_2
Xinput10 io_dbus_rdata[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_4
X_14438_ _14438_/A vssd1 vssd1 vccd1 vccd1 _18706_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput21 io_dbus_rdata[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
Xinput32 io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_2
Xinput43 io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
Xinput54 io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__15468__S _15482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17157_ _17160_/A _17157_/B vssd1 vssd1 vccd1 vccd1 _17158_/A sky130_fd_sc_hd__and2_1
XANTENNA__09974__B _12473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput65 io_ibus_inst[9] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_1
X_14369_ _13940_/X _18677_/Q _14369_/S vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16108_ _16107_/A _16107_/C _13195_/X vssd1 vssd1 vccd1 vccd1 _16108_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_143_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17088_ _19690_/Q _15608_/X _17094_/S vssd1 vssd1 vccd1 vccd1 _17089_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16039_ _16039_/A _19748_/Q _16039_/C vssd1 vssd1 vccd1 vccd1 _16046_/B sky130_fd_sc_hd__or3_1
XFILLER_124_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10903__C1 _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_112_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19729_ _19780_/CLK _19729_/D vssd1 vssd1 vccd1 vccd1 _19729_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15931__S _15937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09413_ _10660_/A vssd1 vssd1 vccd1 vccd1 _10764_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_80_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _17121_/B _11647_/A vssd1 vssd1 vccd1 vccd1 _11620_/A sky130_fd_sc_hd__or2_1
XFILLER_34_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13081__C1 _13080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__B1 _09823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09275_ _16625_/A _12508_/C _12584_/A vssd1 vssd1 vccd1 vccd1 _13356_/B sky130_fd_sc_hd__nor3_4
XANTENNA__11631__B1 _11596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10293__S0 _10286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_106_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10315__S _10315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10050_ _09665_/A _10040_/X _10049_/X _09756_/A _19734_/Q vssd1 vssd1 vccd1 vccd1
+ _10080_/A sky130_fd_sc_hd__a32o_4
XANTENNA__10045__S0 _09441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09405__A _09596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13740_ _13740_/A vssd1 vssd1 vccd1 vccd1 _18437_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10952_ _19304_/Q _18716_/Q _18753_/Q _18327_/Q _09396_/A _10937_/A vssd1 vssd1 vccd1
+ vccd1 _10953_/B sky130_fd_sc_hd__mux4_1
XANTENNA__16928__A2 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17050__A1 _15515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13671_ _13228_/X _18407_/Q _13675_/S vssd1 vssd1 vccd1 vccd1 _13672_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12766__A _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _18782_/Q vssd1 vssd1 vccd1 vccd1 _10883_/X sky130_fd_sc_hd__buf_2
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15410_ _15410_/A vssd1 vssd1 vccd1 vccd1 _19112_/D sky130_fd_sc_hd__clkbuf_1
X_12622_ _12652_/B vssd1 vssd1 vccd1 vccd1 _14518_/B sky130_fd_sc_hd__buf_2
XFILLER_71_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16390_ _16390_/A _16396_/C vssd1 vssd1 vccd1 vccd1 _16390_/Y sky130_fd_sc_hd__nor2_1
XFILLER_25_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15341_ _15387_/S vssd1 vssd1 vccd1 vccd1 _15350_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_169_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ _19623_/Q _18079_/B _12553_/C vssd1 vssd1 vccd1 vccd1 _12553_/X sky130_fd_sc_hd__or3_1
XFILLER_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ _11504_/A vssd1 vssd1 vccd1 vccd1 _18743_/D sky130_fd_sc_hd__clkbuf_1
X_18060_ _18060_/A vssd1 vssd1 vccd1 vccd1 _19799_/D sky130_fd_sc_hd__clkbuf_1
X_15272_ _14557_/X _19051_/Q _15278_/S vssd1 vssd1 vccd1 vccd1 _15273_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _17207_/A vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__clkbuf_2
X_17011_ _19657_/Q _17011_/B vssd1 vssd1 vccd1 vccd1 _17011_/X sky130_fd_sc_hd__or2_1
XFILLER_8_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14223_ _18619_/Q _13981_/X _14231_/S vssd1 vssd1 vccd1 vccd1 _14224_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11435_ _11435_/A _11437_/A _11435_/C vssd1 vssd1 vccd1 vccd1 _11435_/Y sky130_fd_sc_hd__nand3_1
XFILLER_165_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14154_ _18589_/Q _13988_/X _14158_/S vssd1 vssd1 vccd1 vccd1 _14155_/A sky130_fd_sc_hd__mux2_1
X_11366_ _11368_/A _11365_/X _09730_/X vssd1 vssd1 vccd1 vccd1 _11366_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10317_ _18931_/Q _18697_/Q _19379_/Q _19027_/Q _10367_/S _10314_/A vssd1 vssd1 vccd1
+ vccd1 _10317_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13105_ _13105_/A _13105_/B vssd1 vssd1 vccd1 vccd1 _15047_/A sky130_fd_sc_hd__and2_4
XFILLER_125_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18962_ _18964_/CLK _18962_/D vssd1 vssd1 vccd1 vccd1 _18962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_112_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14085_ _13886_/X _18559_/Q _14085_/S vssd1 vssd1 vccd1 vccd1 _14086_/A sky130_fd_sc_hd__mux2_1
X_11297_ _18622_/Q _18957_/Q _11297_/S vssd1 vssd1 vccd1 vccd1 _11298_/B sky130_fd_sc_hd__mux2_1
XANTENNA__14920__S _14926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10036__S0 _09441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ _19190_/Q _18804_/Q _19254_/Q _18373_/Q _10247_/X _10238_/X vssd1 vssd1 vccd1
+ vccd1 _10249_/B sky130_fd_sc_hd__mux4_1
XFILLER_140_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _17673_/X _17384_/X _17912_/Y vssd1 vssd1 vccd1 vccd1 _17913_/Y sky130_fd_sc_hd__o21ai_1
X_13036_ _11538_/X _13034_/X _13035_/X vssd1 vssd1 vccd1 vccd1 _15035_/A sky130_fd_sc_hd__o21a_4
X_18893_ _19373_/CLK _18893_/D vssd1 vssd1 vccd1 vccd1 _18893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_152_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16420__B _16833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13536__S _13545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17844_ _17842_/X _17843_/Y _17844_/S vssd1 vssd1 vccd1 vccd1 _17844_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09751__C1 _09740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10179_ _09762_/X _10165_/X _10177_/X _09835_/X _10178_/Y vssd1 vssd1 vccd1 vccd1
+ _12471_/B sky130_fd_sc_hd__o32a_4
XFILLER_113_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17775_ _17779_/A _17779_/B _17775_/S vssd1 vssd1 vccd1 vccd1 _17775_/X sky130_fd_sc_hd__mux2_1
X_14987_ _14987_/A vssd1 vssd1 vccd1 vccd1 _18939_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16726_ _16762_/A _16731_/C vssd1 vssd1 vccd1 vccd1 _16726_/Y sky130_fd_sc_hd__nor2_1
X_19514_ _19543_/CLK _19514_/D vssd1 vssd1 vccd1 vccd1 _19514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13938_ _13937_/X _18511_/Q _13941_/S vssd1 vssd1 vccd1 vccd1 _13939_/A sky130_fd_sc_hd__mux2_1
X_19445_ _19583_/CLK _19445_/D vssd1 vssd1 vccd1 vccd1 _19445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12098__D _12098_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16657_ _19525_/Q _19524_/Q _16657_/C vssd1 vssd1 vccd1 vccd1 _16659_/C sky130_fd_sc_hd__and3_1
XFILLER_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13869_ _13869_/A vssd1 vssd1 vccd1 vccd1 _18489_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14367__S _14369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11580__A _12442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15608_ _15565_/X _15606_/X _15607_/Y _15549_/X _18277_/Q vssd1 vssd1 vccd1 vccd1
+ _15608_/X sky130_fd_sc_hd__a32o_2
XFILLER_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19376_ _19376_/CLK _19376_/D vssd1 vssd1 vccd1 vccd1 _19376_/Q sky130_fd_sc_hd__dfxtp_1
X_16588_ _19510_/Q _16586_/B _16587_/Y vssd1 vssd1 vccd1 vccd1 _19510_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_16_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10416__A1 _09674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18327_ _19306_/CLK _18327_/D vssd1 vssd1 vccd1 vccd1 _18327_/Q sky130_fd_sc_hd__dfxtp_1
X_15539_ _15539_/A vssd1 vssd1 vccd1 vccd1 _19151_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_147_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18258_ _19720_/CLK _18258_/D vssd1 vssd1 vccd1 vccd1 _18258_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_120_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17209_ _17438_/S vssd1 vssd1 vccd1 vccd1 _17501_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__15198__S _15206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18189_ input36/X _18178_/X _18188_/X _18174_/X _19846_/Q vssd1 vssd1 vccd1 vccd1
+ _18190_/B sky130_fd_sc_hd__a32o_1
XFILLER_156_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11916__A1 _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16314__C _19474_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09990__C1 _09989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14830__S _14832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09962_ _09909_/X _09951_/Y _09957_/X _09961_/Y _09813_/A vssd1 vssd1 vccd1 vccd1
+ _09962_/X sky130_fd_sc_hd__o311a_2
XFILLER_103_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09893_ _09952_/S vssd1 vssd1 vccd1 vccd1 _10166_/S sky130_fd_sc_hd__clkbuf_4
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A1 _12337_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13446__S _13448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10578__S1 _10577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09225__A _11619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12586__A _19506_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16058__A _16086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09327_ _09327_/A vssd1 vssd1 vccd1 vccd1 _17115_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ _19825_/Q vssd1 vssd1 vccd1 vccd1 _09267_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_138_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13357__B1 _12586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09189_ _11511_/A _11511_/B _17184_/A _09188_/X vssd1 vssd1 vccd1 vccd1 _11678_/A
+ sky130_fd_sc_hd__or4b_4
XANTENNA__10834__A _18642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11220_ _11220_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11220_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_134_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12580__A1 _19626_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ _18612_/Q _18947_/Q _11151_/S vssd1 vssd1 vccd1 vccd1 _11151_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14740__S _14748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10102_ _19193_/Q _18807_/Q _19257_/Q _18376_/Q _10093_/S _09715_/A vssd1 vssd1 vccd1
+ vccd1 _10103_/B sky130_fd_sc_hd__mux4_1
XFILLER_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _11026_/A _11081_/X _11042_/X vssd1 vssd1 vccd1 vccd1 _11082_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14910_ _14910_/A vssd1 vssd1 vccd1 vccd1 _18901_/D sky130_fd_sc_hd__clkbuf_1
X_10033_ _09589_/A _10032_/X _09982_/A vssd1 vssd1 vccd1 vccd1 _10033_/X sky130_fd_sc_hd__a21o_1
XFILLER_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15890_ _19281_/Q _14569_/A _15898_/S vssd1 vssd1 vccd1 vccd1 _15891_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14841_ _18871_/Q _14023_/X _14843_/S vssd1 vssd1 vccd1 vccd1 _14842_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input24_A io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10894__A1 _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13880__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17560_ _17563_/A _17563_/B vssd1 vssd1 vccd1 vccd1 _17560_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14772_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14781_/S sky130_fd_sc_hd__buf_4
XFILLER_95_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11984_ _11984_/A _17218_/A vssd1 vssd1 vccd1 vccd1 _11985_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16511_ _19599_/Q _19598_/Q _19600_/Q _16857_/A vssd1 vssd1 vccd1 vccd1 _16865_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_90_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13723_ _13070_/X _18430_/Q _13725_/S vssd1 vssd1 vccd1 vccd1 _13724_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17491_ _17504_/S vssd1 vssd1 vccd1 vccd1 _17716_/S sky130_fd_sc_hd__buf_2
X_10935_ _11011_/A vssd1 vssd1 vccd1 vccd1 _11196_/S sky130_fd_sc_hd__buf_4
XFILLER_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14187__S _14191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__A _17133_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13091__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19230_ _19326_/CLK _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Q sky130_fd_sc_hd__dfxtp_1
X_16442_ _16442_/A _16442_/B _16442_/C vssd1 vssd1 vccd1 vccd1 _19464_/D sky130_fd_sc_hd__nor3_1
XFILLER_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ _13654_/A vssd1 vssd1 vccd1 vccd1 _18399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10866_ _10073_/A _10848_/Y _10859_/X _10865_/Y _09658_/A vssd1 vssd1 vccd1 vccd1
+ _10866_/X sky130_fd_sc_hd__o311a_2
XFILLER_13_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12605_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12605_/Y sky130_fd_sc_hd__nor2_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19161_ _19161_/CLK _19161_/D vssd1 vssd1 vccd1 vccd1 _19161_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16373_ _19440_/Q _16373_/B vssd1 vssd1 vccd1 vccd1 _16379_/C sky130_fd_sc_hd__and2_1
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13585_ _13585_/A vssd1 vssd1 vccd1 vccd1 _18374_/D sky130_fd_sc_hd__clkbuf_1
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10797_ _10798_/A _12454_/A vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__or2_1
XFILLER_158_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18112_ _18112_/A _18116_/B vssd1 vssd1 vccd1 vccd1 _18112_/X sky130_fd_sc_hd__or2_1
XFILLER_13_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15324_ _19074_/Q _15006_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15325_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12536_ _12600_/B _12536_/B vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__nor2_1
X_19092_ _19286_/CLK _19092_/D vssd1 vssd1 vccd1 vccd1 _19092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18043_ _18043_/A vssd1 vssd1 vccd1 vccd1 _19791_/D sky130_fd_sc_hd__clkbuf_1
X_15255_ _15255_/A vssd1 vssd1 vccd1 vccd1 _19043_/D sky130_fd_sc_hd__clkbuf_1
X_12467_ _12468_/A _12467_/B vssd1 vssd1 vccd1 vccd1 _12467_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output92_A _12389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ _14206_/A vssd1 vssd1 vccd1 vccd1 _18611_/D sky130_fd_sc_hd__clkbuf_1
X_11418_ _11418_/A _12479_/B vssd1 vssd1 vccd1 vccd1 _11418_/Y sky130_fd_sc_hd__nor2_1
XFILLER_99_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15186_ _15243_/S vssd1 vssd1 vccd1 vccd1 _15195_/S sky130_fd_sc_hd__buf_2
X_12398_ _18144_/A _11516_/X _12302_/X vssd1 vssd1 vccd1 vccd1 _12398_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_126_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15746__S _15754_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14137_ _14137_/A vssd1 vssd1 vccd1 vccd1 _18581_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14650__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11349_ _11445_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__and2_1
XFILLER_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14068_ _13861_/X _18551_/Q _14074_/S vssd1 vssd1 vccd1 vccd1 _14069_/A sky130_fd_sc_hd__mux2_1
X_18945_ _19736_/CLK _18945_/D vssd1 vssd1 vccd1 vccd1 _18945_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15047__A _15047_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _19748_/Q _19749_/Q _13019_/C vssd1 vssd1 vccd1 vccd1 _13031_/B sky130_fd_sc_hd__and3_1
X_18876_ _19390_/CLK _18876_/D vssd1 vssd1 vccd1 vccd1 _18876_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12874__A2 _12603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__A3 _11191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10885__A1 _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17827_ _17871_/A _17827_/B vssd1 vssd1 vccd1 vccd1 _17827_/X sky130_fd_sc_hd__or2_1
XFILLER_94_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10980__S1 _09513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17758_ _17419_/A _17755_/X _17757_/Y _17541_/A vssd1 vssd1 vccd1 vccd1 _17758_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16709_ _16715_/C _16715_/D _16675_/X vssd1 vssd1 vccd1 vccd1 _16709_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11834__B1 _16086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17689_ _17937_/A vssd1 vssd1 vccd1 vccd1 _17873_/S sky130_fd_sc_hd__clkbuf_2
X_19428_ _19694_/CLK _19428_/D vssd1 vssd1 vccd1 vccd1 _19428_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15576__A1 _15574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19359_ _19660_/CLK _19359_/D vssd1 vssd1 vccd1 vccd1 _19359_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_22_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09112_ _19839_/Q vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_149_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13339__B1 _12521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10654__A _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__S0 _10247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_132_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15656__S _15660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16341__A _16341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09945_ _19290_/Q _19128_/Q _18537_/Q _18307_/Q _10186_/S _09713_/A vssd1 vssd1 vccd1
+ vccd1 _09946_/B sky130_fd_sc_hd__mux4_1
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09876_ _09730_/A _09863_/X _09865_/X _09875_/X _09754_/X vssd1 vssd1 vccd1 vccd1
+ _09876_/X sky130_fd_sc_hd__a311o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17253__A1 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10876__A1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__B1 _19399_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _19180_/Q _18794_/Q _19244_/Q _18363_/Q _10631_/S _10623_/A vssd1 vssd1 vccd1
+ vccd1 _10721_/B sky130_fd_sc_hd__mux4_1
XFILLER_13_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_191_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _10655_/A vssd1 vssd1 vccd1 vccd1 _11298_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_16_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14735__S _14737_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10582_ _10585_/A _10578_/X _10581_/X vssd1 vssd1 vccd1 vccd1 _10582_/Y sky130_fd_sc_hd__o21ai_1
X_13370_ _19770_/Q _13370_/B vssd1 vssd1 vccd1 vccd1 _13370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12321_ _12321_/A _12339_/C vssd1 vssd1 vccd1 vccd1 _12322_/D sky130_fd_sc_hd__nand2_1
XFILLER_166_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12482__C _12482_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__S0 _09700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15040_ _15040_/A vssd1 vssd1 vccd1 vccd1 _18956_/D sky130_fd_sc_hd__clkbuf_1
X_12252_ _12252_/A vssd1 vssd1 vccd1 vccd1 _12252_/Y sky130_fd_sc_hd__inv_2
XFILLER_170_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11203_ _11208_/A _11200_/X _11202_/X _18782_/Q vssd1 vssd1 vccd1 vccd1 _11203_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12183_ _16993_/A _12205_/C vssd1 vssd1 vccd1 vccd1 _12183_/X sky130_fd_sc_hd__or2_1
XFILLER_107_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14470__S _14478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11134_ _18782_/Q vssd1 vssd1 vccd1 vccd1 _11134_/X sky130_fd_sc_hd__clkbuf_2
X_16991_ _19650_/Q _16998_/B vssd1 vssd1 vccd1 vccd1 _16991_/X sky130_fd_sc_hd__or2_1
XFILLER_96_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18730_ _19380_/CLK _18730_/D vssd1 vssd1 vccd1 vccd1 _18730_/Q sky130_fd_sc_hd__dfxtp_1
X_15942_ _13535_/X _19304_/Q _15948_/S vssd1 vssd1 vccd1 vccd1 _15943_/A sky130_fd_sc_hd__mux2_1
X_11065_ _11065_/A vssd1 vssd1 vccd1 vccd1 _11128_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_49_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10016_ _10016_/A vssd1 vssd1 vccd1 vccd1 _10016_/Y sky130_fd_sc_hd__inv_2
XFILLER_76_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18661_ _19249_/CLK _18661_/D vssd1 vssd1 vccd1 vccd1 _18661_/Q sky130_fd_sc_hd__dfxtp_1
X_15873_ _15873_/A vssd1 vssd1 vccd1 vccd1 _19273_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12003__B _17214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13814__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14824_ _18863_/Q _13997_/X _14832_/S vssd1 vssd1 vccd1 vccd1 _14825_/A sky130_fd_sc_hd__mux2_1
X_17612_ _17654_/A _17610_/Y _17611_/X vssd1 vssd1 vccd1 vccd1 _17612_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18592_ _19119_/CLK _18592_/D vssd1 vssd1 vccd1 vccd1 _18592_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12608__A2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ _17532_/X _17538_/X _17540_/Y _17542_/X vssd1 vssd1 vccd1 vccd1 _17543_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10619__A1 _09995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14755_ _14576_/X _18833_/Q _14759_/S vssd1 vssd1 vccd1 vccd1 _14756_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11816__B1 _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11967_ _16974_/A _11994_/C _11966_/Y vssd1 vssd1 vccd1 vccd1 _11974_/A sky130_fd_sc_hd__o21a_1
XFILLER_45_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10739__A _10769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17547__A2 _17430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13706_ _12907_/X _18422_/Q _13714_/S vssd1 vssd1 vccd1 vccd1 _13707_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19312_/CLK sky130_fd_sc_hd__clkbuf_16
X_10918_ _19177_/Q _18791_/Q _19241_/Q _18360_/Q _09625_/A _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10919_/B sky130_fd_sc_hd__mux4_1
X_17474_ _17434_/X _17454_/X _17470_/X _17473_/X vssd1 vssd1 vccd1 vccd1 _17474_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16755__B1 _16718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14686_ _14686_/A vssd1 vssd1 vccd1 vccd1 _18802_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11898_ _11899_/A _17205_/A vssd1 vssd1 vccd1 vccd1 _11900_/A sky130_fd_sc_hd__nand2_1
X_16425_ _16442_/A _16425_/B _16425_/C vssd1 vssd1 vccd1 vccd1 _19458_/D sky130_fd_sc_hd__nor3_1
X_19213_ _19245_/CLK _19213_/D vssd1 vssd1 vccd1 vccd1 _19213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13637_ _13637_/A vssd1 vssd1 vccd1 vccd1 _18391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10849_ _18641_/Q vssd1 vssd1 vccd1 vccd1 _11263_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_60_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19144_ _19421_/CLK _19144_/D vssd1 vssd1 vccd1 vccd1 _19144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15330__A _15387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16356_ _16390_/A _16363_/C vssd1 vssd1 vccd1 vccd1 _16356_/Y sky130_fd_sc_hd__nor2_1
X_13568_ _18369_/Q _13567_/X _13577_/S vssd1 vssd1 vccd1 vccd1 _13569_/A sky130_fd_sc_hd__mux2_1
X_15307_ _14608_/X _19067_/Q _15311_/S vssd1 vssd1 vccd1 vccd1 _15308_/A sky130_fd_sc_hd__mux2_1
XANTENNA__12792__A1 _13399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12519_ _18118_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _13009_/A sky130_fd_sc_hd__nor2_2
X_19075_ _19108_/CLK _19075_/D vssd1 vssd1 vccd1 vccd1 _19075_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16287_ _16287_/A vssd1 vssd1 vccd1 vccd1 _19411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_157_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13499_ _13311_/X _18348_/Q _13503_/S vssd1 vssd1 vccd1 vccd1 _13500_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18026_ _18026_/A vssd1 vssd1 vccd1 vccd1 _19784_/D sky130_fd_sc_hd__clkbuf_1
X_15238_ _15238_/A vssd1 vssd1 vccd1 vccd1 _19036_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14380__S _14384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15169_ _19006_/Q _15095_/X _15171_/S vssd1 vssd1 vccd1 vccd1 _15170_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09730_ _09730_/A vssd1 vssd1 vccd1 vccd1 _09730_/X sky130_fd_sc_hd__clkbuf_2
X_18928_ _19120_/CLK _18928_/D vssd1 vssd1 vccd1 vccd1 _18928_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_86_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09661_ _09617_/X _09642_/X _09659_/X _09579_/A _09660_/Y vssd1 vssd1 vccd1 vccd1
+ _12480_/B sky130_fd_sc_hd__o32a_4
XFILLER_95_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18859_ _19374_/CLK _18859_/D vssd1 vssd1 vccd1 vccd1 _18859_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15505__A hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ _09590_/X _09591_/X _10743_/A vssd1 vssd1 vccd1 vccd1 _09592_/X sky130_fd_sc_hd__a21o_1
XFILLER_82_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12848__B _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09503__A _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11283__B2 _12442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14555__S _14567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12864__A _15009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11035__A1 _11033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10641__S0 _09519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_138_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09928_ _18936_/Q _18702_/Q _19384_/Q _19032_/Q _09840_/S _10090_/A vssd1 vssd1 vccd1
+ vccd1 _09929_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12838__A2 _12784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09859_ _09859_/A _09859_/B _09859_/C vssd1 vssd1 vccd1 vccd1 _09859_/X sky130_fd_sc_hd__or3_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _19592_/Q vssd1 vssd1 vccd1 vccd1 _16845_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11821_/A _11821_/B vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__nor2_2
XFILLER_45_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09413__A _10660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09467__A1 _09726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _14540_/A vssd1 vssd1 vccd1 vccd1 _18752_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11752_ _16951_/A _11810_/S _11750_/X _11751_/Y vssd1 vssd1 vccd1 vccd1 _11752_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_121_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09132__B _18081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ _19717_/Q vssd1 vssd1 vccd1 vccd1 _10703_/Y sky130_fd_sc_hd__inv_2
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14471_ _14471_/A vssd1 vssd1 vccd1 vccd1 _18720_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11683_ _11683_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11683_/X sky130_fd_sc_hd__xor2_4
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16246__A _16848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16210_ _16210_/A vssd1 vssd1 vccd1 vccd1 _19377_/D sky130_fd_sc_hd__clkbuf_1
X_13422_ _16109_/A _13422_/B vssd1 vssd1 vccd1 vccd1 _13423_/B sky130_fd_sc_hd__and2_2
X_17190_ _17190_/A _17432_/B vssd1 vssd1 vccd1 vccd1 _17415_/A sky130_fd_sc_hd__or2_1
X_10634_ _10693_/A _10634_/B vssd1 vssd1 vccd1 vccd1 _10634_/Y sky130_fd_sc_hd__nand2_1
XFILLER_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ _16141_/A vssd1 vssd1 vccd1 vccd1 _19354_/D sky130_fd_sc_hd__clkbuf_1
X_13353_ _19168_/Q _12956_/B _12956_/Y vssd1 vssd1 vccd1 vccd1 _13353_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10294__A _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10565_ _09369_/A _10555_/X _10564_/X _09472_/A _19721_/Q vssd1 vssd1 vccd1 vccd1
+ _10597_/A sky130_fd_sc_hd__a32o_2
XANTENNA__17162__B1 _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12304_ _12301_/X _12476_/B _12303_/Y vssd1 vssd1 vccd1 vccd1 _17867_/A sky130_fd_sc_hd__o21ai_4
X_16072_ _16072_/A vssd1 vssd1 vccd1 vccd1 _19342_/D sky130_fd_sc_hd__clkbuf_1
X_13284_ _19690_/Q _12529_/A _12521_/A _19657_/Q vssd1 vssd1 vccd1 vccd1 _13284_/X
+ sky130_fd_sc_hd__a22o_1
X_10496_ _10496_/A vssd1 vssd1 vccd1 vccd1 _10496_/X sky130_fd_sc_hd__buf_2
XFILLER_170_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13809__S _13809_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15296__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15023_ _18951_/Q _15022_/X _15029_/S vssd1 vssd1 vccd1 vccd1 _15024_/A sky130_fd_sc_hd__mux2_1
X_12235_ _19653_/Q _12256_/C vssd1 vssd1 vccd1 vccd1 _12235_/X sky130_fd_sc_hd__and2_1
X_19831_ _19834_/CLK _19831_/D vssd1 vssd1 vccd1 vccd1 _19831_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12166_ _12167_/A _17202_/A vssd1 vssd1 vccd1 vccd1 _12168_/A sky130_fd_sc_hd__and2_1
XANTENNA__15476__A0 _15475_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14279__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14279__B2 _09351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11117_ _19268_/Q _19106_/Q _18515_/Q _18285_/Q _11112_/X _10910_/A vssd1 vssd1 vccd1
+ vccd1 _11117_/X sky130_fd_sc_hd__mux4_1
XFILLER_2_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19762_ _19793_/CLK _19762_/D vssd1 vssd1 vccd1 vccd1 _19762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16974_ _16974_/A _16984_/B vssd1 vssd1 vccd1 vccd1 _16974_/X sky130_fd_sc_hd__or2_1
X_12097_ _19405_/Q _19406_/Q _12097_/C _12097_/D vssd1 vssd1 vccd1 vccd1 _12098_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18713_ _19205_/CLK _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/Q sky130_fd_sc_hd__dfxtp_1
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11048_/X sky130_fd_sc_hd__or2_1
XFILLER_65_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15925_ _15925_/A vssd1 vssd1 vccd1 vccd1 _19297_/D sky130_fd_sc_hd__clkbuf_1
X_19693_ _19693_/CLK _19693_/D vssd1 vssd1 vccd1 vccd1 _19693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput8 io_dbus_rdata[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15856_ _15924_/S vssd1 vssd1 vccd1 vccd1 _15865_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_37_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18644_ _19711_/CLK _18644_/D vssd1 vssd1 vccd1 vccd1 _18644_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12668__B _18263_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09323__A _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14807_ _14807_/A vssd1 vssd1 vccd1 vccd1 _18855_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15787_ _13519_/X _19235_/Q _15793_/S vssd1 vssd1 vccd1 vccd1 _15788_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18575_ _19296_/CLK _18575_/D vssd1 vssd1 vccd1 vccd1 _18575_/Q sky130_fd_sc_hd__dfxtp_1
X_12999_ _14550_/A vssd1 vssd1 vccd1 vccd1 _12999_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17526_ _17524_/X _17525_/X _17577_/S vssd1 vssd1 vccd1 vccd1 _17526_/X sky130_fd_sc_hd__mux2_1
X_14738_ _14738_/A vssd1 vssd1 vccd1 vccd1 _18825_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16728__B1 _16718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17457_ _17573_/S _17457_/B vssd1 vssd1 vccd1 vccd1 _17457_/X sky130_fd_sc_hd__or2_2
X_14669_ _14669_/A vssd1 vssd1 vccd1 vccd1 _18794_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14203__A1 _13953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16408_ _19452_/Q _16411_/C vssd1 vssd1 vccd1 vccd1 _16409_/B sky130_fd_sc_hd__and2_1
XANTENNA__15060__A _15060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17388_ _17478_/A vssd1 vssd1 vccd1 vccd1 _17597_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_164_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19012_/CLK sky130_fd_sc_hd__clkbuf_16
X_16339_ _16340_/B _16340_/C _19430_/Q vssd1 vssd1 vccd1 vccd1 _16341_/B sky130_fd_sc_hd__a21oi_1
XFILLER_145_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19127_ _19127_/CLK _19127_/D vssd1 vssd1 vccd1 vccd1 _19127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17153__B1 _17140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19058_ _19058_/CLK _19058_/D vssd1 vssd1 vccd1 vccd1 _19058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13719__S _13725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18009_ _18009_/A vssd1 vssd1 vccd1 vccd1 _19776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_179_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19366_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_102_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19581_/CLK sky130_fd_sc_hd__clkbuf_16
X_09713_ _09713_/A vssd1 vssd1 vccd1 vccd1 _09714_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__11179__S1 _11177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09697__A1 _10138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09644_ _09644_/A _09644_/B vssd1 vssd1 vccd1 vccd1 _09644_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09575_ _09575_/A _09575_/B _09230_/B vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__or3b_4
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_117_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19838_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16719__B1 _16718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09544__S1 _09768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_64_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__A1 _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11103__S1 _11020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _10394_/A _10349_/X _10297_/X vssd1 vssd1 vccd1 vccd1 _10350_/X sky130_fd_sc_hd__o21a_1
XFILLER_152_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13629__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ _18405_/Q _18666_/Q _18565_/Q _18900_/Q _10339_/S _10270_/A vssd1 vssd1 vccd1
+ vccd1 _10281_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13181__A1 _19158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _12020_/A vssd1 vssd1 vccd1 vccd1 _12020_/X sky130_fd_sc_hd__buf_2
XFILLER_133_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13181__B2 _19348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__A _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15844__S _15848_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10053__S _10785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13971_ _13971_/A vssd1 vssd1 vccd1 vccd1 _18519_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12769__A _12769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15710_ _15710_/A _16169_/A vssd1 vssd1 vccd1 vccd1 _15767_/A sky130_fd_sc_hd__nand2_4
XFILLER_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12922_ input29/X _12781_/A _12921_/X _12831_/X vssd1 vssd1 vccd1 vccd1 _15019_/A
+ sky130_fd_sc_hd__a22o_2
X_16690_ _16707_/A _16697_/D vssd1 vssd1 vccd1 vccd1 _16690_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15641_ _14519_/X _19170_/Q _15649_/S vssd1 vssd1 vccd1 vccd1 _15642_/A sky130_fd_sc_hd__mux2_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _12853_/A vssd1 vssd1 vccd1 vccd1 _18285_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10289__A _10289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _11743_/C _11804_/B vssd1 vssd1 vccd1 vccd1 _11805_/D sky130_fd_sc_hd__and2b_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18360_ _19239_/CLK _18360_/D vssd1 vssd1 vccd1 vccd1 _18360_/Q sky130_fd_sc_hd__dfxtp_1
X_15572_ _18271_/Q _15572_/B vssd1 vssd1 vccd1 vccd1 _15572_/X sky130_fd_sc_hd__or2_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12895_/A vssd1 vssd1 vccd1 vccd1 _12784_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17311_ _17317_/A _17415_/A _17726_/B vssd1 vssd1 vccd1 vccd1 _17321_/B sky130_fd_sc_hd__or3_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14519_/X _18747_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__mux2_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18291_ _19308_/CLK _18291_/D vssd1 vssd1 vccd1 vccd1 _18291_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _19395_/Q _11736_/C _19396_/Q vssd1 vssd1 vccd1 vccd1 _11737_/A sky130_fd_sc_hd__a21oi_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14195__S _14195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19603_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17242_ _17238_/X _17338_/B _17266_/A vssd1 vssd1 vccd1 vccd1 _17242_/X sky130_fd_sc_hd__mux2_1
X_14454_ _13851_/X _18713_/Q _14456_/S vssd1 vssd1 vccd1 vccd1 _14455_/A sky130_fd_sc_hd__mux2_1
X_11666_ _11662_/Y _11664_/X _11665_/X vssd1 vssd1 vccd1 vccd1 _11666_/Y sky130_fd_sc_hd__o21ai_2
X_13405_ _12230_/X _13404_/X _11706_/B vssd1 vssd1 vccd1 vccd1 _13405_/X sky130_fd_sc_hd__a21bo_1
XFILLER_128_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10617_ _10617_/A _10617_/B vssd1 vssd1 vccd1 vccd1 _10617_/X sky130_fd_sc_hd__or2_1
X_17173_ _17917_/B _17432_/A vssd1 vssd1 vccd1 vccd1 _17173_/X sky130_fd_sc_hd__or2_1
X_14385_ _14385_/A vssd1 vssd1 vccd1 vccd1 _18682_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_167_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11597_ _11672_/S vssd1 vssd1 vccd1 vccd1 _12730_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_116_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _16123_/X _19351_/Q _16140_/S vssd1 vssd1 vccd1 vccd1 _16125_/A sky130_fd_sc_hd__mux2_1
X_13336_ _19768_/Q _13336_/B vssd1 vssd1 vccd1 vccd1 _13362_/B sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_96_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19583_/CLK sky130_fd_sc_hd__clkbuf_16
X_10548_ _09688_/A _10546_/X _11313_/A vssd1 vssd1 vccd1 vccd1 _10548_/X sky130_fd_sc_hd__a21o_1
XFILLER_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13539__S _13545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11970__A2 _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16055_ _16055_/A _16055_/B _16055_/C vssd1 vssd1 vccd1 vccd1 _16064_/B sky130_fd_sc_hd__or3_1
X_13267_ _19449_/Q _12962_/X _13266_/X vssd1 vssd1 vccd1 vccd1 _13267_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10479_ _18497_/Q _18992_/Q _10479_/S vssd1 vssd1 vccd1 vccd1 _10480_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15006_ _15006_/A vssd1 vssd1 vccd1 vccd1 _15006_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12218_ _12220_/A _12219_/A vssd1 vssd1 vccd1 vccd1 _12221_/A sky130_fd_sc_hd__and2_1
XFILLER_170_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13198_ _19685_/Q _12659_/X _12680_/X _19652_/Q vssd1 vssd1 vccd1 vccd1 _13198_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_116_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15754__S _15754_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19814_ _19866_/CLK _19814_/D vssd1 vssd1 vccd1 vccd1 _19814_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_111_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12149_ _12149_/A vssd1 vssd1 vccd1 vccd1 _12149_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_97_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19745_ _19779_/CLK _19745_/D vssd1 vssd1 vccd1 vccd1 _19745_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16957_ _19637_/Q _16957_/B vssd1 vssd1 vccd1 vccd1 _16957_/X sky130_fd_sc_hd__or2_1
XANTENNA__12679__A _13009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15908_ _15908_/A vssd1 vssd1 vccd1 vccd1 _19289_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16949__B1 _16915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19676_ _19695_/CLK _19676_/D vssd1 vssd1 vccd1 vccd1 _19676_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_34_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19088_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_38_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16888_ _16887_/A _16887_/C _19608_/Q vssd1 vssd1 vccd1 vccd1 _16889_/C sky130_fd_sc_hd__a21oi_1
XFILLER_92_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18627_ _18964_/CLK _18627_/D vssd1 vssd1 vccd1 vccd1 _18627_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10694__C1 _09644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15839_ _15839_/A vssd1 vssd1 vccd1 vccd1 _15848_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__15621__A0 _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09360_ _11512_/B _12735_/S _17112_/A _09359_/X vssd1 vssd1 vccd1 vccd1 _09360_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18558_ _19311_/CLK _18558_/D vssd1 vssd1 vccd1 vccd1 _18558_/Q sky130_fd_sc_hd__dfxtp_1
X_17509_ _17372_/X _17374_/X _17509_/S vssd1 vssd1 vccd1 vccd1 _17509_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_49_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19377_/CLK sky130_fd_sc_hd__clkbuf_16
X_09291_ _19699_/Q _19698_/Q _19700_/Q vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__or3b_4
XFILLER_36_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18489_ _19369_/CLK _18489_/D vssd1 vssd1 vccd1 vccd1 _18489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_166_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15929__S _15937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__A1 _09597_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16614__A _16666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10844__S0 _10854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput120 _12443_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[1] sky130_fd_sc_hd__buf_2
Xoutput131 _12444_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[2] sky130_fd_sc_hd__buf_2
Xoutput142 _16241_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[0] sky130_fd_sc_hd__buf_2
XANTENNA__13163__A1 _15566_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput153 _16243_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[1] sky130_fd_sc_hd__buf_2
XFILLER_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput164 _16247_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[2] sky130_fd_sc_hd__buf_2
XFILLER_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16101__A1 _19347_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10072__S1 _09507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12589__A _12589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11021__S0 _09624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09627_ _09645_/S vssd1 vssd1 vccd1 vccd1 _10692_/S sky130_fd_sc_hd__buf_4
XFILLER_83_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09558_ _19327_/Q _18739_/Q _18776_/Q _18350_/Q _10518_/S _10261_/A vssd1 vssd1 vccd1
+ vccd1 _09558_/X sky130_fd_sc_hd__mux4_1
XFILLER_169_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09842__A1 _10138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ _10961_/A vssd1 vssd1 vccd1 vccd1 _10848_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11520_ _17120_/C _11569_/B vssd1 vssd1 vccd1 vccd1 _11523_/C sky130_fd_sc_hd__nand2_1
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11088__S0 _10964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11451_ _11451_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11451_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10402_ _10402_/A _10402_/B vssd1 vssd1 vccd1 vccd1 _11443_/A sky130_fd_sc_hd__nor2_1
X_14170_ _14170_/A vssd1 vssd1 vccd1 vccd1 _18596_/D sky130_fd_sc_hd__clkbuf_1
X_11382_ _09730_/X _11373_/X _11377_/X _11381_/X _09859_/A vssd1 vssd1 vccd1 vccd1
+ _11382_/X sky130_fd_sc_hd__a311o_1
XFILLER_125_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ input8/X _13117_/X _13120_/X vssd1 vssd1 vccd1 vccd1 _13121_/X sky130_fd_sc_hd__a21o_1
X_10333_ _10335_/A _10332_/X _09822_/A vssd1 vssd1 vccd1 vccd1 _10333_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_input54_A io_ibus_inst[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _19601_/Q vssd1 vssd1 vccd1 vccd1 _16871_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10264_ _18932_/Q _18698_/Q _19380_/Q _19028_/Q _10260_/X _10263_/X vssd1 vssd1 vccd1
+ vccd1 _10265_/B sky130_fd_sc_hd__mux4_1
XFILLER_78_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12003_ _12004_/A _17214_/A vssd1 vssd1 vccd1 vccd1 _12005_/A sky130_fd_sc_hd__nand2_1
XFILLER_121_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10195_ _10195_/A _10195_/B vssd1 vssd1 vccd1 vccd1 _10195_/X sky130_fd_sc_hd__or2_1
X_17860_ _17860_/A vssd1 vssd1 vccd1 vccd1 _17860_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_79_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14103__A0 _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_94_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16811_ _19577_/Q vssd1 vssd1 vccd1 vccd1 _16816_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17840__A1 _12252_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17791_ _17586_/X _17788_/Y _17790_/Y vssd1 vssd1 vccd1 vccd1 _17791_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_47_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19530_ _19543_/CLK _19530_/D vssd1 vssd1 vccd1 vccd1 _19530_/Q sky130_fd_sc_hd__dfxtp_1
X_16742_ _16762_/A _16742_/B vssd1 vssd1 vccd1 vccd1 _16742_/Y sky130_fd_sc_hd__nor2_1
XFILLER_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13954_ _18514_/Q _13953_/X _13963_/S vssd1 vssd1 vccd1 vccd1 _13955_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12905_ input28/X _12781_/X _12904_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _15015_/A
+ sky130_fd_sc_hd__a22o_2
X_16673_ _16707_/A _16681_/D vssd1 vssd1 vccd1 vccd1 _16673_/Y sky130_fd_sc_hd__nor2_1
X_19461_ _19594_/CLK _19461_/D vssd1 vssd1 vccd1 vccd1 _19461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17802__B _17802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13885_ _13885_/A vssd1 vssd1 vccd1 vccd1 _18494_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14918__S _14926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__B _19406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15603__A _15603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18412_ _19390_/CLK _18412_/D vssd1 vssd1 vccd1 vccd1 _18412_/Q sky130_fd_sc_hd__dfxtp_1
X_12836_ _18318_/Q _12603_/A _12640_/X _19330_/Q vssd1 vssd1 vccd1 vccd1 _12836_/X
+ sky130_fd_sc_hd__a22o_1
X_15624_ _13344_/X _15613_/Y _18280_/Q vssd1 vssd1 vccd1 vccd1 _15624_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09508__S1 _10261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19392_ _19416_/CLK _19392_/D vssd1 vssd1 vccd1 vccd1 _19392_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_36_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12968__A1 _15505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15555_ _15555_/A vssd1 vssd1 vccd1 vccd1 _19153_/D sky130_fd_sc_hd__clkbuf_1
X_18343_ _19320_/CLK _18343_/D vssd1 vssd1 vccd1 vccd1 _18343_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11850__B _17245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _18274_/Q _12766_/X _11357_/A _12762_/X vssd1 vssd1 vccd1 vccd1 _18274_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17756__A_N _12089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10979__B1 _09561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13123__A _15051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14506_ _14506_/A vssd1 vssd1 vccd1 vccd1 _18736_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09320__B _18071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18274_ _19725_/CLK _18274_/D vssd1 vssd1 vccd1 vccd1 _18274_/Q sky130_fd_sc_hd__dfxtp_1
X_11718_ _12050_/A _11842_/A vssd1 vssd1 vccd1 vccd1 _11725_/A sky130_fd_sc_hd__nor2_1
X_15486_ _15494_/A hold19/A vssd1 vssd1 vccd1 vccd1 _15486_/Y sky130_fd_sc_hd__nand2_1
X_12698_ _12782_/A vssd1 vssd1 vccd1 vccd1 _12939_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11079__S0 _09496_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17225_ _17225_/A vssd1 vssd1 vccd1 vccd1 _17446_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_52_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14437_ _13931_/X _18706_/Q _14439_/S vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__mux2_1
X_11649_ _19394_/Q _11649_/B vssd1 vssd1 vccd1 vccd1 _11649_/Y sky130_fd_sc_hd__nor2_1
Xinput11 io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_4
XFILLER_156_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16434__A _16868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput22 io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
XFILLER_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13393__A1 _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput33 io_dbus_valid vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_4
XFILLER_174_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput44 io_ibus_inst[19] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_2
X_17156_ _17174_/A _17149_/X _17140_/X _19704_/Q vssd1 vssd1 vccd1 vccd1 _17157_/B
+ sky130_fd_sc_hd__a22o_1
Xinput55 io_ibus_inst[29] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
X_14368_ _14368_/A vssd1 vssd1 vccd1 vccd1 _18676_/D sky130_fd_sc_hd__clkbuf_1
Xinput66 io_ibus_valid vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_1
XFILLER_143_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16107_ _16107_/A _19760_/Q _16107_/C vssd1 vssd1 vccd1 vccd1 _16116_/B sky130_fd_sc_hd__or3_1
X_13319_ _19484_/Q vssd1 vssd1 vccd1 vccd1 _16501_/B sky130_fd_sc_hd__clkbuf_2
X_17087_ _17087_/A vssd1 vssd1 vccd1 vccd1 _19689_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10482__A _10482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ _14299_/A _15245_/B vssd1 vssd1 vccd1 vccd1 _14356_/A sky130_fd_sc_hd__nand2_2
XFILLER_6_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13145__A1 input10/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16038_ _16038_/A vssd1 vssd1 vccd1 vccd1 _19336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09444__S0 _09441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_12_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11251__S0 _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17989_ _17989_/A vssd1 vssd1 vccd1 vccd1 _19767_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11003__S0 _10940_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19728_ _19731_/CLK _19728_/D vssd1 vssd1 vccd1 vccd1 _19728_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19659_ _19660_/CLK _19659_/D vssd1 vssd1 vccd1 vccd1 _19659_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14828__S _14832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18096__A _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13732__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ _10872_/S vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__15513__A hold18/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12959__B2 _19336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__B _17250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__A _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _19845_/Q _19844_/Q _19843_/Q _11521_/B vssd1 vssd1 vccd1 vccd1 _11647_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _16625_/A _12508_/C _09274_/C vssd1 vssd1 vccd1 vccd1 _12697_/A sky130_fd_sc_hd__nor3_4
XANTENNA__11631__A1 _19844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16344__A _16344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10293__S1 _10275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15394__S _15400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17175__A _17175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__S1 _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13208__A _15067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ _10951_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _10951_/X sky130_fd_sc_hd__or2_1
XFILLER_16_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13670_ _13670_/A vssd1 vssd1 vccd1 vccd1 _18406_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_71_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10882_ _11138_/A _10882_/B vssd1 vssd1 vccd1 vccd1 _10882_/X sky130_fd_sc_hd__or2_1
X_12621_ _16937_/A _12621_/B _16619_/B vssd1 vssd1 vccd1 vccd1 _12652_/B sky130_fd_sc_hd__or3b_1
XFILLER_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10567__A _10586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15340_ _15340_/A vssd1 vssd1 vccd1 vccd1 _19081_/D sky130_fd_sc_hd__clkbuf_1
X_12552_ _16589_/A vssd1 vssd1 vccd1 vccd1 _18079_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11083__C1 _09553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11503_ _11499_/X _11557_/D _11539_/S vssd1 vssd1 vccd1 vccd1 _11504_/A sky130_fd_sc_hd__mux2_1
X_15271_ _15271_/A vssd1 vssd1 vccd1 vccd1 _19050_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12782__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12483_ _12483_/A vssd1 vssd1 vccd1 vccd1 _12483_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17010_ _17010_/A vssd1 vssd1 vccd1 vccd1 _17010_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14222_ _14268_/S vssd1 vssd1 vccd1 vccd1 _14231_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10808__S0 _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ _11437_/A _11435_/C _11435_/A vssd1 vssd1 vccd1 vccd1 _11434_/X sky130_fd_sc_hd__a21o_1
X_14153_ _14153_/A vssd1 vssd1 vccd1 vccd1 _18588_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11365_ _19329_/Q _18741_/Q _18778_/Q _18352_/Q _09704_/X _09733_/X vssd1 vssd1 vccd1
+ vccd1 _11365_/X sky130_fd_sc_hd__mux4_1
XFILLER_152_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13104_ _13095_/Y _13096_/X _13103_/X _13154_/A _13164_/A vssd1 vssd1 vccd1 vccd1
+ _13105_/B sky130_fd_sc_hd__a221o_1
X_10316_ _09690_/A _10315_/X _10237_/X vssd1 vssd1 vccd1 vccd1 _10316_/X sky130_fd_sc_hd__a21o_1
X_18961_ _19089_/CLK _18961_/D vssd1 vssd1 vccd1 vccd1 _18961_/Q sky130_fd_sc_hd__dfxtp_1
X_14084_ _14084_/A vssd1 vssd1 vccd1 vccd1 _18558_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_output160_A _12328_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11296_ _11460_/A _11462_/A _11459_/B _10751_/A _11295_/Y vssd1 vssd1 vccd1 vccd1
+ _11453_/C sky130_fd_sc_hd__a311o_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17085__A _17085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17912_ _17909_/X _17911_/X _17542_/X vssd1 vssd1 vccd1 vccd1 _17912_/Y sky130_fd_sc_hd__a21oi_1
X_13035_ input3/X _12974_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _13035_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10247_ _10413_/S vssd1 vssd1 vccd1 vccd1 _10247_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__11233__S0 _11074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10036__S1 _10031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18892_ _18894_/CLK _18892_/D vssd1 vssd1 vccd1 vccd1 _18892_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14502__A _14502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_186_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17843_ _17845_/A _17845_/B vssd1 vssd1 vccd1 vccd1 _17843_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10178_ _19729_/Q vssd1 vssd1 vccd1 vccd1 _10178_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09315__B _09315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17774_ _19724_/Q _17570_/X _17773_/X vssd1 vssd1 vccd1 vccd1 _19724_/D sky130_fd_sc_hd__o21a_1
XFILLER_94_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14986_ _18939_/Q vssd1 vssd1 vccd1 vccd1 _14987_/A sky130_fd_sc_hd__clkbuf_1
X_19513_ _19543_/CLK _19513_/D vssd1 vssd1 vccd1 vccd1 _19513_/Q sky130_fd_sc_hd__dfxtp_1
X_16725_ _16754_/C vssd1 vssd1 vccd1 vccd1 _16731_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13937_ _14617_/A vssd1 vssd1 vccd1 vccd1 _13937_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14648__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13552__S _13561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19444_ _19583_/CLK _19444_/D vssd1 vssd1 vccd1 vccd1 _19444_/Q sky130_fd_sc_hd__dfxtp_1
X_16656_ _19523_/Q _19522_/Q _16656_/C vssd1 vssd1 vccd1 vccd1 _16657_/C sky130_fd_sc_hd__and3_1
XFILLER_35_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13868_ _13867_/X _18489_/Q _13871_/S vssd1 vssd1 vccd1 vccd1 _13869_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09331__A _09331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _18317_/Q _12603_/X _12784_/X _19139_/Q _12818_/X vssd1 vssd1 vccd1 vccd1
+ _12819_/X sky130_fd_sc_hd__a221o_1
X_15607_ _15607_/A _18277_/Q vssd1 vssd1 vccd1 vccd1 _15607_/Y sky130_fd_sc_hd__nand2_1
XFILLER_90_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19375_ _19375_/CLK _19375_/D vssd1 vssd1 vccd1 vccd1 _19375_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17329__B1 _09322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16587_ _16610_/A _16596_/C vssd1 vssd1 vccd1 vccd1 _16587_/Y sky130_fd_sc_hd__nor2_1
X_13799_ _13799_/A vssd1 vssd1 vccd1 vccd1 _18463_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18326_ _19305_/CLK _18326_/D vssd1 vssd1 vccd1 vccd1 _18326_/Q sky130_fd_sc_hd__dfxtp_1
X_15538_ _15537_/X _19151_/Q _15544_/S vssd1 vssd1 vccd1 vccd1 _15539_/A sky130_fd_sc_hd__mux2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10821__C1 _09614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15469_ _15468_/X _19139_/Q _15483_/S vssd1 vssd1 vccd1 vccd1 _15470_/A sky130_fd_sc_hd__mux2_1
XFILLER_148_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18257_ _19734_/CLK _18257_/D vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__12692__A _18071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17208_ _17204_/X _17206_/X _17241_/A vssd1 vssd1 vccd1 vccd1 _17208_/X sky130_fd_sc_hd__mux2_1
XFILLER_162_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _18188_/A vssd1 vssd1 vccd1 vccd1 _18188_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_128_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17139_ _17139_/A vssd1 vssd1 vccd1 vccd1 _19699_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09961_ _09964_/A _09958_/X _09960_/X vssd1 vssd1 vccd1 vccd1 _09961_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11129__B1 _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18057__A1 _19419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09892_ _10218_/A vssd1 vssd1 vccd1 vccd1 _10169_/A sky130_fd_sc_hd__clkbuf_4
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09506__A _09506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__B _11918_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__A1 _09765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15815__A0 _13560_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17568__B1 _09322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14558__S _14567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13462__S _13470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12586__B _12586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__A _09241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09326_ _11513_/A vssd1 vssd1 vccd1 vccd1 _11487_/S sky130_fd_sc_hd__buf_2
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09257_ _19823_/Q vssd1 vssd1 vccd1 vccd1 _11803_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09188_ _17145_/B _11541_/A _09188_/C vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__and3_1
XFILLER_135_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16802__A _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14306__A0 _13848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11150_ _10904_/X _11148_/Y _11149_/Y _11020_/X vssd1 vssd1 vccd1 vccd1 _11150_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11383__A3 _09667_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10101_ _09730_/A _10092_/X _10096_/X _10100_/X _09859_/A vssd1 vssd1 vccd1 vccd1
+ _10101_/X sky130_fd_sc_hd__a311o_1
XANTENNA__18048__A1 _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ _18581_/Q _18852_/Q _19076_/Q _18820_/Q _10969_/X _11266_/A vssd1 vssd1 vccd1
+ vccd1 _11081_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11215__S0 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16059__A0 _12669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09416__A _09416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _18508_/Q _19003_/Q _10603_/S vssd1 vssd1 vccd1 vccd1 _10032_/X sky130_fd_sc_hd__mux2_1
XFILLER_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10343__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15852__S _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ _14840_/A vssd1 vssd1 vccd1 vccd1 _18870_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14771_ _14771_/A vssd1 vssd1 vccd1 vccd1 _18840_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_input17_A io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11983_ _11983_/A vssd1 vssd1 vccd1 vccd1 _11985_/A sky130_fd_sc_hd__inv_2
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16510_ _19595_/Q _19597_/Q _19596_/Q _16849_/A vssd1 vssd1 vccd1 vccd1 _16857_/A
+ sky130_fd_sc_hd__and4_1
X_13722_ _13722_/A vssd1 vssd1 vccd1 vccd1 _18429_/D sky130_fd_sc_hd__clkbuf_1
X_10934_ _10934_/A vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10646__A2 _10630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17490_ _17603_/A vssd1 vssd1 vccd1 vccd1 _17490_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16441_ _16440_/A _16440_/C _19464_/Q vssd1 vssd1 vccd1 vccd1 _16442_/C sky130_fd_sc_hd__a21oi_1
X_13653_ _13090_/X _18399_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13654_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10865_ _10839_/A _10860_/X _10864_/X vssd1 vssd1 vccd1 vccd1 _10865_/Y sky130_fd_sc_hd__o21ai_1
X_12604_ _19667_/Q _17028_/A _12603_/X _18319_/Q vssd1 vssd1 vccd1 vccd1 _12604_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12399__A2 _12480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16372_ _16388_/A _16372_/B _16373_/B vssd1 vssd1 vccd1 vccd1 _19439_/D sky130_fd_sc_hd__nor3_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19160_ _19598_/CLK _19160_/D vssd1 vssd1 vccd1 vccd1 _19160_/Q sky130_fd_sc_hd__dfxtp_1
X_13584_ _18374_/Q _13583_/X _13593_/S vssd1 vssd1 vccd1 vccd1 _13585_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10796_ _09617_/A _10782_/X _10794_/X _09578_/A _10795_/Y vssd1 vssd1 vccd1 vccd1
+ _12454_/A sky130_fd_sc_hd__o32a_4
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18111_ _19819_/Q _18106_/X hold23/X _18110_/X vssd1 vssd1 vccd1 vccd1 _19819_/D
+ sky130_fd_sc_hd__o211a_1
X_15323_ _15323_/A vssd1 vssd1 vccd1 vccd1 _19073_/D sky130_fd_sc_hd__clkbuf_1
X_12535_ _19623_/Q _12496_/C _12565_/A _19647_/Q _12534_/X vssd1 vssd1 vccd1 vccd1
+ _12535_/X sky130_fd_sc_hd__a221o_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19091_ _19091_/CLK _19091_/D vssd1 vssd1 vccd1 vccd1 _19091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15254_ _14531_/X _19043_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15255_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18042_ _19791_/Q _19412_/Q _18050_/S vssd1 vssd1 vccd1 vccd1 _18043_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12466_ _12468_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _12466_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_144_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14205_ _18611_/Q _13956_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14206_/A sky130_fd_sc_hd__mux2_1
X_11417_ _11417_/A vssd1 vssd1 vccd1 vccd1 _11417_/Y sky130_fd_sc_hd__inv_2
X_15185_ _15185_/A vssd1 vssd1 vccd1 vccd1 _19012_/D sky130_fd_sc_hd__clkbuf_1
X_12397_ _12391_/A _12319_/X _12393_/X _12396_/Y vssd1 vssd1 vccd1 vccd1 _12397_/X
+ sky130_fd_sc_hd__o22a_4
XFILLER_126_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14136_ _18581_/Q _13962_/X _14136_/S vssd1 vssd1 vccd1 vccd1 _14137_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output85_A _12225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11348_ _10599_/Y _11452_/B _11450_/A _10598_/A vssd1 vssd1 vccd1 vccd1 _11448_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_125_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14067_ _14067_/A vssd1 vssd1 vccd1 vccd1 _18550_/D sky130_fd_sc_hd__clkbuf_1
X_18944_ _19361_/CLK _18944_/D vssd1 vssd1 vccd1 vccd1 _18944_/Q sky130_fd_sc_hd__dfxtp_1
X_11279_ _18449_/Q _19040_/Q _19202_/Q _18417_/Q _10962_/S _11220_/A vssd1 vssd1 vccd1
+ vccd1 _11279_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13520__A1 _13519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13018_ _12994_/A _13019_/C _19749_/Q vssd1 vssd1 vccd1 vccd1 _13020_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12323__A2 _12317_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18875_ _19390_/CLK _18875_/D vssd1 vssd1 vccd1 vccd1 _18875_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17826_ _17673_/X _17648_/X _17825_/Y vssd1 vssd1 vccd1 vccd1 _17826_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13284__B1 _12521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14378__S _14384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17757_ _17812_/A _17752_/X _17756_/X vssd1 vssd1 vccd1 vccd1 _17757_/Y sky130_fd_sc_hd__a21oi_1
X_14969_ _14969_/A vssd1 vssd1 vccd1 vccd1 _18930_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15063__A _15063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16708_ _19545_/Q _16712_/D _16707_/Y vssd1 vssd1 vccd1 vccd1 _19545_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17688_ _17477_/X _17683_/Y _17687_/X _17518_/X _11932_/Y vssd1 vssd1 vccd1 vccd1
+ _17688_/X sky130_fd_sc_hd__a32o_2
XFILLER_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19427_ _19694_/CLK _19427_/D vssd1 vssd1 vccd1 vccd1 _19427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15998__A _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16639_ _16650_/C _16639_/B vssd1 vssd1 vccd1 vccd1 _19523_/D sky130_fd_sc_hd__nor2_1
XFILLER_35_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19358_ _19660_/CLK _19358_/D vssd1 vssd1 vccd1 vccd1 _19358_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_148_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11598__A0 _09331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09111_ _09182_/B vssd1 vssd1 vccd1 vccd1 _18081_/A sky130_fd_sc_hd__buf_2
X_18309_ _19292_/CLK _18309_/D vssd1 vssd1 vccd1 vccd1 _18309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19289_ _19291_/CLK _19289_/D vssd1 vssd1 vccd1 vccd1 _19289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15937__S _15937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10248__S1 _10238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14841__S _14843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16622__A _16622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _18473_/Q _19064_/Q _19226_/Q _18441_/Q _10137_/S _09714_/A vssd1 vssd1 vccd1
+ vccd1 _09944_/X sky130_fd_sc_hd__mux4_1
XFILLER_98_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _10105_/A _09872_/X _09874_/X _09857_/X vssd1 vssd1 vccd1 vccd1 _09875_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input9_A io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10420__S1 _09674_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12597__A _18234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__A1 _11826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_134_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ _10824_/S vssd1 vssd1 vccd1 vccd1 _10650_/X sky130_fd_sc_hd__buf_4
XFILLER_55_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09309_ _19707_/Q vssd1 vssd1 vccd1 vccd1 _09309_/X sky130_fd_sc_hd__buf_6
XFILLER_110_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10487__S1 _10347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10581_ _11335_/A _10580_/X _10074_/A vssd1 vssd1 vccd1 vccd1 _10581_/X sky130_fd_sc_hd__o21a_1
XFILLER_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12320_ _12321_/A _12339_/C vssd1 vssd1 vccd1 vccd1 _12322_/C sky130_fd_sc_hd__or2_1
XFILLER_6_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09629__S0 _10692_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12251_ _12251_/A _12251_/B vssd1 vssd1 vccd1 vccd1 _12252_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12002__A1 _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10239__S1 _10238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14751__S _14759_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16532__A _16714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ _18781_/Q _11202_/B vssd1 vssd1 vccd1 vccd1 _11202_/X sky130_fd_sc_hd__or2_1
XFILLER_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12182_ _19651_/Q vssd1 vssd1 vccd1 vccd1 _16993_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_123_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10564__A1 _09995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11133_ _11248_/A _11133_/B vssd1 vssd1 vccd1 vccd1 _11133_/X sky130_fd_sc_hd__or2_1
XFILLER_150_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16990_ _12593_/B _16983_/X _16989_/X _16981_/X vssd1 vssd1 vccd1 vccd1 _19649_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09146__A _18146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15941_ _15941_/A vssd1 vssd1 vccd1 vccd1 _19303_/D sky130_fd_sc_hd__clkbuf_1
X_11064_ _11064_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11064_/X sky130_fd_sc_hd__or2_1
XFILLER_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10316__A1 _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_59_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10015_ _18507_/Q _19002_/Q _10572_/S vssd1 vssd1 vccd1 vccd1 _10016_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18660_ _18894_/CLK _18660_/D vssd1 vssd1 vccd1 vccd1 _18660_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15872_ _19273_/Q _14544_/A _15876_/S vssd1 vssd1 vccd1 vccd1 _15873_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17611_ _11669_/B _17305_/B _17399_/Y vssd1 vssd1 vccd1 vccd1 _17611_/X sky130_fd_sc_hd__o21a_1
XFILLER_91_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14823_ _14845_/A vssd1 vssd1 vccd1 vccd1 _14832_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13266__B1 _13264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18591_ _19086_/CLK _18591_/D vssd1 vssd1 vccd1 vccd1 _18591_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17542_ _17633_/A vssd1 vssd1 vccd1 vccd1 _17542_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ _16974_/A _11994_/C _16114_/A vssd1 vssd1 vccd1 vccd1 _11966_/Y sky130_fd_sc_hd__a21oi_1
X_14754_ _14754_/A vssd1 vssd1 vccd1 vccd1 _18832_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10175__S0 _10114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13115__B _19723_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13705_ _13762_/S vssd1 vssd1 vccd1 vccd1 _13714_/S sky130_fd_sc_hd__buf_2
X_10917_ _10903_/X _10908_/Y _10912_/Y _10916_/Y _09553_/A vssd1 vssd1 vccd1 vccd1
+ _10917_/X sky130_fd_sc_hd__o221a_1
X_14685_ _14579_/X _18802_/Q _14687_/S vssd1 vssd1 vccd1 vccd1 _14686_/A sky130_fd_sc_hd__mux2_1
X_17473_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17473_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17810__B _17810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16755__A1 _16760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ _19781_/Q _10749_/B _12028_/S vssd1 vssd1 vccd1 vccd1 _17205_/A sky130_fd_sc_hd__mux2_2
XANTENNA__14926__S _14926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19212_ _19247_/CLK _19212_/D vssd1 vssd1 vccd1 vccd1 _19212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16424_ _16423_/A _16423_/B _19458_/Q vssd1 vssd1 vccd1 vccd1 _16425_/C sky130_fd_sc_hd__a21oi_1
X_13636_ _12924_/X _18391_/Q _13642_/S vssd1 vssd1 vccd1 vccd1 _13637_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10848_ _10848_/A _10848_/B vssd1 vssd1 vccd1 vccd1 _10848_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19143_ _19421_/CLK _19143_/D vssd1 vssd1 vccd1 vccd1 _19143_/Q sky130_fd_sc_hd__dfxtp_1
X_16355_ _19434_/Q _19433_/Q _19432_/Q _16355_/D vssd1 vssd1 vccd1 vccd1 _16363_/C
+ sky130_fd_sc_hd__and4_1
X_13567_ _15051_/A vssd1 vssd1 vccd1 vccd1 _13567_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10755__A _11313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ _10779_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _10779_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09642__C1 _09572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12518_ _12518_/A vssd1 vssd1 vccd1 vccd1 _12518_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10252__B1 _09728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15306_ _15306_/A vssd1 vssd1 vccd1 vccd1 _19066_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16286_ _16298_/A _16286_/B vssd1 vssd1 vccd1 vccd1 _16287_/A sky130_fd_sc_hd__and2_1
X_19074_ _19074_/CLK _19074_/D vssd1 vssd1 vccd1 vccd1 _19074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13498_ _13498_/A vssd1 vssd1 vccd1 vccd1 _18347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15757__S _15765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18025_ _19784_/Q _12011_/A _18027_/S vssd1 vssd1 vccd1 vccd1 _18026_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ _12450_/A _12449_/B vssd1 vssd1 vccd1 vccd1 _12449_/Y sky130_fd_sc_hd__nor2_1
X_15237_ _19036_/Q _15089_/X _15239_/S vssd1 vssd1 vccd1 vccd1 _15238_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16442__A _16442_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15168_ _15168_/A vssd1 vssd1 vccd1 vccd1 _19005_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10555__A1 _09995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14119_ _14119_/A vssd1 vssd1 vccd1 vccd1 _18574_/D sky130_fd_sc_hd__clkbuf_1
X_15099_ _18975_/Q _15098_/X _15099_/S vssd1 vssd1 vccd1 vccd1 _15100_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18927_ _19261_/CLK _18927_/D vssd1 vssd1 vccd1 vccd1 _18927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09660_ _19737_/Q vssd1 vssd1 vccd1 vccd1 _09660_/Y sky130_fd_sc_hd__inv_2
XFILLER_68_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18858_ _18974_/CLK _18858_/D vssd1 vssd1 vccd1 vccd1 _18858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17809_ _17810_/A _17810_/B _17842_/S vssd1 vssd1 vccd1 vccd1 _17809_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15505__B _15505_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09591_ _18639_/Q _18974_/Q _10764_/S vssd1 vssd1 vccd1 vccd1 _09591_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18789_ _19239_/CLK _18789_/D vssd1 vssd1 vccd1 vccd1 _18789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__A2 _13619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10665__A _11313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15667__S _15671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14571__S _14583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_145_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10641__S1 _10705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _09927_/A vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_60_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09858_ _10150_/A _09847_/X _09856_/X _09857_/X vssd1 vssd1 vccd1 vccd1 _09859_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_74_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09789_ _10014_/A vssd1 vssd1 vccd1 vccd1 _10277_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16985__A1 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11850_/A _17245_/A vssd1 vssd1 vccd1 vccd1 _11821_/B sky130_fd_sc_hd__nor2_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10157__S0 _10114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ _11750_/A _11750_/B _11708_/A vssd1 vssd1 vccd1 vccd1 _11751_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14746__S _14748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17630__B _17630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _11456_/A _12457_/B vssd1 vssd1 vccd1 vccd1 _11453_/B sky130_fd_sc_hd__nand2_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _13873_/X _18720_/Q _14478_/S vssd1 vssd1 vccd1 vccd1 _14471_/A sky130_fd_sc_hd__mux2_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11682_ _11638_/A _11638_/B _11681_/Y vssd1 vssd1 vccd1 vccd1 _11683_/B sky130_fd_sc_hd__o21ai_4
XFILLER_14_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13421_/A vssd1 vssd1 vccd1 vccd1 _18318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10633_ _18621_/Q _18956_/Q _10633_/S vssd1 vssd1 vccd1 vccd1 _10634_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10575__A _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16140_ _16139_/X _19354_/Q _16140_/S vssd1 vssd1 vccd1 vccd1 _16141_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12774__A2 _12773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13352_ input24/X _13166_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__a21oi_1
XFILLER_6_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10564_ _09995_/X _10557_/X _10559_/X _10563_/X _09752_/A vssd1 vssd1 vccd1 vccd1
+ _10564_/X sky130_fd_sc_hd__a311o_4
XFILLER_154_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17162__A1 _17175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12303_ _18135_/A _11516_/A _12302_/X vssd1 vssd1 vccd1 vccd1 _12303_/Y sky130_fd_sc_hd__o21ai_1
X_16071_ _16070_/X _19342_/Q _16083_/S vssd1 vssd1 vccd1 vccd1 _16072_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13886__A _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13283_ _19546_/Q vssd1 vssd1 vccd1 vccd1 _16715_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14481__S _14489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10495_ _10495_/A _10495_/B vssd1 vssd1 vccd1 vccd1 _11448_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13184__C1 _13183_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15022_ _15022_/A vssd1 vssd1 vccd1 vccd1 _15022_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12234_ _19653_/Q _12256_/C vssd1 vssd1 vccd1 vccd1 _12234_/Y sky130_fd_sc_hd__nor2_1
XFILLER_136_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19830_ _19830_/CLK _19830_/D vssd1 vssd1 vccd1 vccd1 _19830_/Q sky130_fd_sc_hd__dfxtp_1
X_12165_ _19791_/Q _10303_/A _12423_/S vssd1 vssd1 vccd1 vccd1 _17202_/A sky130_fd_sc_hd__mux2_2
XFILLER_123_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11116_ _11116_/A _11116_/B vssd1 vssd1 vccd1 vccd1 _11116_/Y sky130_fd_sc_hd__nor2_1
XFILLER_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19761_ _19793_/CLK _19761_/D vssd1 vssd1 vccd1 vccd1 _19761_/Q sky130_fd_sc_hd__dfxtp_1
X_16973_ _17013_/A vssd1 vssd1 vccd1 vccd1 _16984_/B sky130_fd_sc_hd__clkbuf_1
X_12096_ _19398_/Q _19399_/Q _19402_/Q _19403_/Q vssd1 vssd1 vccd1 vccd1 _12097_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18712_ _19268_/CLK _18712_/D vssd1 vssd1 vccd1 vccd1 _18712_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13825__S _13831_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _18916_/Q _18682_/Q _19364_/Q _19012_/Q _11196_/S _10990_/A vssd1 vssd1 vccd1
+ vccd1 _11048_/B sky130_fd_sc_hd__mux4_1
X_15924_ _19297_/Q _14620_/A _15924_/S vssd1 vssd1 vccd1 vccd1 _15925_/A sky130_fd_sc_hd__mux2_1
X_19692_ _19693_/CLK _19692_/D vssd1 vssd1 vccd1 vccd1 _19692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 io_dbus_rdata[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
X_18643_ _19724_/CLK _18643_/D vssd1 vssd1 vccd1 vccd1 _18643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15855_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15924_/S sky130_fd_sc_hd__buf_6
XANTENNA__10170__C1 _09964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14806_ _18855_/Q _13972_/X _14810_/S vssd1 vssd1 vccd1 vccd1 _14807_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18574_ _19324_/CLK _18574_/D vssd1 vssd1 vccd1 vccd1 _18574_/Q sky130_fd_sc_hd__dfxtp_1
X_15786_ _15786_/A vssd1 vssd1 vccd1 vccd1 _19234_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12998_ _15028_/A vssd1 vssd1 vccd1 vccd1 _14550_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17525_ _17279_/X _17288_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17525_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16728__A1 _16731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14737_ _14550_/X _18825_/Q _14737_/S vssd1 vssd1 vccd1 vccd1 _14738_/A sky130_fd_sc_hd__mux2_1
X_11949_ _11949_/A vssd1 vssd1 vccd1 vccd1 _12111_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15341__A _15387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17456_ _17396_/B _17341_/X _17456_/S vssd1 vssd1 vccd1 vccd1 _17456_/X sky130_fd_sc_hd__mux2_1
X_14668_ _14553_/X _18794_/Q _14676_/S vssd1 vssd1 vccd1 vccd1 _14669_/A sky130_fd_sc_hd__mux2_1
X_16407_ _16442_/A _16407_/B _16411_/C vssd1 vssd1 vccd1 vccd1 _19451_/D sky130_fd_sc_hd__nor3_1
X_13619_ _13619_/A _14371_/B _13619_/C _14642_/C vssd1 vssd1 vccd1 vccd1 _14299_/A
+ sky130_fd_sc_hd__and4_2
XFILLER_32_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17387_ _17404_/C _17387_/B _17404_/B vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__and3b_1
XANTENNA__09615__C1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14599_ _14598_/X _18771_/Q _14599_/S vssd1 vssd1 vccd1 vccd1 _14600_/A sky130_fd_sc_hd__mux2_1
X_19126_ _19127_/CLK _19126_/D vssd1 vssd1 vccd1 vccd1 _19126_/Q sky130_fd_sc_hd__dfxtp_1
X_16338_ _16340_/B _16340_/C _16337_/Y vssd1 vssd1 vccd1 vccd1 _19429_/D sky130_fd_sc_hd__o21a_1
XFILLER_9_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17153__A1 _17122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__S0 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19057_ _19315_/CLK _19057_/D vssd1 vssd1 vccd1 vccd1 _19057_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14391__S _14395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16269_ _16981_/A vssd1 vssd1 vccd1 vccd1 _16269_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_161_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18008_ _19776_/Q _19397_/Q _18016_/S vssd1 vssd1 vccd1 vccd1 _18009_/A sky130_fd_sc_hd__mux2_1
XFILLER_133_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10528__A1 _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16900__A _16915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18099__A _18099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09712_ _09712_/A vssd1 vssd1 vccd1 vccd1 _09713_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12150__B1 _19411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09643_ _18942_/Q _18708_/Q _19390_/Q _19038_/Q _10572_/S _09542_/A vssd1 vssd1 vccd1
+ vccd1 _09644_/B sky130_fd_sc_hd__mux4_1
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10700__A1 _09829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09574_ _18742_/Q vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__inv_2
XFILLER_24_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13470__S _13470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12756__A2 _12752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17178__A _17203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10280_ _10433_/S vssd1 vssd1 vccd1 vccd1 _10339_/S sky130_fd_sc_hd__buf_4
XFILLER_117_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_151_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17906__A _17907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16810__A _16838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19248_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11192__B2 _19710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13645__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14130__A1 _13953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13970_ _18519_/Q _13969_/X _13979_/S vssd1 vssd1 vccd1 vccd1 _13971_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12921_ _12912_/X _12920_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12921_/X sky130_fd_sc_hd__mux2_1
XFILLER_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16958__A1 _15495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15640_ _15708_/S vssd1 vssd1 vccd1 vccd1 _15649_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12851_/X _18285_/Q _12887_/S vssd1 vssd1 vccd1 vccd1 _12853_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15630__A1 hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11803_ _11803_/A vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ _19552_/Q vssd1 vssd1 vccd1 vccd1 _16731_/B sky130_fd_sc_hd__buf_2
X_15571_ _15571_/A vssd1 vssd1 vccd1 vccd1 _19157_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14476__S _14478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__C1 _09844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16257__A _16848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17310_ _17387_/B _17319_/B vssd1 vssd1 vccd1 vccd1 _17726_/B sky130_fd_sc_hd__nand2_2
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11734_/A vssd1 vssd1 vccd1 vccd1 _11734_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522_ _14621_/S vssd1 vssd1 vccd1 vccd1 _14535_/S sky130_fd_sc_hd__clkbuf_4
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18290_ _19305_/CLK _18290_/D vssd1 vssd1 vccd1 vccd1 _18290_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10550__S0 _09415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17241_ _17241_/A vssd1 vssd1 vccd1 vccd1 _17266_/A sky130_fd_sc_hd__clkbuf_2
X_11665_ _11887_/A vssd1 vssd1 vccd1 vccd1 _11665_/X sky130_fd_sc_hd__clkbuf_2
X_14453_ _14453_/A vssd1 vssd1 vccd1 vccd1 _18712_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10207__B1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13404_ _13398_/X _13399_/X _13402_/Y _13403_/X hold21/X vssd1 vssd1 vccd1 vccd1
+ _13404_/X sky130_fd_sc_hd__a32o_4
X_10616_ _19278_/Q _19116_/Q _18525_/Q _18295_/Q _10670_/S _09443_/A vssd1 vssd1 vccd1
+ vccd1 _10617_/B sky130_fd_sc_hd__mux4_1
X_14384_ _13854_/X _18682_/Q _14384_/S vssd1 vssd1 vccd1 vccd1 _14385_/A sky130_fd_sc_hd__mux2_1
X_17172_ _17917_/B _17432_/A vssd1 vssd1 vccd1 vccd1 _17172_/Y sky130_fd_sc_hd__nand2_1
X_11596_ _11596_/A vssd1 vssd1 vccd1 vccd1 _11723_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12009__B _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16123_ _12689_/X _16122_/Y _16156_/S vssd1 vssd1 vccd1 vccd1 _16123_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13335_ _16159_/A _13336_/B vssd1 vssd1 vccd1 vccd1 _13335_/Y sky130_fd_sc_hd__nor2_1
X_10547_ _10547_/A vssd1 vssd1 vccd1 vccd1 _11313_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_143_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13266_ _19577_/Q _13055_/X _13264_/X _13265_/X vssd1 vssd1 vccd1 vccd1 _13266_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_142_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16054_ _16054_/A vssd1 vssd1 vccd1 vccd1 _19339_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10478_ _10471_/Y _10473_/Y _10475_/Y _10477_/Y _09830_/A vssd1 vssd1 vccd1 vccd1
+ _10478_/X sky130_fd_sc_hd__o221a_4
XFILLER_136_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15005_ _15005_/A vssd1 vssd1 vccd1 vccd1 _18945_/D sky130_fd_sc_hd__clkbuf_1
X_12217_ _19793_/Q _10181_/A _12357_/S vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__mux2_4
XFILLER_142_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13197_ _13195_/X _13213_/C _13196_/Y vssd1 vssd1 vccd1 vccd1 _13197_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19813_ _19866_/CLK _19813_/D vssd1 vssd1 vccd1 vccd1 _19813_/Q sky130_fd_sc_hd__dfxtp_1
X_12148_ _12148_/A _12148_/B vssd1 vssd1 vccd1 vccd1 _12149_/A sky130_fd_sc_hd__xnor2_2
XFILLER_116_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11864__A _16963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13555__S _13561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ _19779_/CLK _19744_/D vssd1 vssd1 vccd1 vccd1 _19744_/Q sky130_fd_sc_hd__dfxtp_1
X_16956_ _16970_/A vssd1 vssd1 vccd1 vccd1 _16956_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12079_ _12075_/X _12076_/Y _12104_/B _12440_/A vssd1 vssd1 vccd1 vccd1 _12079_/Y
+ sky130_fd_sc_hd__o31ai_2
XFILLER_111_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15907_ _19289_/Q _14595_/A _15909_/S vssd1 vssd1 vccd1 vccd1 _15908_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09334__A _19864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19675_ _19694_/CLK _19675_/D vssd1 vssd1 vccd1 vccd1 _19675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11486__A2 _11492_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16949__A1 _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16887_ _16887_/A _19608_/Q _16887_/C vssd1 vssd1 vccd1 vccd1 _16889_/B sky130_fd_sc_hd__and3_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15770__S _15776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18626_ _19089_/CLK _18626_/D vssd1 vssd1 vccd1 vccd1 _18626_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15838_ _15838_/A vssd1 vssd1 vccd1 vccd1 _19258_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_25_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15621__A1 _15620_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18557_ _18894_/CLK _18557_/D vssd1 vssd1 vccd1 vccd1 _18557_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15769_ _15769_/A vssd1 vssd1 vccd1 vccd1 _19227_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17508_ _17508_/A vssd1 vssd1 vccd1 vccd1 _17508_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_33_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ _12543_/B _16624_/A _12548_/A vssd1 vssd1 vccd1 vccd1 _16937_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12986__A2 _12817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18488_ _19365_/CLK _18488_/D vssd1 vssd1 vccd1 vccd1 _18488_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17439_ _17439_/A vssd1 vssd1 vccd1 vccd1 _17439_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_159_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19109_ _19109_/CLK _19109_/D vssd1 vssd1 vccd1 vccd1 _19109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_opt_2_0_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15010__S _15013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09509__A _09557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput110 _12456_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[10] sky130_fd_sc_hd__buf_2
XFILLER_161_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11838__A2_N _12453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput121 _12468_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[20] sky130_fd_sc_hd__buf_2
Xoutput132 _12480_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[30] sky130_fd_sc_hd__buf_2
Xoutput143 _16264_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[10] sky130_fd_sc_hd__buf_2
XFILLER_115_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput154 _16288_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[20] sky130_fd_sc_hd__buf_2
Xoutput165 _12418_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[30] sky130_fd_sc_hd__buf_2
XFILLER_142_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15246__A _15302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11021__S1 _11020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15680__S _15682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09626_ _09626_/A vssd1 vssd1 vccd1 vccd1 _09645_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_56_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10780__S0 _09519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ _09557_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09557_/Y sky130_fd_sc_hd__nor2_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09488_ _11232_/A vssd1 vssd1 vccd1 vccd1 _10961_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10988__A1 _10895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11450_ _11450_/A vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__inv_2
XFILLER_109_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11088__S1 _11033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10401_ _10401_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _10402_/B sky130_fd_sc_hd__nor2_1
XFILLER_109_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17668__A2 _17658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _09732_/A _11378_/X _11380_/X _09740_/X vssd1 vssd1 vccd1 vccd1 _11381_/X
+ sky130_fd_sc_hd__o211a_1
X_13120_ _13167_/A vssd1 vssd1 vccd1 vccd1 _13120_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10332_ _19317_/Q _18729_/Q _18766_/Q _18340_/Q _10286_/X _10382_/A vssd1 vssd1 vccd1
+ vccd1 _10332_/X sky130_fd_sc_hd__mux4_1
XFILLER_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11668__B _11668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09419__A _09419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18078__C1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ _13051_/A vssd1 vssd1 vccd1 vccd1 _13051_/X sky130_fd_sc_hd__buf_2
X_10263_ _10482_/A vssd1 vssd1 vccd1 vccd1 _10263_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16540__A _19494_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12002_ _19785_/Q _10597_/A _12143_/S vssd1 vssd1 vccd1 vccd1 _17214_/A sky130_fd_sc_hd__mux2_2
XANTENNA__09453__S1 _09390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_120_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input47_A io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _19319_/Q _18731_/Q _18768_/Q _18342_/Q _09854_/X _09676_/A vssd1 vssd1 vccd1
+ vccd1 _10195_/B sky130_fd_sc_hd__mux4_1
XFILLER_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16810_ _16838_/A _16810_/B _16810_/C vssd1 vssd1 vccd1 vccd1 _19576_/D sky130_fd_sc_hd__nor3_1
XANTENNA__11684__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17790_ _17790_/A _17790_/B vssd1 vssd1 vccd1 vccd1 _17790_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16741_ _19557_/Q _16752_/D _16741_/C vssd1 vssd1 vccd1 vccd1 _16742_/B sky130_fd_sc_hd__and3_1
XFILLER_120_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13953_ _14525_/A vssd1 vssd1 vccd1 vccd1 _13953_/X sky130_fd_sc_hd__buf_2
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_163_clock clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 _19734_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19460_ _19607_/CLK _19460_/D vssd1 vssd1 vccd1 vccd1 _19460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ _12892_/Y _12902_/X _12942_/S vssd1 vssd1 vccd1 vccd1 _12904_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16672_ _19533_/Q _19532_/Q _19531_/Q _16672_/D vssd1 vssd1 vccd1 vccd1 _16681_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_35_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13884_ _13883_/X _18494_/Q _13887_/S vssd1 vssd1 vccd1 vccd1 _13885_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18411_ _19387_/CLK _18411_/D vssd1 vssd1 vccd1 vccd1 _18411_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15623_ _15623_/A vssd1 vssd1 vccd1 vccd1 _19166_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _19554_/Q vssd1 vssd1 vccd1 vccd1 _16736_/B sky130_fd_sc_hd__buf_2
XFILLER_46_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19391_ _19391_/CLK _19391_/D vssd1 vssd1 vccd1 vccd1 _19391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _19619_/CLK _18342_/D vssd1 vssd1 vccd1 vccd1 _18342_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_178_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19272_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15554_ hold9/X _19153_/Q _15570_/S vssd1 vssd1 vccd1 vccd1 _15555_/A sky130_fd_sc_hd__mux2_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12773_/A vssd1 vssd1 vccd1 vccd1 _12766_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14505_ _13925_/X _18736_/Q _14511_/S vssd1 vssd1 vccd1 vccd1 _14506_/A sky130_fd_sc_hd__mux2_1
X_18273_ _19162_/CLK _18273_/D vssd1 vssd1 vccd1 vccd1 _18273_/Q sky130_fd_sc_hd__dfxtp_1
X_11717_ _11717_/A vssd1 vssd1 vccd1 vccd1 _11842_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_182_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12697_ _12697_/A vssd1 vssd1 vccd1 vccd1 _12697_/X sky130_fd_sc_hd__buf_2
X_15485_ hold19/A _15485_/B vssd1 vssd1 vccd1 vccd1 _15485_/X sky130_fd_sc_hd__or2_1
X_17224_ _17220_/X _17223_/X _17241_/A vssd1 vssd1 vccd1 vccd1 _17224_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11648_ _19394_/Q _11649_/B vssd1 vssd1 vccd1 vccd1 _11736_/C sky130_fd_sc_hd__and2_1
X_14436_ _14436_/A vssd1 vssd1 vccd1 vccd1 _18705_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_101_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19635_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_174_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput12 io_dbus_rdata[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
Xinput23 io_dbus_rdata[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_4
Xinput34 io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
X_17155_ _17155_/A vssd1 vssd1 vccd1 vccd1 _19703_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14367_ _13937_/X _18676_/Q _14369_/S vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__mux2_1
X_11579_ _19842_/Q _11542_/A _11572_/X _11578_/X vssd1 vssd1 vccd1 vccd1 _11579_/X
+ sky130_fd_sc_hd__o22a_1
Xinput56 io_ibus_inst[2] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__clkbuf_1
Xinput67 io_irq_motor_irq vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_2
XFILLER_143_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16106_ _16106_/A vssd1 vssd1 vccd1 vccd1 _19348_/D sky130_fd_sc_hd__clkbuf_1
X_13318_ _19616_/Q vssd1 vssd1 vccd1 vccd1 _16912_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_143_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17086_ _19689_/Q _15600_/X _17094_/S vssd1 vssd1 vccd1 vccd1 _17087_/A sky130_fd_sc_hd__mux2_1
X_14298_ _14298_/A vssd1 vssd1 vccd1 vccd1 _15245_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_170_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15765__S _15765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_116_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19699_/CLK sky130_fd_sc_hd__clkbuf_16
X_16037_ _16036_/X _19336_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16038_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13249_ _13249_/A _13249_/B vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__and2_2
XANTENNA__09444__S1 _09443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10364__C1 _09753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10903__A1 _10965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16095__A1 _19346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17292__A0 _17232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11594__A _11668_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17988_ _19767_/Q _19799_/Q _17990_/S vssd1 vssd1 vccd1 vccd1 _17989_/A sky130_fd_sc_hd__mux2_1
XFILLER_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19727_ _19731_/CLK _19727_/D vssd1 vssd1 vccd1 vccd1 _19727_/Q sky130_fd_sc_hd__dfxtp_2
X_16939_ _16939_/A _18071_/S _12565_/X vssd1 vssd1 vccd1 vccd1 _16946_/A sky130_fd_sc_hd__or3b_1
XANTENNA__12656__A1 _16341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__S1 _10990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19658_ _19660_/CLK _19658_/D vssd1 vssd1 vccd1 vccd1 _19658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17595__A1 _19713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18096__B _18142_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ _10873_/S vssd1 vssd1 vccd1 vccd1 _10872_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_80_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18609_ _19361_/CLK _18609_/D vssd1 vssd1 vccd1 vccd1 _18609_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15513__B _15513_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19589_ _19594_/CLK _19589_/D vssd1 vssd1 vccd1 vccd1 _19589_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10938__A _18779_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _18107_/A _19846_/Q vssd1 vssd1 vccd1 vccd1 _11521_/B sky130_fd_sc_hd__or2_1
XANTENNA__12959__A2 _17028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17347__A1 _17294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ _12494_/A _12522_/A _12605_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _16937_/B
+ sky130_fd_sc_hd__nor4b_4
XFILLER_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16307__C1 _12556_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_134_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_162_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12344__B1 _16086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17283__A0 _12289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19162_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_29_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13923__S _13935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ _19176_/Q _18790_/Q _19240_/Q _18359_/Q _09396_/A _10937_/A vssd1 vssd1 vccd1
+ vccd1 _10951_/B sky130_fd_sc_hd__mux4_1
XFILLER_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_95_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19448_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09702__A _09840_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09609_ _10614_/A _09607_/X _09995_/A vssd1 vssd1 vccd1 vccd1 _09609_/X sky130_fd_sc_hd__o21a_1
X_10881_ _18392_/Q _18653_/Q _18552_/Q _18887_/Q _10878_/A _10817_/A vssd1 vssd1 vccd1
+ vccd1 _10882_/B sky130_fd_sc_hd__mux4_1
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12620_ _16935_/A _12598_/X _12716_/S vssd1 vssd1 vccd1 vccd1 _12620_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12551_ _16245_/A vssd1 vssd1 vccd1 vccd1 _16589_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11502_ _17981_/A vssd1 vssd1 vccd1 vccd1 _11539_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_40_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15270_ _14553_/X _19050_/Q _15278_/S vssd1 vssd1 vccd1 vccd1 _15271_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12482_ _12482_/A _12482_/B _12482_/C vssd1 vssd1 vccd1 vccd1 _12483_/A sky130_fd_sc_hd__and3_1
XFILLER_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14221_ _14221_/A vssd1 vssd1 vccd1 vccd1 _18618_/D sky130_fd_sc_hd__clkbuf_1
X_11433_ _11433_/A _11433_/B vssd1 vssd1 vccd1 vccd1 _11433_/Y sky130_fd_sc_hd__nand2_1
XFILLER_138_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10808__S1 _10802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _18569_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14152_ _18588_/Q _13985_/X _14158_/S vssd1 vssd1 vccd1 vccd1 _14153_/A sky130_fd_sc_hd__mux2_1
X_11364_ _11373_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__or2_1
XFILLER_138_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10315_ _18500_/Q _18995_/Q _10315_/S vssd1 vssd1 vccd1 vccd1 _10315_/X sky130_fd_sc_hd__mux2_1
X_13103_ _19722_/Q _15546_/B _13103_/S vssd1 vssd1 vccd1 vccd1 _13103_/X sky130_fd_sc_hd__mux2_1
X_18960_ _19088_/CLK _18960_/D vssd1 vssd1 vccd1 vccd1 _18960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14083_ _13883_/X _18558_/Q _14085_/S vssd1 vssd1 vccd1 vccd1 _14084_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_98_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11295_ _11456_/A _12457_/B vssd1 vssd1 vccd1 vccd1 _11295_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ _17907_/B _17906_/B _17494_/X _17910_/Y vssd1 vssd1 vccd1 vccd1 _17911_/X
+ sky130_fd_sc_hd__o211a_1
X_13034_ _13030_/Y _13064_/C _13032_/X _13234_/A vssd1 vssd1 vccd1 vccd1 _13034_/X
+ sky130_fd_sc_hd__a2bb2o_1
X_10246_ _10406_/A vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18891_ _19310_/CLK _18891_/D vssd1 vssd1 vccd1 vccd1 _18891_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_129_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11233__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19091_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16077__A1 _19343_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17842_ _17845_/A _17845_/B _17842_/S vssd1 vssd1 vccd1 vccd1 _17842_/X sky130_fd_sc_hd__mux2_1
XFILLER_152_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10177_ _10170_/X _10172_/Y _10174_/Y _10176_/Y _09813_/X vssd1 vssd1 vccd1 vccd1
+ _10177_/X sky130_fd_sc_hd__o221a_2
XANTENNA__17813__A2 _17810_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17773_ _12092_/Y _17427_/X _17772_/X _09359_/X vssd1 vssd1 vccd1 vccd1 _17773_/X
+ sky130_fd_sc_hd__a211o_1
X_14985_ _14985_/A vssd1 vssd1 vccd1 vccd1 _18938_/D sky130_fd_sc_hd__clkbuf_1
X_19512_ _19543_/CLK _19512_/D vssd1 vssd1 vccd1 vccd1 _19512_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13833__S _13835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16724_ _19551_/Q _19550_/Q _16724_/C _16724_/D vssd1 vssd1 vccd1 vccd1 _16754_/C
+ sky130_fd_sc_hd__and4_2
X_13936_ _13936_/A vssd1 vssd1 vccd1 vccd1 _18510_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10744__S0 _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19443_ _19583_/CLK _19443_/D vssd1 vssd1 vccd1 vccd1 _19443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16655_ _19529_/Q _16655_/B vssd1 vssd1 vccd1 vccd1 _16660_/B sky130_fd_sc_hd__nor2_1
XFILLER_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13867_ _14547_/A vssd1 vssd1 vccd1 vccd1 _13867_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10664__A3 _18827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15606_ _18277_/Q _15606_/B vssd1 vssd1 vccd1 vccd1 _15606_/X sky130_fd_sc_hd__or2_1
XANTENNA__13134__A _13166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12818_ _19665_/Q _12817_/X _12704_/X _19632_/Q vssd1 vssd1 vccd1 vccd1 _12818_/X
+ sky130_fd_sc_hd__a22o_1
X_19374_ _19374_/CLK _19374_/D vssd1 vssd1 vccd1 vccd1 _19374_/Q sky130_fd_sc_hd__dfxtp_1
X_16586_ _19510_/Q _16586_/B vssd1 vssd1 vccd1 vccd1 _16596_/C sky130_fd_sc_hd__and2_1
XANTENNA__17329__A1 _12488_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13798_ _13090_/X _18463_/Q _13798_/S vssd1 vssd1 vccd1 vccd1 _13799_/A sky130_fd_sc_hd__mux2_1
X_18325_ _19302_/CLK _18325_/D vssd1 vssd1 vccd1 vccd1 _18325_/Q sky130_fd_sc_hd__dfxtp_1
X_15537_ _19720_/Q _15536_/X _15543_/S vssd1 vssd1 vccd1 vccd1 _15537_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _18262_/Q _12744_/X _10677_/A _12747_/X vssd1 vssd1 vccd1 vccd1 _18262_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18256_ _19734_/CLK _18256_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_2
X_15468_ _09315_/B _13410_/X _15482_/S vssd1 vssd1 vccd1 vccd1 _15468_/X sky130_fd_sc_hd__mux2_1
XFILLER_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17207_ _17207_/A vssd1 vssd1 vccd1 vccd1 _17241_/A sky130_fd_sc_hd__clkbuf_2
X_14419_ _14430_/A vssd1 vssd1 vccd1 vccd1 _14428_/S sky130_fd_sc_hd__buf_4
X_18187_ _18187_/A vssd1 vssd1 vccd1 vccd1 _19845_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10493__A _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15399_ _15399_/A vssd1 vssd1 vccd1 vccd1 _19107_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17138_ _17142_/A _17138_/B vssd1 vssd1 vccd1 vccd1 _17139_/A sky130_fd_sc_hd__and2_1
XFILLER_144_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17069_ _17069_/A vssd1 vssd1 vccd1 vccd1 _19681_/D sky130_fd_sc_hd__clkbuf_1
X_09960_ _10209_/A _09959_/X _09909_/A vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__o21a_1
XFILLER_104_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11129__A1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12877__A1 _16752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09891_ _09891_/A vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__buf_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17265__A0 _17779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12213__A _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14839__S _14843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13743__S _13747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17568__A1 _11765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__A _10854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09241__B _17133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _09325_/A vssd1 vssd1 vccd1 vccd1 _11565_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_159_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14574__S _14583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09256_ _19824_/Q vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13357__A2 _12584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09187_ _09171_/B _09124_/A _09124_/B _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1
+ _09188_/C sky130_fd_sc_hd__o2111a_1
XFILLER_107_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17186__A _17190_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10100_ _10105_/A _10097_/X _10099_/X _09857_/X vssd1 vssd1 vccd1 vccd1 _10100_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_1_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11080_ _11085_/A _11080_/B vssd1 vssd1 vccd1 vccd1 _11080_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10328__C1 _09754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_130_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10031_ _10031_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10031_/X sky130_fd_sc_hd__and2_1
XFILLER_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13653__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14770_ _14598_/X _18840_/Q _14770_/S vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11982_ _11984_/A _17218_/A vssd1 vssd1 vccd1 vccd1 _11983_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13721_ _13048_/X _18429_/Q _13725_/S vssd1 vssd1 vccd1 vccd1 _13722_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11681__B _17239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__A _09432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10933_ _10933_/A vssd1 vssd1 vccd1 vccd1 _10934_/A sky130_fd_sc_hd__buf_4
XFILLER_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10646__A3 _10644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__S _11173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16440_ _16440_/A _19464_/Q _16440_/C vssd1 vssd1 vccd1 vccd1 _16442_/B sky130_fd_sc_hd__and3_1
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13652_ _13652_/A vssd1 vssd1 vccd1 vccd1 _18398_/D sky130_fd_sc_hd__clkbuf_1
X_10864_ _10977_/A _10863_/X _09482_/A vssd1 vssd1 vccd1 vccd1 _10864_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13045__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12603_ _12603_/A vssd1 vssd1 vccd1 vccd1 _12603_/X sky130_fd_sc_hd__buf_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16371_ _19439_/Q _19438_/Q _16371_/C vssd1 vssd1 vccd1 vccd1 _16373_/B sky130_fd_sc_hd__and3_1
XFILLER_158_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14793__A1 _13953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13583_ _15067_/A vssd1 vssd1 vccd1 vccd1 _13583_/X sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10795_ _19716_/Q vssd1 vssd1 vccd1 vccd1 _10795_/Y sky130_fd_sc_hd__inv_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18110_ _18136_/A vssd1 vssd1 vccd1 vccd1 _18110_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_55_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _19073_/Q _15003_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15323_/A sky130_fd_sc_hd__mux2_1
XFILLER_40_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12534_ _19628_/Q _16931_/A _12526_/X _19154_/Q _12533_/X vssd1 vssd1 vccd1 vccd1
+ _12534_/X sky130_fd_sc_hd__a221o_1
X_19090_ _19091_/CLK _19090_/D vssd1 vssd1 vccd1 vccd1 _19090_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18041_ _18188_/A vssd1 vssd1 vccd1 vccd1 _18050_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15253_ _15253_/A vssd1 vssd1 vccd1 vccd1 _19042_/D sky130_fd_sc_hd__clkbuf_1
X_12465_ _12468_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _12465_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14204_ _14204_/A vssd1 vssd1 vccd1 vccd1 _18610_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11416_ _11416_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _11417_/A sky130_fd_sc_hd__and2_1
XFILLER_126_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12396_ _12416_/B _12395_/Y _12440_/A vssd1 vssd1 vccd1 vccd1 _12396_/Y sky130_fd_sc_hd__o21ai_2
X_15184_ _19012_/Q _15012_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__mux2_1
XFILLER_125_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14135_ _14135_/A vssd1 vssd1 vccd1 vccd1 _18580_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11347_ _11347_/A _12462_/A vssd1 vssd1 vccd1 vccd1 _11450_/A sky130_fd_sc_hd__and2_1
XFILLER_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_152_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11278_ _11278_/A _11278_/B vssd1 vssd1 vccd1 vccd1 _11278_/Y sky130_fd_sc_hd__nor2_1
X_14066_ _13857_/X _18550_/Q _14074_/S vssd1 vssd1 vccd1 vccd1 _14067_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output78_A _12063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18943_ _19391_/CLK _18943_/D vssd1 vssd1 vccd1 vccd1 _18943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17764__B_N _17215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _10229_/A vssd1 vssd1 vccd1 vccd1 _10229_/X sky130_fd_sc_hd__buf_2
X_13017_ _19717_/Q _15520_/B _13381_/S vssd1 vssd1 vccd1 vccd1 _13017_/X sky130_fd_sc_hd__mux2_1
X_18874_ _19098_/CLK _18874_/D vssd1 vssd1 vccd1 vccd1 _18874_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17798__A1 _17802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17825_ _17822_/X _17824_/X _17646_/A vssd1 vssd1 vccd1 vccd1 _17825_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17756_ _12089_/X _17756_/B vssd1 vssd1 vccd1 vccd1 _17756_/X sky130_fd_sc_hd__and2b_1
X_14968_ _18930_/Q vssd1 vssd1 vccd1 vccd1 _14969_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_48_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12687__B _12687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16707_ _16707_/A _16715_/D vssd1 vssd1 vccd1 vccd1 _16707_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09342__A _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13919_ _13918_/X _18505_/Q _13919_/S vssd1 vssd1 vccd1 vccd1 _13920_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17687_ _17852_/A _17687_/B vssd1 vssd1 vccd1 vccd1 _17687_/X sky130_fd_sc_hd__or2_1
X_14899_ _14899_/A vssd1 vssd1 vccd1 vccd1 _18896_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19426_ _19694_/CLK _19426_/D vssd1 vssd1 vccd1 vccd1 _19426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16638_ _19523_/Q _16635_/B _12556_/X vssd1 vssd1 vccd1 vccd1 _16639_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__13036__A1 _11538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19357_ _19357_/CLK _19357_/D vssd1 vssd1 vccd1 vccd1 _19357_/Q sky130_fd_sc_hd__dfxtp_1
X_16569_ _19504_/Q _16569_/B vssd1 vssd1 vccd1 vccd1 _16575_/C sky130_fd_sc_hd__and2_1
XANTENNA__11598__A1 _09194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09110_ _09182_/C vssd1 vssd1 vccd1 vccd1 _18083_/A sky130_fd_sc_hd__buf_2
X_18308_ _19197_/CLK _18308_/D vssd1 vssd1 vccd1 vccd1 _18308_/Q sky130_fd_sc_hd__dfxtp_1
X_19288_ _19290_/CLK _19288_/D vssd1 vssd1 vccd1 vccd1 _19288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18239_ _18248_/A _18239_/B vssd1 vssd1 vccd1 vccd1 _18240_/A sky130_fd_sc_hd__and2_1
XFILLER_163_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16930__C1 _16269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11112__A _11219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16622__B _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17486__A0 _17504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_104_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09517__A _10056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09943_ _10108_/A _09943_/B vssd1 vssd1 vccd1 vccd1 _09943_/X sky130_fd_sc_hd__or2_1
XANTENNA__11482__C_N _11481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15953__S _15959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09874_ _10197_/A _09874_/B vssd1 vssd1 vccd1 vccd1 _09874_/X sky130_fd_sc_hd__or2_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13473__S _13481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10398__A _19725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12786__B1 _12784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ _19708_/Q vssd1 vssd1 vccd1 vccd1 _09315_/B sky130_fd_sc_hd__buf_6
XFILLER_142_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10580_ _18591_/Q _18862_/Q _19086_/Q _18830_/Q _10579_/X _10060_/A vssd1 vssd1 vccd1
+ vccd1 _10580_/X sky130_fd_sc_hd__mux4_1
XFILLER_166_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__15724__A0 _13531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09239_ _11755_/A vssd1 vssd1 vccd1 vccd1 _12159_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_166_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09629__S1 _09628_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12250_ _12223_/A _12224_/A _12223_/B _12221_/A vssd1 vssd1 vccd1 vccd1 _12251_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_170_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17628__B _17630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ _18386_/Q _18647_/Q _18546_/Q _18881_/Q _11065_/A _11124_/A vssd1 vssd1 vccd1
+ vccd1 _11202_/B sky130_fd_sc_hd__mux4_1
XFILLER_135_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12181_ _11794_/A _12175_/Y _12179_/X _12180_/Y vssd1 vssd1 vccd1 vccd1 _12181_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16024__S _16024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11132_ _18387_/Q _18648_/Q _18547_/Q _18882_/Q _11123_/A _10933_/A vssd1 vssd1 vccd1
+ vccd1 _11133_/B sky130_fd_sc_hd__mux4_1
XFILLER_123_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09427__A _10667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_110_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15863__S _15865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15940_ _13531_/X _19303_/Q _15948_/S vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__mux2_1
X_11063_ _18453_/Q _19044_/Q _19206_/Q _18421_/Q _11011_/X _11012_/X vssd1 vssd1 vccd1
+ vccd1 _11064_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10014_ _10014_/A _10014_/B vssd1 vssd1 vccd1 vccd1 _10014_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15871_ _15871_/A vssd1 vssd1 vccd1 vccd1 _19272_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17610_ _17609_/A _17499_/Y _17609_/Y vssd1 vssd1 vccd1 vccd1 _17610_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_92_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14822_ _14822_/A vssd1 vssd1 vccd1 vccd1 _18862_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14463__A0 _13864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18590_ _19085_/CLK _18590_/D vssd1 vssd1 vccd1 vccd1 _18590_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09565__S0 _10479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17541_ _17541_/A vssd1 vssd1 vccd1 vccd1 _17633_/A sky130_fd_sc_hd__clkbuf_2
X_14753_ _14573_/X _18832_/Q _14759_/S vssd1 vssd1 vccd1 vccd1 _14754_/A sky130_fd_sc_hd__mux2_1
X_11965_ _12074_/A vssd1 vssd1 vccd1 vccd1 _16114_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13704_ _13704_/A vssd1 vssd1 vccd1 vccd1 _18421_/D sky130_fd_sc_hd__clkbuf_1
X_10916_ _11164_/A _10913_/X _10915_/X vssd1 vssd1 vccd1 vccd1 _10916_/Y sky130_fd_sc_hd__o21ai_1
X_17472_ _17860_/A vssd1 vssd1 vccd1 vccd1 _17592_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14684_ _14684_/A vssd1 vssd1 vccd1 vccd1 _18801_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11896_ _11925_/S vssd1 vssd1 vccd1 vccd1 _12028_/S sky130_fd_sc_hd__clkbuf_2
X_19211_ _19243_/CLK _19211_/D vssd1 vssd1 vccd1 vccd1 _19211_/Q sky130_fd_sc_hd__dfxtp_1
X_16423_ _16423_/A _16423_/B _19458_/Q vssd1 vssd1 vccd1 vccd1 _16425_/B sky130_fd_sc_hd__and3_1
XFILLER_60_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ _13635_/A vssd1 vssd1 vccd1 vccd1 _18390_/D sky130_fd_sc_hd__clkbuf_1
X_10847_ _18920_/Q _18686_/Q _19368_/Q _19016_/Q _09626_/A _10837_/X vssd1 vssd1 vccd1
+ vccd1 _10848_/B sky130_fd_sc_hd__mux4_1
X_19142_ _19635_/CLK _19142_/D vssd1 vssd1 vccd1 vccd1 _19142_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12777__B1 _12422_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16354_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16390_/A sky130_fd_sc_hd__buf_2
XFILLER_9_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13566_ _13566_/A vssd1 vssd1 vccd1 vccd1 _18368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10778_ _19275_/Q _19113_/Q _18522_/Q _18292_/Q _10633_/S _09628_/X vssd1 vssd1 vccd1
+ vccd1 _10779_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17704__B2 _11968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10252__A1 _10323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15715__A0 _13519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15305_ _14605_/X _19066_/Q _15311_/S vssd1 vssd1 vccd1 vccd1 _15306_/A sky130_fd_sc_hd__mux2_1
X_12517_ _13055_/A vssd1 vssd1 vccd1 vccd1 _12518_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19073_ _19267_/CLK _19073_/D vssd1 vssd1 vccd1 vccd1 _19073_/Q sky130_fd_sc_hd__dfxtp_1
X_16285_ _16301_/A vssd1 vssd1 vccd1 vccd1 _16298_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17819__A _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16723__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13497_ _13294_/X _18347_/Q _13503_/S vssd1 vssd1 vccd1 vccd1 _13498_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18024_ _18024_/A vssd1 vssd1 vccd1 vccd1 _19783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15236_ _15236_/A vssd1 vssd1 vccd1 vccd1 _19035_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _12450_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12448_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13558__S _13561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11867__A _11890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ _19005_/Q _15092_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15168_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12379_ _17312_/A vssd1 vssd1 vccd1 vccd1 _17404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_5_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09337__A _18146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ _13934_/X _18574_/Q _14118_/S vssd1 vssd1 vccd1 vccd1 _14119_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15098_ _15098_/A vssd1 vssd1 vccd1 vccd1 _15098_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18926_ _19086_/CLK _18926_/D vssd1 vssd1 vccd1 vccd1 _18926_/Q sky130_fd_sc_hd__dfxtp_1
X_14049_ _18544_/Q _14048_/X _14049_/S vssd1 vssd1 vccd1 vccd1 _14050_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14389__S _14395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18857_ _19081_/CLK _18857_/D vssd1 vssd1 vccd1 vccd1 _18857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold18_A hold18/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12698__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09590_ _09590_/A vssd1 vssd1 vccd1 vccd1 _09590_/X sky130_fd_sc_hd__clkbuf_4
X_17808_ _10300_/Y _12727_/X _17807_/X vssd1 vssd1 vccd1 vccd1 _19727_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__14454__A0 _13851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18788_ _19237_/CLK _18788_/D vssd1 vssd1 vccd1 vccd1 _18788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13306__B _13306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17739_ _17309_/B _17738_/X _17739_/S vssd1 vssd1 vccd1 vccd1 _17739_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09556__S0 _10479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19409_ _19699_/CLK _19409_/D vssd1 vssd1 vccd1 vccd1 _19409_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__15521__B hold16/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11115__S0 _11149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12768__B1 _10087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15013__S _15013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14852__S _14854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11991__A1 _11988_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13193__A0 _13191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13468__S _13470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09926_ _09975_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _09926_/Y sky130_fd_sc_hd__nand2_1
XFILLER_131_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09164__A2 _18100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _09857_/A vssd1 vssd1 vccd1 vccd1 _09857_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_100_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09788_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13248__B2 _13144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10157__S1 _09888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15712__A _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16198__A0 _13554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ _11750_/A _11750_/B vssd1 vssd1 vccd1 vccd1 _11750_/X sky130_fd_sc_hd__and2_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09710__A _09710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14748__A1 _18830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10701_ _10678_/Y _09833_/A _09760_/A _10700_/X vssd1 vssd1 vccd1 vccd1 _12457_/B
+ sky130_fd_sc_hd__o22ai_4
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11681_ _11681_/A _17239_/A vssd1 vssd1 vccd1 vccd1 _11681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_42_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11106__S0 _11074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13420_ _13419_/Y _18318_/Q _13424_/S vssd1 vssd1 vccd1 vccd1 _13421_/A sky130_fd_sc_hd__mux2_1
X_10632_ _10632_/A vssd1 vssd1 vccd1 vccd1 _10632_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10234__A1 _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13351_ _13351_/A vssd1 vssd1 vccd1 vccd1 _18312_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10563_ _10559_/A _10560_/X _10562_/X _09989_/X vssd1 vssd1 vccd1 vccd1 _10563_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14762__S _14770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12302_ _12302_/A vssd1 vssd1 vccd1 vccd1 _12302_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16070_ _15542_/X _16069_/Y _16082_/S vssd1 vssd1 vccd1 vccd1 _16070_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _10494_/A _12464_/B vssd1 vssd1 vccd1 vccd1 _10495_/B sky130_fd_sc_hd__nor2_1
X_13282_ _13315_/C _13281_/Y _11499_/X vssd1 vssd1 vccd1 vccd1 _13282_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_136_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_170_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11687__A _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15021_ _15021_/A vssd1 vssd1 vccd1 vccd1 _18950_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12233_ _16114_/A vssd1 vssd1 vccd1 vccd1 _12233_/X sky130_fd_sc_hd__buf_2
XFILLER_136_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ _17802_/A _12164_/B vssd1 vssd1 vccd1 vccd1 _12167_/A sky130_fd_sc_hd__xor2_1
XFILLER_162_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11115_ _18451_/Q _19042_/Q _19204_/Q _18419_/Q _11149_/A _09512_/A vssd1 vssd1 vccd1
+ vccd1 _11116_/B sky130_fd_sc_hd__mux4_1
XFILLER_123_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_150_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16972_ _12651_/X _16970_/X _16971_/X _16968_/X vssd1 vssd1 vccd1 vccd1 _19642_/D
+ sky130_fd_sc_hd__o211a_1
X_12095_ _19400_/Q _19401_/Q _19404_/Q _19407_/Q vssd1 vssd1 vccd1 vccd1 _12097_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_122_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19760_ _19793_/CLK _19760_/D vssd1 vssd1 vccd1 vccd1 _19760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_104_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09591__S _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18711_ _19299_/CLK _18711_/D vssd1 vssd1 vccd1 vccd1 _18711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11046_ _09477_/A _11029_/X _11044_/Y _09577_/A _11045_/Y vssd1 vssd1 vccd1 vccd1
+ _12448_/B sky130_fd_sc_hd__o32a_4
X_15923_ _15923_/A vssd1 vssd1 vccd1 vccd1 _19296_/D sky130_fd_sc_hd__clkbuf_1
X_19691_ _19693_/CLK _19691_/D vssd1 vssd1 vccd1 vccd1 _19691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15606__B _15606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18642_ _19740_/CLK _18642_/D vssd1 vssd1 vccd1 vccd1 _18642_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14002__S _14011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ _15854_/A _15854_/B vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__nor2_4
XFILLER_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14805_ _14805_/A vssd1 vssd1 vccd1 vccd1 _18854_/D sky130_fd_sc_hd__clkbuf_1
X_18573_ _19326_/CLK _18573_/D vssd1 vssd1 vccd1 vccd1 _18573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15785_ _13509_/X _19234_/Q _15793_/S vssd1 vssd1 vccd1 vccd1 _15786_/A sky130_fd_sc_hd__mux2_1
XFILLER_52_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12997_ _12997_/A _12997_/B vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__and2_2
XANTENNA__16718__A _16812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17524_ _17269_/X _17227_/X _17524_/S vssd1 vssd1 vccd1 vccd1 _17524_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16189__A0 _13541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14736_ _14736_/A vssd1 vssd1 vccd1 vccd1 _18824_/D sky130_fd_sc_hd__clkbuf_1
X_11948_ _12025_/A vssd1 vssd1 vccd1 vccd1 _17696_/A sky130_fd_sc_hd__buf_2
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17925__A1 _19738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17455_ _17504_/S vssd1 vssd1 vccd1 vccd1 _17738_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14667_ _14713_/S vssd1 vssd1 vccd1 vccd1 _14676_/S sky130_fd_sc_hd__buf_2
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11879_ _11879_/A _19401_/Q _11879_/C vssd1 vssd1 vccd1 vccd1 _11969_/D sky130_fd_sc_hd__and3_2
XFILLER_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16406_ _19451_/Q _19450_/Q _16406_/C vssd1 vssd1 vccd1 vccd1 _16411_/C sky130_fd_sc_hd__and3_1
XFILLER_60_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13618_ _19811_/Q _14787_/B vssd1 vssd1 vccd1 vccd1 _15926_/A sky130_fd_sc_hd__nor2_4
XFILLER_158_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17386_ _17386_/A vssd1 vssd1 vccd1 vccd1 _17386_/X sky130_fd_sc_hd__clkbuf_2
X_14598_ _14598_/A vssd1 vssd1 vccd1 vccd1 _14598_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19125_ _19287_/CLK _19125_/D vssd1 vssd1 vccd1 vccd1 _19125_/Q sky130_fd_sc_hd__dfxtp_1
X_16337_ _16340_/B _16340_/C _16293_/X vssd1 vssd1 vccd1 vccd1 _16337_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15768__S _15776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13549_ _18363_/Q _13547_/X _13561_/S vssd1 vssd1 vccd1 vccd1 _13550_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14672__S _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19056_ _19314_/CLK _19056_/D vssd1 vssd1 vccd1 vccd1 _19056_/Q sky130_fd_sc_hd__dfxtp_1
X_16268_ _18172_/A vssd1 vssd1 vccd1 vccd1 _16981_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_69_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18007_ _18029_/A vssd1 vssd1 vccd1 vccd1 _18016_/S sky130_fd_sc_hd__clkbuf_2
X_15219_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15228_/S sky130_fd_sc_hd__clkbuf_8
X_16199_ _16199_/A vssd1 vssd1 vccd1 vccd1 _19372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09217__D _19855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_177_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09711_ _10238_/A vssd1 vssd1 vccd1 vccd1 _09712_/A sky130_fd_sc_hd__buf_2
X_18909_ _19292_/CLK _18909_/D vssd1 vssd1 vccd1 vccd1 _18909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12150__A1 _12126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09642_ _09619_/Y _09631_/Y _09634_/Y _09641_/Y _09572_/A vssd1 vssd1 vccd1 vccd1
+ _09642_/X sky130_fd_sc_hd__o221a_2
XFILLER_95_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09573_ _09557_/Y _09564_/Y _09566_/Y _09568_/Y _09829_/A vssd1 vssd1 vccd1 vccd1
+ _09573_/X sky130_fd_sc_hd__o221a_2
XANTENNA__18169__B2 _18083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__S0 _10633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17916__A1 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15678__S _15682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16104__A0 _15574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_104_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13926__S _13935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09909_ _09909_/A vssd1 vssd1 vccd1 vccd1 _09909_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09705__A _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13227__A _15070_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ _19713_/Q _15493_/B _13103_/S vssd1 vssd1 vccd1 vccd1 _12920_/X sky130_fd_sc_hd__mux2_1
XFILLER_74_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12851_ _14528_/A vssd1 vssd1 vccd1 vccd1 _12851_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_62_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14757__S _14759_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11327__S0 _10579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11802_ _11802_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11809_/A sky130_fd_sc_hd__or2_1
XANTENNA__15630__A2 _13359_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15570_ _15569_/X _19157_/Q _15570_/S vssd1 vssd1 vccd1 vccd1 _15571_/A sky130_fd_sc_hd__mux2_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12782_ _12782_/A vssd1 vssd1 vccd1 vccd1 _12782_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09440__A _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14621_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__09940__S0 _10137_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11733_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10586__A _10586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17240_ _17463_/B _12383_/A _17240_/S vssd1 vssd1 vccd1 vccd1 _17338_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10550__S1 _09443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14452_ _13848_/X _18712_/Q _14456_/S vssd1 vssd1 vccd1 vccd1 _14453_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15394__A1 _15003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _19633_/Q _11696_/B _11810_/S _12074_/A vssd1 vssd1 vccd1 vccd1 _11664_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_30_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13403_ _15549_/A vssd1 vssd1 vccd1 vccd1 _13403_/X sky130_fd_sc_hd__buf_2
X_10615_ _18461_/Q _19052_/Q _19214_/Q _18429_/Q _10763_/S _09590_/X vssd1 vssd1 vccd1
+ vccd1 _10615_/X sky130_fd_sc_hd__mux4_1
X_17171_ _17404_/B vssd1 vssd1 vccd1 vccd1 _17432_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__14492__S _14500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14383_ _14383_/A vssd1 vssd1 vccd1 vccd1 _18681_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11595_ _09210_/X _09211_/Y _09168_/X _17145_/A _17145_/B vssd1 vssd1 vccd1 vccd1
+ _11596_/A sky130_fd_sc_hd__o2111a_2
XFILLER_167_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16122_ _16126_/A _16126_/C vssd1 vssd1 vccd1 vccd1 _16122_/Y sky130_fd_sc_hd__xnor2_1
X_13334_ _19768_/Q vssd1 vssd1 vccd1 vccd1 _16159_/A sky130_fd_sc_hd__clkbuf_2
X_10546_ _18495_/Q _18990_/Q _10546_/S vssd1 vssd1 vccd1 vccd1 _10546_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_3_4_0_clock clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_9_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16053_ _16052_/X _19339_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__mux2_1
X_13265_ _13265_/A vssd1 vssd1 vccd1 vccd1 _13265_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10477_ _10535_/A _10476_/X _09821_/A vssd1 vssd1 vccd1 vccd1 _10477_/Y sky130_fd_sc_hd__o21ai_1
X_15004_ _18945_/Q _15003_/X _15013_/S vssd1 vssd1 vccd1 vccd1 _15005_/A sky130_fd_sc_hd__mux2_1
X_12216_ _12404_/S vssd1 vssd1 vccd1 vccd1 _12357_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__10066__S0 _09500_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13196_ _13195_/X _13213_/C _12848_/A vssd1 vssd1 vccd1 vccd1 _13196_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19812_ _19866_/CLK _19812_/D vssd1 vssd1 vccd1 vccd1 _19812_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12147_ _12122_/A _12122_/B _12118_/A vssd1 vssd1 vccd1 vccd1 _12148_/B sky130_fd_sc_hd__a21bo_1
XFILLER_97_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14521__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19743_ _19779_/CLK _19743_/D vssd1 vssd1 vccd1 vccd1 _19743_/Q sky130_fd_sc_hd__dfxtp_1
X_16955_ _15487_/X _16943_/X _16953_/Y _16954_/X vssd1 vssd1 vccd1 vccd1 _19636_/D
+ sky130_fd_sc_hd__o211a_1
X_12078_ _12078_/A vssd1 vssd1 vccd1 vccd1 _12440_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13137__A _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15906_ _15906_/A vssd1 vssd1 vccd1 vccd1 _19288_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09334__B _19863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ _11019_/Y _11023_/Y _11026_/Y _11028_/Y _11044_/A vssd1 vssd1 vccd1 vccd1
+ _11029_/X sky130_fd_sc_hd__o221a_1
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19674_ _19687_/CLK _19674_/D vssd1 vssd1 vccd1 vccd1 _19674_/Q sky130_fd_sc_hd__dfxtp_1
X_16886_ _16887_/A _16887_/C _16885_/Y vssd1 vssd1 vccd1 vccd1 _19607_/D sky130_fd_sc_hd__o21a_1
XFILLER_38_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15837_ _13592_/X _19258_/Q _15837_/S vssd1 vssd1 vccd1 vccd1 _15838_/A sky130_fd_sc_hd__mux2_1
X_18625_ _19089_/CLK _18625_/D vssd1 vssd1 vccd1 vccd1 _18625_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10694__A1 _09547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12976__A _12976_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13571__S _13577_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18556_ _19310_/CLK _18556_/D vssd1 vssd1 vccd1 vccd1 _18556_/Q sky130_fd_sc_hd__dfxtp_1
X_15768_ _13595_/X _19227_/Q _15776_/S vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__mux2_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09350__A _17125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17507_ _17509_/S _17371_/X _17506_/Y vssd1 vssd1 vccd1 vccd1 _17508_/A sky130_fd_sc_hd__a21oi_2
X_14719_ _14719_/A vssd1 vssd1 vccd1 vccd1 _18816_/D sky130_fd_sc_hd__clkbuf_1
X_18487_ _19367_/CLK _18487_/D vssd1 vssd1 vccd1 vccd1 _18487_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15699_ _15699_/A vssd1 vssd1 vccd1 vccd1 _19196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17438_ _17208_/X _17224_/X _17438_/S vssd1 vssd1 vccd1 vccd1 _17439_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17369_ _17506_/B _17368_/Y _17407_/A vssd1 vssd1 vccd1 vccd1 _17369_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19108_ _19108_/CLK _19108_/D vssd1 vssd1 vccd1 vccd1 _19108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19039_ _19383_/CLK _19039_/D vssd1 vssd1 vccd1 vccd1 _19039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput100 _11824_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[7] sky130_fd_sc_hd__buf_2
Xoutput111 _12458_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[11] sky130_fd_sc_hd__buf_2
XANTENNA__11120__A _19709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput122 _12470_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[21] sky130_fd_sc_hd__buf_2
XFILLER_115_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput133 _12483_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[31] sky130_fd_sc_hd__buf_2
XFILLER_126_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput144 _16266_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[11] sky130_fd_sc_hd__buf_2
XFILLER_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput155 _16290_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[21] sky130_fd_sc_hd__buf_2
XFILLER_82_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput166 _12441_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[31] sky130_fd_sc_hd__buf_2
XFILLER_99_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09525__A _10055_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__B1 _12521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13047__A _15038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09625_ _09625_/A vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__buf_2
XFILLER_55_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14577__S _14583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13481__S _13481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16270__C1 _16269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10780__S1 _09506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09556_ _19199_/Q _18813_/Q _19263_/Q _18382_/Q _10479_/S _09768_/A vssd1 vssd1 vccd1
+ vccd1 _09557_/B sky130_fd_sc_hd__mux4_1
XFILLER_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10437__A1 _10275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09487_ _10968_/A vssd1 vssd1 vccd1 vccd1 _11232_/A sky130_fd_sc_hd__buf_2
XFILLER_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10988__A2 _12450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12825__S _13144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11398__C1 _09813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10400_ _10401_/A _12466_/B vssd1 vssd1 vccd1 vccd1 _10402_/A sky130_fd_sc_hd__and2_1
X_11380_ _11380_/A _11380_/B vssd1 vssd1 vccd1 vccd1 _11380_/X sky130_fd_sc_hd__or2_1
XFILLER_164_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10331_ _10390_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10331_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17917__A _17917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12126__A _12126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11030__A _11033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10262_ _10262_/A vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__buf_2
X_13050_ _13050_/A vssd1 vssd1 vccd1 vccd1 _18295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16540__B _16540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13656__S _13664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ _12028_/S vssd1 vssd1 vccd1 vccd1 _12143_/S sky130_fd_sc_hd__clkbuf_2
X_10193_ _09844_/X _10184_/X _10188_/X _10192_/X _09670_/A vssd1 vssd1 vccd1 vccd1
+ _10193_/X sky130_fd_sc_hd__a311o_2
XFILLER_79_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11684__B _18125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16740_ _16752_/D _16741_/C _16739_/Y vssd1 vssd1 vccd1 vccd1 _19556_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17652__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13952_ _13952_/A vssd1 vssd1 vccd1 vccd1 _18513_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11322__C1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17053__A1 _15522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10220__S0 _10112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12903_ _13065_/A vssd1 vssd1 vccd1 vccd1 _12942_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16671_ _16714_/A vssd1 vssd1 vccd1 vccd1 _16707_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_100_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10676__B2 _19718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14487__S _14489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ _14563_/A vssd1 vssd1 vccd1 vccd1 _13883_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16268__A _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12796__A _18744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15622_ _15621_/X _19166_/Q _15627_/S vssd1 vssd1 vccd1 vccd1 _15623_/A sky130_fd_sc_hd__mux2_1
X_18410_ _19197_/CLK _18410_/D vssd1 vssd1 vccd1 vccd1 _18410_/Q sky130_fd_sc_hd__dfxtp_1
X_12834_ _19426_/Q vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_19390_ _19390_/CLK _19390_/D vssd1 vssd1 vccd1 vccd1 _19390_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _19319_/CLK _18341_/D vssd1 vssd1 vccd1 vccd1 _18341_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15603_/A vssd1 vssd1 vccd1 vccd1 _15570_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09913__S0 _09904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12765_ _18273_/Q _12759_/X _10181_/A _12762_/X vssd1 vssd1 vccd1 vccd1 _18273_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_125_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14504_ _14504_/A vssd1 vssd1 vccd1 vccd1 _18735_/D sky130_fd_sc_hd__clkbuf_1
X_18272_ _19162_/CLK _18272_/D vssd1 vssd1 vccd1 vccd1 _18272_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15900__A _15911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11716_ _11668_/B _17256_/A _17393_/A _11716_/D vssd1 vssd1 vccd1 vccd1 _11717_/A
+ sky130_fd_sc_hd__and4b_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15484_ _15484_/A vssd1 vssd1 vccd1 vccd1 _19142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12696_/A input70/X vssd1 vssd1 vccd1 vccd1 _12696_/X sky130_fd_sc_hd__or2_1
XFILLER_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17223_ _17696_/B _17790_/B _17263_/A vssd1 vssd1 vccd1 vccd1 _17223_/X sky130_fd_sc_hd__mux2_1
XFILLER_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14435_ _13928_/X _18705_/Q _14439_/S vssd1 vssd1 vccd1 vccd1 _14436_/A sky130_fd_sc_hd__mux2_1
X_11647_ _11647_/A _11647_/B _11647_/C vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__or3_2
XFILLER_156_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16207__S _16213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput13 io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10287__S0 _10286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput24 io_dbus_rdata[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_4
X_17154_ _17160_/A _17154_/B vssd1 vssd1 vccd1 vccd1 _17155_/A sky130_fd_sc_hd__and2_1
Xinput35 io_ibus_inst[10] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14366_ _14366_/A vssd1 vssd1 vccd1 vccd1 _18675_/D sky130_fd_sc_hd__clkbuf_1
Xinput46 io_ibus_inst[20] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_2
X_11578_ _11575_/X _11577_/X _19855_/Q _11571_/Y vssd1 vssd1 vccd1 vccd1 _11578_/X
+ sky130_fd_sc_hd__o211a_1
Xinput57 io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_2
XFILLER_171_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput68 io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_1
XFILLER_155_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16105_ _16104_/X _19348_/Q _16112_/S vssd1 vssd1 vccd1 vccd1 _16106_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13317_ _13336_/B _13316_/Y _11499_/X vssd1 vssd1 vccd1 vccd1 _13317_/Y sky130_fd_sc_hd__o21ai_1
X_17085_ _17085_/A vssd1 vssd1 vccd1 vccd1 _17094_/S sky130_fd_sc_hd__clkbuf_2
X_10529_ _10522_/X _10524_/Y _10526_/Y _10528_/Y _09812_/A vssd1 vssd1 vccd1 vccd1
+ _10529_/X sky130_fd_sc_hd__o221a_4
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14297_ _18089_/A _14297_/B vssd1 vssd1 vccd1 vccd1 _14298_/A sky130_fd_sc_hd__and2_1
XANTENNA__16731__A _19553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _15509_/X _16035_/Y _16052_/S vssd1 vssd1 vccd1 vccd1 _16036_/X sky130_fd_sc_hd__mux2_1
X_13248_ _13245_/Y _13246_/X _13247_/X _13144_/S _13164_/A vssd1 vssd1 vccd1 vccd1
+ _13249_/B sky130_fd_sc_hd__a221o_1
XFILLER_170_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12353__A1 _18140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13179_ _13179_/A vssd1 vssd1 vccd1 vccd1 _13179_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17292__A1 _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17987_ _17987_/A vssd1 vssd1 vccd1 vccd1 _19766_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_96_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13302__B1 _13301_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19726_ _19740_/CLK _19726_/D vssd1 vssd1 vccd1 vccd1 _19726_/Q sky130_fd_sc_hd__dfxtp_4
X_16938_ _16959_/A vssd1 vssd1 vccd1 vccd1 _16957_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17044__A1 _15495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19657_ _19660_/CLK _19657_/D vssd1 vssd1 vccd1 vccd1 _19657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16869_ _16871_/A _16871_/C _16868_/X vssd1 vssd1 vccd1 vccd1 _16869_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09410_ _09410_/A vssd1 vssd1 vccd1 vccd1 _10873_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_53_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18608_ _19297_/CLK _18608_/D vssd1 vssd1 vccd1 vccd1 _18608_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19588_ _19594_/CLK _19588_/D vssd1 vssd1 vccd1 vccd1 _19588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09341_ _09341_/A vssd1 vssd1 vccd1 vccd1 _18107_/A sky130_fd_sc_hd__buf_4
XFILLER_80_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18539_ _19292_/CLK _18539_/D vssd1 vssd1 vccd1 vccd1 _18539_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16906__A _16914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09272_ _16622_/A _12602_/B vssd1 vssd1 vccd1 vccd1 _12817_/A sky130_fd_sc_hd__nor2_1
XFILLER_20_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_174_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15691__S _15693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17035__A1 _13418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09608_ _09608_/A vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ _11248_/A vssd1 vssd1 vccd1 vccd1 _11138_/A sky130_fd_sc_hd__buf_2
XFILLER_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09539_ _09539_/A vssd1 vssd1 vccd1 vccd1 _10479_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_19_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ _12542_/X _12544_/X _12547_/Y _12549_/X hold8/X vssd1 vssd1 vccd1 vccd1 _12550_/X
+ sky130_fd_sc_hd__a32o_4
XFILLER_12_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11501_ _12720_/A vssd1 vssd1 vccd1 vccd1 _17981_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_156_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12481_ _17105_/A vssd1 vssd1 vccd1 vccd1 _12482_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_156_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _18618_/Q _13978_/X _14220_/S vssd1 vssd1 vccd1 vccd1 _14221_/A sky130_fd_sc_hd__mux2_1
X_11432_ _11435_/A _11437_/A _11435_/C _10182_/A vssd1 vssd1 vccd1 vccd1 _11432_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_165_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14151_ _14151_/A vssd1 vssd1 vccd1 vccd1 _18587_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14770__S _14770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11363_ _19201_/Q _18815_/Q _19265_/Q _18384_/Q _09704_/X _09733_/X vssd1 vssd1 vccd1
+ vccd1 _11364_/B sky130_fd_sc_hd__mux4_1
XFILLER_164_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_152_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13102_ _19603_/Q _12697_/X _12503_/A _19471_/Q _13101_/X vssd1 vssd1 vccd1 vccd1
+ _15546_/B sky130_fd_sc_hd__a221o_2
X_10314_ _10314_/A _10314_/B vssd1 vssd1 vccd1 vccd1 _10314_/X sky130_fd_sc_hd__and2_1
X_14082_ _14082_/A vssd1 vssd1 vccd1 vccd1 _18557_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11294_ _11462_/B _11461_/A _11461_/B vssd1 vssd1 vccd1 vccd1 _11459_/B sky130_fd_sc_hd__nand3_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17910_ _17910_/A _17910_/B vssd1 vssd1 vccd1 vccd1 _17910_/Y sky130_fd_sc_hd__nand2_1
X_13033_ _13033_/A vssd1 vssd1 vccd1 vccd1 _13234_/A sky130_fd_sc_hd__clkbuf_2
X_10245_ _09844_/A _10231_/X _10235_/X _10244_/X _09670_/A vssd1 vssd1 vccd1 vccd1
+ _10245_/X sky130_fd_sc_hd__a311o_4
XFILLER_65_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18890_ _19311_/CLK _18890_/D vssd1 vssd1 vccd1 vccd1 _18890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10176_ _10158_/A _10175_/X _09909_/X vssd1 vssd1 vccd1 vccd1 _10176_/Y sky130_fd_sc_hd__o21ai_1
X_17841_ _19730_/Q _17831_/X _17840_/X vssd1 vssd1 vccd1 vccd1 _19730_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_51_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output146_A _16272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17772_ _17571_/X _17721_/Y _17771_/Y _17592_/X vssd1 vssd1 vccd1 vccd1 _17772_/X
+ sky130_fd_sc_hd__o211a_1
X_14984_ _18938_/Q vssd1 vssd1 vccd1 vccd1 _14985_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17026__A1 _16935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19511_ _19543_/CLK _19511_/D vssd1 vssd1 vccd1 vccd1 _19511_/Q sky130_fd_sc_hd__dfxtp_1
X_16723_ _16737_/A _16723_/B _16750_/B vssd1 vssd1 vccd1 vccd1 _19550_/D sky130_fd_sc_hd__nor3_1
X_13935_ _13934_/X _18510_/Q _13935_/S vssd1 vssd1 vccd1 vccd1 _13936_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13415__A _18253_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15106__S _15112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19442_ _19583_/CLK _19442_/D vssd1 vssd1 vccd1 vccd1 _19442_/Q sky130_fd_sc_hd__dfxtp_1
X_16654_ _19528_/Q _16663_/D _16653_/Y vssd1 vssd1 vccd1 vccd1 _19528_/D sky130_fd_sc_hd__o21a_1
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13866_ _13866_/A vssd1 vssd1 vccd1 vccd1 _18488_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15605_ _15605_/A vssd1 vssd1 vccd1 vccd1 _19163_/D sky130_fd_sc_hd__clkbuf_1
X_12817_ _12817_/A vssd1 vssd1 vccd1 vccd1 _12817_/X sky130_fd_sc_hd__buf_2
X_16585_ _16585_/A _16585_/B _16586_/B vssd1 vssd1 vccd1 vccd1 _19509_/D sky130_fd_sc_hd__nor3_1
X_19373_ _19373_/CLK _19373_/D vssd1 vssd1 vccd1 vccd1 _19373_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13797_ _13797_/A vssd1 vssd1 vccd1 vccd1 _18462_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17329__A2 _17328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16726__A _16762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15536_ _15519_/X _15534_/X _15535_/Y _15508_/X hold11/X vssd1 vssd1 vccd1 vccd1
+ _15536_/X sky130_fd_sc_hd__a32o_4
X_18324_ _19237_/CLK _18324_/D vssd1 vssd1 vccd1 vccd1 _18324_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ hold16/A _12744_/X _10749_/B _12747_/X vssd1 vssd1 vccd1 vccd1 _18261_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10821__A1 _09432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18255_ _19786_/CLK _18255_/D vssd1 vssd1 vccd1 vccd1 _18255_/Q sky130_fd_sc_hd__dfxtp_2
X_15467_ _15467_/A vssd1 vssd1 vccd1 vccd1 _19138_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ _13009_/A vssd1 vssd1 vccd1 vccd1 _12680_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_129_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17206_ _17662_/B _12195_/A _17263_/A vssd1 vssd1 vccd1 vccd1 _17206_/X sky130_fd_sc_hd__mux2_1
X_14418_ _14418_/A vssd1 vssd1 vccd1 vccd1 _18697_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18186_ _18190_/A _18186_/B vssd1 vssd1 vccd1 vccd1 _18187_/A sky130_fd_sc_hd__and2_1
X_15398_ _19107_/Q _15009_/X _15400_/S vssd1 vssd1 vccd1 vccd1 _15399_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10493__B _12464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17137_ _12482_/A _17115_/X _17149_/A _17140_/A _12543_/B vssd1 vssd1 vccd1 vccd1
+ _17138_/B sky130_fd_sc_hd__a32o_1
XFILLER_7_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15776__S _15776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14349_ _14349_/A vssd1 vssd1 vccd1 vccd1 _18667_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_17068_ _19681_/Q _12577_/B _17072_/S vssd1 vssd1 vccd1 vccd1 _17069_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16019_ _16018_/X _19333_/Q _16025_/S vssd1 vssd1 vccd1 vccd1 _16020_/A sky130_fd_sc_hd__mux2_1
XFILLER_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10337__B1 _09765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09890_ _09890_/A _09890_/B vssd1 vssd1 vccd1 vccd1 _09890_/Y sky130_fd_sc_hd__nor2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17265__A1 _17709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10014__A _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17017__A1 _15620_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09803__A _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19709_ _19712_/CLK _19709_/D vssd1 vssd1 vccd1 vccd1 _19709_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_26_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10949__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17568__A2 _17328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15540__A hold13/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09324_ _17534_/A vssd1 vssd1 vccd1 vccd1 _11512_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__12262__B1 _17305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09255_ _19826_/Q vssd1 vssd1 vccd1 vccd1 _12494_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10684__A _10684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09186_ _09186_/A _09186_/B _11585_/C _11646_/B vssd1 vssd1 vccd1 vccd1 _11573_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_135_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_162_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19736_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14590__S _14599_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15503__A1 _19145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_177_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _18824_/CLK sky130_fd_sc_hd__clkbuf_16
X_10030_ _18636_/Q _18971_/Q _10030_/S vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__mux2_1
XFILLER_89_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_3_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_100_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19669_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _19784_/Q _11342_/A _12028_/S vssd1 vssd1 vccd1 vccd1 _17218_/A sky130_fd_sc_hd__mux2_2
XFILLER_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13720_ _13720_/A vssd1 vssd1 vccd1 vccd1 _18428_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10932_ _09477_/A _10917_/X _10930_/X _09577_/A _10931_/Y vssd1 vssd1 vccd1 vccd1
+ _12450_/B sky130_fd_sc_hd__o32a_4
XFILLER_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_140_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13651_ _13070_/X _18398_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13652_/A sky130_fd_sc_hd__mux2_1
X_10863_ _18393_/Q _18654_/Q _18553_/Q _18888_/Q _10862_/X _09513_/A vssd1 vssd1 vccd1
+ vccd1 _10863_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16546__A _16546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_115_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19649_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_25_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _12606_/A _12602_/B vssd1 vssd1 vccd1 vccd1 _12603_/A sky130_fd_sc_hd__nor2_1
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11056__A1 _11064_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16370_ _19438_/Q _16371_/C _19439_/Q vssd1 vssd1 vccd1 vccd1 _16372_/B sky130_fd_sc_hd__a21oi_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13582_ _13582_/A vssd1 vssd1 vccd1 vccd1 _18373_/D sky130_fd_sc_hd__clkbuf_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10794_ _10787_/X _10789_/Y _10791_/Y _10793_/Y _09658_/X vssd1 vssd1 vccd1 vccd1
+ _10794_/X sky130_fd_sc_hd__o221a_2
XANTENNA__11193__A2_N _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15321_/A vssd1 vssd1 vccd1 vccd1 _19072_/D sky130_fd_sc_hd__clkbuf_1
X_12533_ _19680_/Q _12601_/A _12532_/X _19344_/Q vssd1 vssd1 vccd1 vccd1 _12533_/X
+ sky130_fd_sc_hd__a22o_1
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10594__A _19721_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _18040_/A vssd1 vssd1 vccd1 vccd1 _18188_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_8_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ _14528_/X _19042_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15253_/A sky130_fd_sc_hd__mux2_1
X_12464_ _12468_/A _12464_/B vssd1 vssd1 vccd1 vccd1 _12464_/Y sky130_fd_sc_hd__nor2_1
XFILLER_138_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ _18610_/Q _13953_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14204_/A sky130_fd_sc_hd__mux2_1
X_11415_ _11415_/A _11420_/A _11468_/B _11414_/Y vssd1 vssd1 vccd1 vccd1 _11415_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_137_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15183_ _15183_/A vssd1 vssd1 vccd1 vccd1 _19011_/D sky130_fd_sc_hd__clkbuf_1
X_12395_ _19660_/Q _12368_/X _12130_/X vssd1 vssd1 vccd1 vccd1 _12395_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14134_ _18580_/Q _13959_/X _14136_/S vssd1 vssd1 vccd1 vccd1 _14135_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17495__A1 _17466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _11453_/A _11453_/B _11453_/C _11344_/Y _11345_/Y vssd1 vssd1 vccd1 vccd1
+ _11452_/B sky130_fd_sc_hd__a41o_1
XFILLER_152_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12308__A1 _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ _14122_/S vssd1 vssd1 vccd1 vccd1 _14074_/S sky130_fd_sc_hd__clkbuf_4
X_18942_ _18974_/CLK _18942_/D vssd1 vssd1 vccd1 vccd1 _18942_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10319__B1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14005__S _14011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11277_ _19266_/Q _19104_/Q _18513_/Q _18283_/Q _11112_/X _10910_/A vssd1 vssd1 vccd1
+ vccd1 _11278_/B sky130_fd_sc_hd__mux4_1
XFILLER_79_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13016_ _16862_/B _12950_/X _12951_/X _16450_/B _13015_/X vssd1 vssd1 vccd1 vccd1
+ _15520_/B sky130_fd_sc_hd__a221o_2
X_10228_ _10413_/S vssd1 vssd1 vccd1 vccd1 _10315_/S sky130_fd_sc_hd__clkbuf_4
X_18873_ _19197_/CLK _18873_/D vssd1 vssd1 vccd1 vccd1 _18873_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17824_ _17820_/B _17819_/B _17419_/A _17823_/Y vssd1 vssd1 vccd1 vccd1 _17824_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10159_ _19288_/Q _19126_/Q _18535_/Q _18305_/Q _09782_/A _09956_/A vssd1 vssd1 vccd1
+ vccd1 _10159_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16220__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09623__A _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11872__B _17195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14967_ _14967_/A vssd1 vssd1 vccd1 vccd1 _18929_/D sky130_fd_sc_hd__clkbuf_1
X_17755_ _17844_/S _17752_/X _17754_/X _17626_/A vssd1 vssd1 vccd1 vccd1 _17755_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10769__A _10769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16706_ _19545_/Q _19544_/Q _16706_/C _16706_/D vssd1 vssd1 vccd1 vccd1 _16715_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__09342__B _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12492__B1 _12548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13918_ _14598_/A vssd1 vssd1 vccd1 vccd1 _13918_/X sky130_fd_sc_hd__clkbuf_2
X_14898_ _18896_/Q _14001_/X _14904_/S vssd1 vssd1 vccd1 vccd1 _14899_/A sky130_fd_sc_hd__mux2_1
X_17686_ _17684_/Y _17685_/X _17739_/S vssd1 vssd1 vccd1 vccd1 _17687_/B sky130_fd_sc_hd__mux2_1
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19425_ _19694_/CLK _19425_/D vssd1 vssd1 vccd1 vccd1 _19425_/Q sky130_fd_sc_hd__dfxtp_1
X_16637_ _19523_/Q _19522_/Q _16659_/A _16659_/B vssd1 vssd1 vccd1 vccd1 _16650_/C
+ sky130_fd_sc_hd__and4_1
X_13849_ _13848_/X _18483_/Q _13855_/S vssd1 vssd1 vccd1 vccd1 _13850_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19356_ _19356_/CLK _19356_/D vssd1 vssd1 vccd1 vccd1 _19356_/Q sky130_fd_sc_hd__dfxtp_1
X_16568_ _16585_/A _16568_/B _16569_/B vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__nor3_1
X_18307_ _19096_/CLK _18307_/D vssd1 vssd1 vccd1 vccd1 _18307_/Q sky130_fd_sc_hd__dfxtp_1
X_15519_ _15565_/A vssd1 vssd1 vccd1 vccd1 _15519_/X sky130_fd_sc_hd__clkbuf_2
X_16499_ _16501_/B _16501_/C _16489_/X vssd1 vssd1 vccd1 vccd1 _16499_/Y sky130_fd_sc_hd__a21oi_1
X_19287_ _19287_/CLK _19287_/D vssd1 vssd1 vccd1 vccd1 _19287_/Q sky130_fd_sc_hd__dfxtp_1
X_18238_ input54/X _14274_/X _18229_/X _18234_/X _18140_/A vssd1 vssd1 vccd1 vccd1
+ _18239_/B sky130_fd_sc_hd__a32o_1
XFILLER_163_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09948__C1 _09754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18169_ input62/X _18155_/X _18168_/X _12657_/X _18083_/A vssd1 vssd1 vccd1 vccd1
+ _18170_/B sky130_fd_sc_hd__a32o_1
XFILLER_8_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10009__A _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_94_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19524_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_144_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11539__S _11539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09942_ _19194_/Q _18808_/Q _19258_/Q _18377_/Q _09840_/S _10090_/A vssd1 vssd1 vccd1
+ vccd1 _09943_/B sky130_fd_sc_hd__mux4_1
XANTENNA__17238__A1 _12358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10405__S0 _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09873_ _19291_/Q _19129_/Q _18538_/Q _18308_/Q _09931_/S _09871_/A vssd1 vssd1 vccd1
+ vccd1 _09874_/B sky130_fd_sc_hd__mux4_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13754__S _13758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10708__S1 _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_32_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _18902_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11286__B2 _12445_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11286__A1_N _11070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09307_ _09305_/B _09303_/Y _13166_/A vssd1 vssd1 vccd1 vccd1 _11699_/A sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_47_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _18964_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_10_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09238_ _11560_/B _18083_/A _09172_/C vssd1 vssd1 vccd1 vccd1 _11755_/A sky130_fd_sc_hd__or3b_4
XFILLER_10_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09939__C1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13929__S _13935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ _17168_/A _09169_/B _09169_/C _09168_/X vssd1 vssd1 vccd1 vccd1 _11511_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_163_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ _18578_/Q _18849_/Q _19073_/Q _18817_/Q _11128_/S _10801_/A vssd1 vssd1 vccd1
+ vccd1 _11200_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09708__A _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ _19348_/Q _12068_/A _13411_/A vssd1 vssd1 vccd1 vccd1 _12180_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_107_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_163_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ _18579_/Q _18850_/Q _19074_/Q _18818_/Q _10878_/A _10817_/A vssd1 vssd1 vccd1
+ vccd1 _11131_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_107_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12134__A _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11062_ _11188_/A _11061_/X _11007_/X vssd1 vssd1 vccd1 vccd1 _11062_/X sky130_fd_sc_hd__o21a_1
XFILLER_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13664__S _13664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ _18938_/Q _18704_/Q _19386_/Q _19034_/Q _09539_/A _09547_/X vssd1 vssd1 vccd1
+ vccd1 _10014_/B sky130_fd_sc_hd__mux4_1
X_15870_ _19272_/Q _14541_/A _15876_/S vssd1 vssd1 vccd1 vccd1 _15871_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input22_A io_dbus_rdata[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _18862_/Q _13994_/X _14821_/S vssd1 vssd1 vccd1 vccd1 _14822_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14752_ _14752_/A vssd1 vssd1 vccd1 vccd1 _18831_/D sky130_fd_sc_hd__clkbuf_1
X_17540_ _17468_/A _17533_/X _17539_/X vssd1 vssd1 vccd1 vccd1 _17540_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_151_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11964_ _19643_/Q vssd1 vssd1 vccd1 vccd1 _16974_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09565__S1 _09768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13703_ _12886_/X _18421_/Q _13703_/S vssd1 vssd1 vccd1 vccd1 _13704_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10915_ _11042_/A vssd1 vssd1 vccd1 vccd1 _10915_/X sky130_fd_sc_hd__clkbuf_2
X_17471_ _17471_/A _17471_/B vssd1 vssd1 vccd1 vccd1 _17860_/A sky130_fd_sc_hd__and2_1
XFILLER_60_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11372__S1 _09715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14683_ _14576_/X _18801_/Q _14687_/S vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11895_ _17662_/A _11895_/B vssd1 vssd1 vccd1 vccd1 _11899_/A sky130_fd_sc_hd__xnor2_1
XFILLER_60_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19210_ _19243_/CLK _19210_/D vssd1 vssd1 vccd1 vccd1 _19210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16422_ _16423_/A _16423_/B _16421_/Y vssd1 vssd1 vccd1 vccd1 _19457_/D sky130_fd_sc_hd__o21a_1
X_13634_ _12907_/X _18390_/Q _13642_/S vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__mux2_1
X_10846_ _10839_/Y _10841_/Y _10843_/Y _10845_/Y _09571_/A vssd1 vssd1 vccd1 vccd1
+ _10846_/X sky130_fd_sc_hd__o221a_2
XFILLER_158_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19141_ _19635_/CLK _19141_/D vssd1 vssd1 vccd1 vccd1 _19141_/Q sky130_fd_sc_hd__dfxtp_1
X_16353_ _16589_/A vssd1 vssd1 vccd1 vccd1 _16868_/A sky130_fd_sc_hd__buf_2
X_13565_ _18368_/Q _13563_/X _13577_/S vssd1 vssd1 vccd1 vccd1 _13566_/A sky130_fd_sc_hd__mux2_1
X_10777_ _09632_/A _10776_/X _09563_/A vssd1 vssd1 vccd1 vccd1 _10777_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12309__A _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ _15304_/A vssd1 vssd1 vccd1 vccd1 _19065_/D sky130_fd_sc_hd__clkbuf_1
X_12516_ _12606_/A _12536_/B vssd1 vssd1 vccd1 vccd1 _13055_/A sky130_fd_sc_hd__nor2_2
XFILLER_9_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19072_ _19267_/CLK _19072_/D vssd1 vssd1 vccd1 vccd1 _19072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_157_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16284_ _12126_/A _16278_/X _12129_/X _12135_/X _16280_/X vssd1 vssd1 vccd1 vccd1
+ _19410_/D sky130_fd_sc_hd__o221a_1
XFILLER_158_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17819__B _17819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13496_ _13496_/A vssd1 vssd1 vccd1 vccd1 _18346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_157_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_145_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15235_ _19035_/Q _15086_/X _15239_/S vssd1 vssd1 vccd1 vccd1 _15236_/A sky130_fd_sc_hd__mux2_1
X_18023_ _19783_/Q _11969_/C _18027_/S vssd1 vssd1 vccd1 vccd1 _18024_/A sky130_fd_sc_hd__mux2_1
X_12447_ _12447_/A _12447_/B vssd1 vssd1 vccd1 vccd1 _12447_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output90_A _12337_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15166_ _15166_/A vssd1 vssd1 vccd1 vccd1 _19004_/D sky130_fd_sc_hd__clkbuf_1
X_12378_ _12301_/X _12479_/B _12377_/Y vssd1 vssd1 vccd1 vccd1 _17899_/A sky130_fd_sc_hd__o21ai_4
XFILLER_141_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14117_ _14117_/A vssd1 vssd1 vccd1 vccd1 _18573_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11322_/X _11324_/Y _11326_/Y _11328_/Y _09658_/X vssd1 vssd1 vccd1 vccd1
+ _11329_/X sky130_fd_sc_hd__o221a_2
XANTENNA__09337__B _18144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15097_ _15097_/A vssd1 vssd1 vccd1 vccd1 _18974_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_119_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18925_ _19373_/CLK _18925_/D vssd1 vssd1 vccd1 vccd1 _18925_/Q sky130_fd_sc_hd__dfxtp_1
X_14048_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14048_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_141_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13574__S _13577_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17046__S _17050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18856_ _19081_/CLK _18856_/D vssd1 vssd1 vccd1 vccd1 _18856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17807_ _12174_/A _17737_/X _17806_/X _17761_/X vssd1 vssd1 vccd1 vccd1 _17807_/X
+ sky130_fd_sc_hd__o211a_4
X_18787_ _19237_/CLK _18787_/D vssd1 vssd1 vccd1 vccd1 _18787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15999_ _12071_/X _15998_/Y _13419_/B vssd1 vssd1 vccd1 vccd1 _15999_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17570__A _17831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17738_ _17614_/Y _17610_/Y _17738_/S vssd1 vssd1 vccd1 vccd1 _17738_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09556__S1 _09768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17669_ _17646_/X _17656_/X _17668_/X _17386_/X vssd1 vssd1 vccd1 vccd1 _17669_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15403__A0 _19109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19408_ _19802_/CLK _19408_/D vssd1 vssd1 vccd1 vccd1 _19408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11115__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19339_ _19356_/CLK _19339_/D vssd1 vssd1 vccd1 vccd1 _19339_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_leaf_173_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17156__B1 _17140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16914__A _16914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12219__A _12219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18105__C1 _18097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10626__S0 _10022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15964__S _15970_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_105_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09925_ _09762_/X _09912_/X _09923_/X _09835_/X _09924_/Y vssd1 vssd1 vccd1 vccd1
+ _12474_/B sky130_fd_sc_hd__o32a_4
XFILLER_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13484__S _13492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09856_ _10184_/A _09856_/B vssd1 vssd1 vccd1 vccd1 _09856_/X sky130_fd_sc_hd__or2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_98_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _18637_/Q _18972_/Q _11387_/A vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__mux2_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11259__A1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13513__A _19701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15204__S _15206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _09829_/A _10687_/X _10699_/X vssd1 vssd1 vccd1 vccd1 _10700_/X sky130_fd_sc_hd__a21o_2
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _11730_/A _17237_/A vssd1 vssd1 vccd1 vccd1 _11683_/A sky130_fd_sc_hd__xor2_4
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11106__S1 _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10631_ _18493_/Q _18988_/Q _10631_/S vssd1 vssd1 vccd1 vccd1 _10632_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11033__A _11033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ _13349_/X _18312_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _13351_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10562_ _10617_/A _10562_/B vssd1 vssd1 vccd1 vccd1 _10562_/X sky130_fd_sc_hd__or2_1
XFILLER_155_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12301_ _12301_/A vssd1 vssd1 vccd1 vccd1 _12301_/X sky130_fd_sc_hd__buf_4
XFILLER_139_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13281_ _16142_/A _13281_/B vssd1 vssd1 vccd1 vccd1 _13281_/Y sky130_fd_sc_hd__nor2_1
X_10493_ _10494_/A _12464_/B vssd1 vssd1 vccd1 vccd1 _10495_/A sky130_fd_sc_hd__and2_1
X_15020_ _18950_/Q _15019_/X _15029_/S vssd1 vssd1 vccd1 vccd1 _15021_/A sky130_fd_sc_hd__mux2_1
X_12232_ _11794_/X _12225_/Y _12229_/X _12231_/Y vssd1 vssd1 vccd1 vccd1 _12232_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09438__A _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12163_ _12142_/A _12141_/B _12241_/A vssd1 vssd1 vccd1 vccd1 _12164_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__09157__B _18102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11114_ _11116_/A _11113_/X _11022_/X vssd1 vssd1 vccd1 vccd1 _11114_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16971_ _19642_/Q _16971_/B vssd1 vssd1 vccd1 vccd1 _16971_/X sky130_fd_sc_hd__or2_1
XFILLER_110_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12094_ _19409_/Q _12176_/B vssd1 vssd1 vccd1 vccd1 _12099_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18710_ _19268_/CLK _18710_/D vssd1 vssd1 vccd1 vccd1 _18710_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15175__A _15243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ _19712_/Q vssd1 vssd1 vccd1 vccd1 _11045_/Y sky130_fd_sc_hd__inv_2
X_15922_ _19296_/Q _14617_/A _15924_/S vssd1 vssd1 vccd1 vccd1 _15923_/A sky130_fd_sc_hd__mux2_1
XFILLER_89_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19690_ _19693_/CLK _19690_/D vssd1 vssd1 vccd1 vccd1 _19690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_103_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18641_ _19711_/CLK _18641_/D vssd1 vssd1 vccd1 vccd1 _18641_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_162_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15853_ _15853_/A vssd1 vssd1 vccd1 vccd1 _19265_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10170__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_0_0_clock clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA__11208__A _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ _18854_/Q _13969_/X _14810_/S vssd1 vssd1 vccd1 vccd1 _14805_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18572_ _19035_/CLK _18572_/D vssd1 vssd1 vccd1 vccd1 _18572_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15784_ _15852_/S vssd1 vssd1 vccd1 vccd1 _15793_/S sky130_fd_sc_hd__clkbuf_4
X_12996_ _13154_/A _12992_/X _12994_/Y _12995_/X _13164_/A vssd1 vssd1 vccd1 vccd1
+ _12997_/B sky130_fd_sc_hd__a221o_1
XFILLER_80_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17523_ _17481_/X _17522_/X _17577_/S vssd1 vssd1 vccd1 vccd1 _17674_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14735_ _14547_/X _18824_/Q _14737_/S vssd1 vssd1 vccd1 vccd1 _14736_/A sky130_fd_sc_hd__mux2_1
X_11947_ _12020_/A _12459_/A _11946_/Y vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__a21oi_1
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17925__A2 _17430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _17444_/Y _17452_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17454_/X sky130_fd_sc_hd__mux2_1
X_14666_ _14666_/A vssd1 vssd1 vccd1 vccd1 _18793_/D sky130_fd_sc_hd__clkbuf_1
X_11878_ _11879_/A _11879_/C _19401_/Q vssd1 vssd1 vccd1 vccd1 _11880_/A sky130_fd_sc_hd__a21oi_1
X_16405_ _19450_/Q _16406_/C _19451_/Q vssd1 vssd1 vccd1 vccd1 _16407_/B sky130_fd_sc_hd__a21oi_1
X_13617_ _14297_/B vssd1 vssd1 vccd1 vccd1 _14787_/B sky130_fd_sc_hd__buf_6
XFILLER_20_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10829_ _18393_/Q _18654_/Q _18553_/Q _18888_/Q _11049_/S _10817_/X vssd1 vssd1 vccd1
+ vccd1 _10830_/B sky130_fd_sc_hd__mux4_1
X_14597_ _14597_/A vssd1 vssd1 vccd1 vccd1 _18770_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17385_ _17471_/A _17471_/B vssd1 vssd1 vccd1 vccd1 _17386_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12039__A _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19124_ _19124_/CLK _19124_/D vssd1 vssd1 vccd1 vccd1 _19124_/Q sky130_fd_sc_hd__dfxtp_1
X_16336_ _19428_/Q _16332_/C _16335_/Y vssd1 vssd1 vccd1 vccd1 _19428_/D sky130_fd_sc_hd__o21a_1
X_13548_ _13615_/S vssd1 vssd1 vccd1 vccd1 _13561_/S sky130_fd_sc_hd__buf_2
XFILLER_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16267_ _16267_/A vssd1 vssd1 vccd1 vccd1 _19403_/D sky130_fd_sc_hd__clkbuf_1
X_19055_ _19249_/CLK _19055_/D vssd1 vssd1 vccd1 vccd1 _19055_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10630__C1 _09572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13479_ _13148_/X _18339_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _13480_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15218_ _15218_/A vssd1 vssd1 vccd1 vccd1 _19027_/D sky130_fd_sc_hd__clkbuf_1
X_18006_ _18006_/A vssd1 vssd1 vccd1 vccd1 _19775_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09348__A _19864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16198_ _13554_/X _19372_/Q _16202_/S vssd1 vssd1 vccd1 vccd1 _16199_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11186__B1 _11007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12922__A1 input29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ _15149_/A vssd1 vssd1 vccd1 vccd1 _18996_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09710_ _09710_/A vssd1 vssd1 vccd1 vccd1 _10238_/A sky130_fd_sc_hd__clkbuf_4
X_18908_ _19325_/CLK _18908_/D vssd1 vssd1 vccd1 vccd1 _18908_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12502__A _13356_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09641_ _11331_/A _09639_/X _09640_/X vssd1 vssd1 vccd1 vccd1 _09641_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18839_ _19256_/CLK _18839_/D vssd1 vssd1 vccd1 vccd1 _18839_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15624__A0 _13344_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17504__S _17504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09572_ _09572_/A vssd1 vssd1 vccd1 vccd1 _09829_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10022__A _10631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09811__A _09811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__S1 _10060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17916__A2 _17430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15959__S _15959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10168__S _10168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14863__S _14871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16644__A _16666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13479__S _13481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10924__B1 _09561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11192__A3 _11191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09908_ _18602_/Q _18873_/Q _19097_/Q _18841_/Q _10112_/S _09905_/A vssd1 vssd1 vccd1
+ vccd1 _09908_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10631__S _10631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14103__S _14107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09839_ _09839_/A _09839_/B vssd1 vssd1 vccd1 vccd1 _09839_/X sky130_fd_sc_hd__and2_1
XFILLER_101_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _15006_/A vssd1 vssd1 vccd1 vccd1 _14528_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15723__A _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _19637_/Q _11801_/B vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11327__S1 _10705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12781_/A vssd1 vssd1 vccd1 vccd1 _12781_/X sky130_fd_sc_hd__clkbuf_4
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10867__A _19715_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14520_ _15926_/B _16169_/A vssd1 vssd1 vccd1 vccd1 _14602_/A sky130_fd_sc_hd__nand2_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ _11788_/A _11788_/B vssd1 vssd1 vccd1 vccd1 _11732_/X sky130_fd_sc_hd__xor2_4
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14451_ _14451_/A vssd1 vssd1 vccd1 vccd1 _18711_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _12184_/A vssd1 vssd1 vccd1 vccd1 _12074_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14773__S _14781_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13402_ _15494_/A hold21/A vssd1 vssd1 vccd1 vccd1 _13402_/Y sky130_fd_sc_hd__nand2_1
XFILLER_174_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10614_ _10614_/A _10614_/B vssd1 vssd1 vccd1 vccd1 _10614_/X sky130_fd_sc_hd__or2_1
X_17170_ _17319_/B vssd1 vssd1 vccd1 vccd1 _17404_/B sky130_fd_sc_hd__clkbuf_2
X_14382_ _13851_/X _18681_/Q _14384_/S vssd1 vssd1 vccd1 vccd1 _14383_/A sky130_fd_sc_hd__mux2_1
XFILLER_167_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11594_ _11668_/B vssd1 vssd1 vccd1 vccd1 _17207_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16121_ _16121_/A vssd1 vssd1 vccd1 vccd1 _19350_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13333_ input22/X _13166_/A _13254_/X vssd1 vssd1 vccd1 vccd1 _13333_/X sky130_fd_sc_hd__a21o_1
X_10545_ _18623_/Q _18958_/Q _10602_/S vssd1 vssd1 vccd1 vccd1 _10545_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14354__A0 _13918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16052_ _12651_/X _16051_/Y _16052_/S vssd1 vssd1 vccd1 vccd1 _16052_/X sky130_fd_sc_hd__mux2_1
X_13264_ _19163_/Q _13007_/X _12532_/X _19353_/Q _13263_/X vssd1 vssd1 vccd1 vccd1
+ _13264_/X sky130_fd_sc_hd__a221o_2
XFILLER_108_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10476_ _19314_/Q _18726_/Q _18763_/Q _18337_/Q _10260_/A _10521_/A vssd1 vssd1 vccd1
+ vccd1 _10476_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15003_ _15003_/A vssd1 vssd1 vccd1 vccd1 _15003_/X sky130_fd_sc_hd__buf_2
X_12215_ _12242_/B _12215_/B vssd1 vssd1 vccd1 vccd1 _12220_/A sky130_fd_sc_hd__nor2_1
XFILLER_124_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13195_ _19760_/Q vssd1 vssd1 vccd1 vccd1 _13195_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10066__S1 _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19811_ _19866_/CLK _19811_/D vssd1 vssd1 vccd1 vccd1 _19811_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_97_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12380__A2 _17886_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__and2_1
XFILLER_97_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_121_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13418__A _13418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19742_ _19779_/CLK _19742_/D vssd1 vssd1 vccd1 vccd1 _19742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16954_ _16981_/A vssd1 vssd1 vccd1 vccd1 _16954_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_12077_ _19647_/Q _12105_/C vssd1 vssd1 vccd1 vccd1 _12104_/B sky130_fd_sc_hd__and2_1
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_110_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15905_ _19288_/Q _14592_/A _15909_/S vssd1 vssd1 vccd1 vccd1 _15906_/A sky130_fd_sc_hd__mux2_1
X_11028_ _11111_/A _11027_/X _09481_/A vssd1 vssd1 vccd1 vccd1 _11028_/Y sky130_fd_sc_hd__o21ai_1
X_19673_ _19695_/CLK _19673_/D vssd1 vssd1 vccd1 vccd1 _19673_/Q sky130_fd_sc_hd__dfxtp_1
X_16885_ _16887_/A _16887_/C _16868_/X vssd1 vssd1 vccd1 vccd1 _16885_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18624_ _19088_/CLK _18624_/D vssd1 vssd1 vccd1 vccd1 _18624_/Q sky130_fd_sc_hd__dfxtp_1
X_15836_ _15836_/A vssd1 vssd1 vccd1 vccd1 _19257_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18555_ _19311_/CLK _18555_/D vssd1 vssd1 vccd1 vccd1 _18555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12979_ _11538_/X _12973_/X _12978_/X vssd1 vssd1 vccd1 vccd1 _15025_/A sky130_fd_sc_hd__o21a_2
XFILLER_92_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15767_ _15767_/A vssd1 vssd1 vccd1 vccd1 _15776_/S sky130_fd_sc_hd__buf_4
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17506_ _17509_/S _17506_/B vssd1 vssd1 vccd1 vccd1 _17506_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09350__B _18140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A2 _10432_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14718_ _14519_/X _18816_/Q _14726_/S vssd1 vssd1 vccd1 vccd1 _14719_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16031__A0 _16919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18486_ _18917_/CLK _18486_/D vssd1 vssd1 vccd1 vccd1 _18486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15698_ _14605_/X _19196_/Q _15704_/S vssd1 vssd1 vccd1 vccd1 _15699_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17437_ _17397_/Y _17436_/Y _17572_/S vssd1 vssd1 vccd1 vccd1 _17437_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14683__S _14687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14649_ _14649_/A vssd1 vssd1 vccd1 vccd1 _18785_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_46_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10829__S0 _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17368_ _17368_/A vssd1 vssd1 vccd1 vccd1 _17368_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19107_ _19108_/CLK _19107_/D vssd1 vssd1 vccd1 vccd1 _19107_/Q sky130_fd_sc_hd__dfxtp_1
X_16319_ _16324_/D vssd1 vssd1 vccd1 vccd1 _16504_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_118_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17299_ _17393_/A vssd1 vssd1 vccd1 vccd1 _17550_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_174_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19038_ _19390_/CLK _19038_/D vssd1 vssd1 vccd1 vccd1 _19038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_133_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput101 _11855_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[8] sky130_fd_sc_hd__buf_2
XFILLER_133_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput112 _12459_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[12] sky130_fd_sc_hd__buf_2
XFILLER_133_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput123 _12471_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[22] sky130_fd_sc_hd__buf_2
Xoutput134 _12446_/X vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[3] sky130_fd_sc_hd__buf_2
Xoutput145 _11975_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[12] sky130_fd_sc_hd__buf_2
Xoutput156 _12237_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[22] sky130_fd_sc_hd__buf_2
Xoutput167 _16249_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[3] sky130_fd_sc_hd__buf_2
XFILLER_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11006__S0 _10940_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14858__S _14858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13762__S _13762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09624_ _09624_/A vssd1 vssd1 vccd1 vccd1 _09625_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09555_ _10296_/A _09509_/Y _09528_/X _09550_/Y _09811_/A vssd1 vssd1 vccd1 vccd1
+ _09555_/X sky130_fd_sc_hd__o311a_4
XFILLER_71_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _18643_/Q vssd1 vssd1 vccd1 vccd1 _10968_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_52_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15689__S _15693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14593__S _14599_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10330_ _19189_/Q _18803_/Q _19253_/Q _18372_/Q _10286_/X _10382_/A vssd1 vssd1 vccd1
+ vccd1 _10331_/B sky130_fd_sc_hd__mux4_1
XFILLER_139_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10261_ _10261_/A vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_106_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12000_ _17722_/A _12000_/B vssd1 vssd1 vccd1 vccd1 _12004_/A sky130_fd_sc_hd__xor2_1
XFILLER_132_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10192_ _10195_/A _10189_/X _10191_/X _09740_/A vssd1 vssd1 vccd1 vccd1 _10192_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14639__A1 input44/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14639__B2 _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13951_ _18513_/Q _13943_/X _13963_/S vssd1 vssd1 vccd1 vccd1 _13952_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14768__S _14770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09610__S0 _09599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16549__A _16549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _19712_/Q _15485_/B _13103_/S vssd1 vssd1 vccd1 vccd1 _12902_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16670_ _16696_/A _16670_/B _16679_/D vssd1 vssd1 vccd1 vccd1 _19532_/D sky130_fd_sc_hd__nor3_1
XANTENNA__10220__S1 _09905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13882_ _13882_/A vssd1 vssd1 vccd1 vccd1 _18493_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10676__A2 _10663_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12833_ _19490_/Q vssd1 vssd1 vccd1 vccd1 _16529_/B sky130_fd_sc_hd__clkbuf_2
X_15621_ _19735_/Q _15620_/X _15626_/S vssd1 vssd1 vccd1 vccd1 _15621_/X sky130_fd_sc_hd__mux2_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10597__A _10597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _19378_/CLK _18340_/D vssd1 vssd1 vccd1 vccd1 _18340_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _19722_/Q _15550_/X _15569_/S vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__mux2_1
X_12764_ _18272_/Q _12759_/X _11354_/A _12762_/X vssd1 vssd1 vccd1 vccd1 _18272_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09913__S1 _09905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11723_/S _12445_/B _11674_/X vssd1 vssd1 vccd1 vccd1 _17393_/A sky130_fd_sc_hd__o21ai_2
X_14503_ _13921_/X _18735_/Q _14511_/S vssd1 vssd1 vccd1 vccd1 _14504_/A sky130_fd_sc_hd__mux2_1
X_15483_ _15482_/X _19142_/Q _15483_/S vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__mux2_1
X_18271_ _19162_/CLK _18271_/D vssd1 vssd1 vccd1 vccd1 _18271_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12674_/X _12675_/X _12691_/X _12694_/X vssd1 vssd1 vccd1 vccd1 _19584_/D
+ sky130_fd_sc_hd__o22a_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17222_ _17222_/A vssd1 vssd1 vccd1 vccd1 _17790_/B sky130_fd_sc_hd__buf_2
XFILLER_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14434_ _14434_/A vssd1 vssd1 vccd1 vccd1 _18704_/D sky130_fd_sc_hd__clkbuf_1
X_11646_ _19842_/Q _11646_/B _11646_/C _11569_/B vssd1 vssd1 vccd1 vccd1 _11647_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_156_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 io_dbus_rdata[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
Xinput25 io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_4
X_17153_ _17122_/A _17149_/X _17140_/X _12975_/B vssd1 vssd1 vccd1 vccd1 _17154_/B
+ sky130_fd_sc_hd__a22o_1
X_14365_ _13934_/X _18675_/Q _14365_/S vssd1 vssd1 vccd1 vccd1 _14366_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10287__S1 _10275_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__S _14011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput36 io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
X_11577_ _17166_/B _11577_/B _11577_/C _17183_/B vssd1 vssd1 vccd1 vccd1 _11577_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__09451__C1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput47 io_ibus_inst[21] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_2
XFILLER_116_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput58 io_ibus_inst[31] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_2
XFILLER_116_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16104_ _15574_/X _16103_/Y _16156_/S vssd1 vssd1 vccd1 vccd1 _16104_/X sky130_fd_sc_hd__mux2_1
X_13316_ _16142_/B _13315_/C _19767_/Q vssd1 vssd1 vccd1 vccd1 _13316_/Y sky130_fd_sc_hd__a21oi_1
Xinput69 io_irq_uart_irq vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_1
X_17084_ _17084_/A vssd1 vssd1 vccd1 vccd1 _19688_/D sky130_fd_sc_hd__clkbuf_1
X_10528_ _10535_/A _10527_/X _10297_/A vssd1 vssd1 vccd1 vccd1 _10528_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_170_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14296_ _14296_/A vssd1 vssd1 vccd1 vccd1 _18645_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16731__B _16731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16035_ _16039_/A _16039_/C vssd1 vssd1 vccd1 vccd1 _16035_/Y sky130_fd_sc_hd__xnor2_2
X_13247_ _19731_/Q _12712_/B _13247_/S vssd1 vssd1 vccd1 vccd1 _13247_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10459_ _09727_/A _10449_/X _10453_/X _10458_/X _09669_/A vssd1 vssd1 vccd1 vccd1
+ _10459_/X sky130_fd_sc_hd__a311o_4
XFILLER_171_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17816__A1 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _19540_/Q vssd1 vssd1 vccd1 vccd1 _16697_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_170_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10271__S _10381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _19346_/Q _12069_/X _12128_/X _12075_/X vssd1 vssd1 vccd1 vccd1 _12129_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09345__B _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17986_ _16142_/B _19798_/Q _17990_/S vssd1 vssd1 vccd1 vccd1 _17987_/A sky130_fd_sc_hd__mux2_1
XFILLER_97_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19725_ _19725_/CLK _19725_/D vssd1 vssd1 vccd1 vccd1 _19725_/Q sky130_fd_sc_hd__dfxtp_2
X_16937_ _16937_/A _16937_/B _16937_/C _16937_/D vssd1 vssd1 vccd1 vccd1 _16959_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__10116__A1 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09601__S0 _09599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18241__A1 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19656_ _19693_/CLK _19656_/D vssd1 vssd1 vccd1 vccd1 _19656_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18241__B2 _17125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16868_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16868_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18607_ _19113_/CLK _18607_/D vssd1 vssd1 vccd1 vccd1 _18607_/Q sky130_fd_sc_hd__dfxtp_1
X_15819_ _15819_/A vssd1 vssd1 vccd1 vccd1 _19249_/D sky130_fd_sc_hd__clkbuf_1
X_19587_ _19807_/CLK _19587_/D vssd1 vssd1 vccd1 vccd1 _19587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16799_ _16799_/A _16799_/B _16807_/C vssd1 vssd1 vccd1 vccd1 _19573_/D sky130_fd_sc_hd__nor3_1
XFILLER_18_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09340_ _11574_/A vssd1 vssd1 vccd1 vccd1 _17121_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18538_ _19197_/CLK _18538_/D vssd1 vssd1 vccd1 vccd1 _18538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _12782_/A _13391_/B _12956_/A _09271_/D vssd1 vssd1 vccd1 vccd1 _09271_/X
+ sky130_fd_sc_hd__and4b_1
X_18469_ _19287_/CLK _18469_/D vssd1 vssd1 vccd1 vccd1 _18469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13611__A _15095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__A1 _12035_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12227__A _19414_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11227__S0 _11074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10970__A _18642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17753__A _17753_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13492__S _13492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09607_ _19328_/Q _18740_/Q _18777_/Q _18351_/Q _09599_/X _09977_/A vssd1 vssd1 vccd1
+ vccd1 _09607_/X sky130_fd_sc_hd__mux4_1
XFILLER_113_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09538_ _09538_/A vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__buf_2
XFILLER_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09469_ _09469_/A vssd1 vssd1 vccd1 vccd1 _09470_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12280__A1 _18132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ _11508_/A _11943_/A vssd1 vssd1 vccd1 vccd1 _11557_/D sky130_fd_sc_hd__nand2_4
XFILLER_157_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12480_ _12480_/A _12480_/B vssd1 vssd1 vccd1 vccd1 _12480_/Y sky130_fd_sc_hd__nor2_1
XFILLER_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11431_ _11431_/A _11433_/A _11431_/C vssd1 vssd1 vccd1 vccd1 _11431_/Y sky130_fd_sc_hd__nand3_1
XFILLER_11_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11041__A _11232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14150_ _18587_/Q _13981_/X _14158_/S vssd1 vssd1 vccd1 vccd1 _14151_/A sky130_fd_sc_hd__mux2_1
X_11362_ _11416_/A _12478_/B _11415_/A vssd1 vssd1 vccd1 vccd1 _11362_/X sky130_fd_sc_hd__or3_1
X_13101_ _19535_/Q _12939_/S _12953_/A _19503_/Q _13100_/X vssd1 vssd1 vccd1 vccd1
+ _13101_/X sky130_fd_sc_hd__a221o_1
XFILLER_125_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10313_ _18628_/Q _18963_/Q _10315_/S vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__mux2_1
XANTENNA__13667__S _13675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14081_ _13880_/X _18557_/Q _14085_/S vssd1 vssd1 vccd1 vccd1 _14082_/A sky130_fd_sc_hd__mux2_1
X_11293_ _11463_/A _11463_/B _11463_/C vssd1 vssd1 vccd1 vccd1 _11461_/B sky130_fd_sc_hd__a21o_1
XFILLER_4_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13032_ _19718_/Q _12649_/B _13345_/S vssd1 vssd1 vccd1 vccd1 _13032_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input52_A io_ibus_inst[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _10237_/X _10239_/X _10242_/X _10243_/X vssd1 vssd1 vccd1 vccd1 _10244_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09446__A _18782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17840_ _12252_/Y _17786_/X _17839_/X _17795_/X vssd1 vssd1 vccd1 vccd1 _17840_/X
+ sky130_fd_sc_hd__a211o_1
X_10175_ _18599_/Q _18870_/Q _19094_/Q _18838_/Q _10114_/S _09956_/A vssd1 vssd1 vccd1
+ vccd1 _10175_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17771_ _17771_/A _17771_/B vssd1 vssd1 vccd1 vccd1 _17771_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14498__S _14500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14983_ _14983_/A vssd1 vssd1 vccd1 vccd1 _18937_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16279__A _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19510_ _19540_/CLK _19510_/D vssd1 vssd1 vccd1 vccd1 _19510_/Q sky130_fd_sc_hd__dfxtp_1
X_16722_ _19550_/Q _19549_/Q _19548_/Q _16722_/D vssd1 vssd1 vccd1 vccd1 _16750_/B
+ sky130_fd_sc_hd__and4_2
X_13934_ _14614_/A vssd1 vssd1 vccd1 vccd1 _13934_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_93_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19441_ _19448_/CLK _19441_/D vssd1 vssd1 vccd1 vccd1 _19441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16653_ _16666_/A _16655_/B vssd1 vssd1 vccd1 vccd1 _16653_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13415__B _13415_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13865_ _13864_/X _18488_/Q _13871_/S vssd1 vssd1 vccd1 vccd1 _13866_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15604_ _15602_/X _19163_/Q _15627_/S vssd1 vssd1 vccd1 vccd1 _15605_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15911__A _15911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ _19457_/Q vssd1 vssd1 vccd1 vccd1 _16423_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19372_ _19374_/CLK _19372_/D vssd1 vssd1 vccd1 vccd1 _19372_/Q sky130_fd_sc_hd__dfxtp_1
X_16584_ _19509_/Q _19508_/Q _16584_/C vssd1 vssd1 vccd1 vccd1 _16586_/B sky130_fd_sc_hd__and3_1
XFILLER_90_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13796_ _13070_/X _18462_/Q _13798_/S vssd1 vssd1 vccd1 vccd1 _13797_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18323_ _19300_/CLK _18323_/D vssd1 vssd1 vccd1 vccd1 _18323_/Q sky130_fd_sc_hd__dfxtp_1
X_15535_ _15541_/A hold11/A vssd1 vssd1 vccd1 vccd1 _15535_/Y sky130_fd_sc_hd__nand2_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16537__A1 _16540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12747_/A vssd1 vssd1 vccd1 vccd1 _12747_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16218__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10282__B1 _09764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18254_ _19786_/CLK _18254_/D vssd1 vssd1 vccd1 vccd1 _18254_/Q sky130_fd_sc_hd__dfxtp_1
X_15466_ _15461_/X _19138_/Q _15483_/S vssd1 vssd1 vccd1 vccd1 _15467_/A sky130_fd_sc_hd__mux2_1
X_12678_ _19161_/Q _13179_/A _12677_/X _19351_/Q vssd1 vssd1 vccd1 vccd1 _12678_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_129_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17205_ _17205_/A vssd1 vssd1 vccd1 vccd1 _17662_/B sky130_fd_sc_hd__clkbuf_2
X_14417_ _13902_/X _18697_/Q _14417_/S vssd1 vssd1 vccd1 vccd1 _14418_/A sky130_fd_sc_hd__mux2_1
X_11629_ _19852_/Q vssd1 vssd1 vccd1 vccd1 _18112_/A sky130_fd_sc_hd__buf_4
XFILLER_8_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12023__A1 _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18185_ input35/X _18178_/X _18168_/X _18174_/X _19845_/Q vssd1 vssd1 vccd1 vccd1
+ _18186_/B sky130_fd_sc_hd__a32o_1
XFILLER_128_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16742__A _16762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15397_ _15397_/A vssd1 vssd1 vccd1 vccd1 _19106_/D sky130_fd_sc_hd__clkbuf_1
X_17136_ _17136_/A vssd1 vssd1 vccd1 vccd1 _19698_/D sky130_fd_sc_hd__clkbuf_1
X_14348_ _13909_/X _18667_/Q _14354_/S vssd1 vssd1 vccd1 vccd1 _14349_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13577__S _13577_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11209__S0 _11128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17067_ _17067_/A vssd1 vssd1 vccd1 vccd1 _19680_/D sky130_fd_sc_hd__clkbuf_1
X_14279_ input46/X _14274_/X _14277_/X _14278_/X _09351_/A vssd1 vssd1 vccd1 vccd1
+ _18216_/B sky130_fd_sc_hd__a32o_2
XFILLER_144_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13118__A4 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13523__A1 _13522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16018_ _15487_/X _16017_/Y _16024_/S vssd1 vssd1 vccd1 vccd1 _16018_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10337__A1 _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17670__C1 _17831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _17969_/A vssd1 vssd1 vccd1 vccd1 _19758_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_84_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19708_ _19740_/CLK _19708_/D vssd1 vssd1 vccd1 vccd1 _19708_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11837__A1 _19399_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14201__S _14209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10196__S0 _09854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19639_ _19645_/CLK _19639_/D vssd1 vssd1 vccd1 vccd1 _19639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11126__A _11138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09889__S0 _10114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ _17753_/A vssd1 vssd1 vccd1 vccd1 _17534_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10965__A _10965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09254_ _09270_/B vssd1 vssd1 vccd1 vccd1 _12602_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_166_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14871__S _14871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ _09185_/A _11574_/A _11560_/B vssd1 vssd1 vccd1 vccd1 _11573_/A sky130_fd_sc_hd__or3_2
XFILLER_119_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09966__B1 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11796__A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10328__A1 _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_168_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_124_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13516__A _13615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11828__A1 _11824_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11980_ _17709_/A _11980_/B vssd1 vssd1 vccd1 vccd1 _11984_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10931_ _19714_/Q vssd1 vssd1 vccd1 vccd1 _10931_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13650_ _13650_/A vssd1 vssd1 vccd1 vccd1 _18397_/D sky130_fd_sc_hd__clkbuf_1
X_10862_ _11071_/S vssd1 vssd1 vccd1 vccd1 _10862_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ _12601_/A vssd1 vssd1 vccd1 vccd1 _17028_/A sky130_fd_sc_hd__buf_2
XFILLER_25_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13581_ _18373_/Q _13579_/X _13593_/S vssd1 vssd1 vccd1 vccd1 _13582_/A sky130_fd_sc_hd__mux2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10875__A _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10793_ _11335_/A _10792_/X _09484_/A vssd1 vssd1 vccd1 vccd1 _10793_/Y sky130_fd_sc_hd__o21ai_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _12958_/A vssd1 vssd1 vccd1 vccd1 _12532_/X sky130_fd_sc_hd__clkbuf_2
X_15320_ _19072_/Q _14996_/X _15328_/S vssd1 vssd1 vccd1 vccd1 _15321_/A sky130_fd_sc_hd__mux2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15251_ _15251_/A vssd1 vssd1 vccd1 vccd1 _19041_/D sky130_fd_sc_hd__clkbuf_1
X_12463_ _12475_/A vssd1 vssd1 vccd1 vccd1 _12468_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14781__S _14781_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14202_ _14202_/A vssd1 vssd1 vccd1 vccd1 _18609_/D sky130_fd_sc_hd__clkbuf_1
X_11414_ _11416_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _11414_/Y sky130_fd_sc_hd__nor2_1
X_15182_ _19011_/Q _15009_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15183_/A sky130_fd_sc_hd__mux2_1
X_12394_ _19660_/Q _19659_/Q _12394_/C vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__and3_1
XFILLER_126_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14133_ _14133_/A vssd1 vssd1 vccd1 vccd1 _18579_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11345_ _11342_/Y _10649_/A _11343_/A vssd1 vssd1 vccd1 vccd1 _11345_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_99_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _14064_/A vssd1 vssd1 vccd1 vccd1 _18549_/D sky130_fd_sc_hd__clkbuf_1
X_18941_ _19389_/CLK _18941_/D vssd1 vssd1 vccd1 vccd1 _18941_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10319__A1 _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11276_ _09531_/A _11275_/X _11022_/X vssd1 vssd1 vccd1 vccd1 _11276_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_141_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13015_ _19530_/Q _13004_/X _12953_/X _19498_/Q _13014_/X vssd1 vssd1 vccd1 vccd1
+ _13015_/X sky130_fd_sc_hd__a221o_2
X_10227_ _11354_/A _12470_/B vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__or2_1
X_18872_ _19096_/CLK _18872_/D vssd1 vssd1 vccd1 vccd1 _18872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10115__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17823_ _17920_/B _17823_/B vssd1 vssd1 vccd1 vccd1 _17823_/Y sky130_fd_sc_hd__nand2_1
X_10158_ _10158_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10158_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA__14021__S _14027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17754_ _17753_/A _12089_/X _17462_/A _17753_/Y vssd1 vssd1 vccd1 vccd1 _17754_/X
+ sky130_fd_sc_hd__o211a_1
X_14966_ _18929_/Q vssd1 vssd1 vccd1 vccd1 _14967_/A sky130_fd_sc_hd__clkbuf_1
X_10089_ _10089_/A _11431_/A vssd1 vssd1 vccd1 vccd1 _11423_/A sky130_fd_sc_hd__or2b_1
XFILLER_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16705_ _16737_/A _16705_/B _16712_/D vssd1 vssd1 vccd1 vccd1 _19544_/D sky130_fd_sc_hd__nor3_1
XFILLER_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13917_ _13917_/A vssd1 vssd1 vccd1 vccd1 _18504_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12492__A1 _12543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17685_ _17514_/B _17500_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17685_/X sky130_fd_sc_hd__mux2_1
XANTENNA__16737__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14897_ _14897_/A vssd1 vssd1 vccd1 vccd1 _18895_/D sky130_fd_sc_hd__clkbuf_1
X_19424_ _19694_/CLK _19424_/D vssd1 vssd1 vccd1 vccd1 _19424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16636_ _19522_/Q _16633_/C _16635_/Y vssd1 vssd1 vccd1 vccd1 _19522_/D sky130_fd_sc_hd__o21a_1
X_13848_ _14528_/A vssd1 vssd1 vccd1 vccd1 _13848_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19355_ _19357_/CLK _19355_/D vssd1 vssd1 vccd1 vccd1 _19355_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12244__A1 _11357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ _19503_/Q hold1/X _16567_/C vssd1 vssd1 vccd1 vccd1 _16569_/B sky130_fd_sc_hd__and3_1
X_13779_ _12907_/X _18454_/Q _13787_/S vssd1 vssd1 vccd1 vccd1 _13780_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18306_ _19127_/CLK _18306_/D vssd1 vssd1 vccd1 vccd1 _18306_/Q sky130_fd_sc_hd__dfxtp_1
X_15518_ _15518_/A vssd1 vssd1 vccd1 vccd1 _19147_/D sky130_fd_sc_hd__clkbuf_1
X_19286_ _19286_/CLK _19286_/D vssd1 vssd1 vccd1 vccd1 _19286_/Q sky130_fd_sc_hd__dfxtp_1
X_16498_ _19483_/Q _16495_/B _16497_/Y vssd1 vssd1 vccd1 vccd1 _19483_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15787__S _15793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18237_ _18237_/A vssd1 vssd1 vccd1 vccd1 _19862_/D sky130_fd_sc_hd__clkbuf_1
X_15449_ _19130_/Q _15083_/X _15455_/S vssd1 vssd1 vccd1 vccd1 _15450_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16930__A1 _19628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__B1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18168_ _18188_/A vssd1 vssd1 vccd1 vccd1 _18168_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10102__S0 _10093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _17114_/A _17120_/D _17115_/X _17907_/A _17118_/X vssd1 vssd1 vccd1 vccd1
+ _17119_/X sky130_fd_sc_hd__a311o_1
XFILLER_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18099_ _18099_/A vssd1 vssd1 vccd1 vccd1 _18128_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_117_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15497__A1 _19144_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09941_ _09941_/A _09941_/B vssd1 vssd1 vccd1 vccd1 _09941_/X sky130_fd_sc_hd__or2_1
XFILLER_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10405__S1 _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09872_ _18474_/Q _19065_/Q _19227_/Q _18442_/Q _09930_/S _09871_/X vssd1 vssd1 vccd1
+ vccd1 _09872_/X sky130_fd_sc_hd__mux4_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15535__B hold11/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13770__S _13776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15551__A _15601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09306_ _09306_/A vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__buf_2
XANTENNA__12786__A2 _12603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09237_ _11569_/A _11569_/B vssd1 vssd1 vccd1 vccd1 _11943_/A sky130_fd_sc_hd__nand2_4
XFILLER_166_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_94_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09168_ _09328_/A _11566_/C _09208_/A _17165_/B _17165_/A vssd1 vssd1 vccd1 vccd1
+ _09168_/X sky130_fd_sc_hd__o32a_2
XANTENNA__10549__A1 _10310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09099_ _19836_/Q vssd1 vssd1 vccd1 vccd1 _09236_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11130_ _09416_/A _11127_/X _11129_/X vssd1 vssd1 vccd1 vccd1 _11130_/X sky130_fd_sc_hd__a21o_1
XFILLER_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_134_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11061_ _19302_/Q _18714_/Q _18751_/Q _18325_/Q _11011_/X _11012_/X vssd1 vssd1 vccd1
+ vccd1 _11061_/X sky130_fd_sc_hd__mux4_1
XFILLER_62_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18102__A _18102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14630__A _14630_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10012_ _10004_/Y _10007_/Y _10009_/Y _10011_/Y _09829_/A vssd1 vssd1 vccd1 vccd1
+ _10012_/X sky130_fd_sc_hd__o221a_4
XFILLER_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16988__A1 _12577_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820_ _14820_/A vssd1 vssd1 vccd1 vccd1 _18861_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_92_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input15_A io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13671__A0 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ _14569_/X _18831_/Q _14759_/S vssd1 vssd1 vccd1 vccd1 _14752_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11963_ _16278_/A vssd1 vssd1 vccd1 vccd1 _11963_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_56_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13680__S _13686_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13702_ _13702_/A vssd1 vssd1 vccd1 vccd1 _18420_/D sky130_fd_sc_hd__clkbuf_1
X_17470_ _17390_/X _17459_/Y _17469_/X _17333_/X vssd1 vssd1 vccd1 vccd1 _17470_/X
+ sky130_fd_sc_hd__a211o_1
X_10914_ _10914_/A vssd1 vssd1 vccd1 vccd1 _11042_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14682_ _14682_/A vssd1 vssd1 vccd1 vccd1 _18800_/D sky130_fd_sc_hd__clkbuf_1
X_11894_ _11950_/A _11950_/C _11949_/A vssd1 vssd1 vccd1 vccd1 _11895_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__16276__B _16276_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10580__S0 _10579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16421_ _16423_/A _16423_/B _16402_/X vssd1 vssd1 vccd1 vccd1 _16421_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13633_ _13690_/S vssd1 vssd1 vccd1 vccd1 _13642_/S sky130_fd_sc_hd__buf_2
X_10845_ _10839_/A _10844_/X _09630_/A vssd1 vssd1 vccd1 vccd1 _10845_/Y sky130_fd_sc_hd__o21ai_1
X_19140_ _19635_/CLK _19140_/D vssd1 vssd1 vccd1 vccd1 _19140_/Q sky130_fd_sc_hd__dfxtp_1
X_16352_ _16388_/A _16352_/B _16352_/C vssd1 vssd1 vccd1 vccd1 _19433_/D sky130_fd_sc_hd__nor3_1
XANTENNA__12777__A2 _12773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ _13596_/A vssd1 vssd1 vccd1 vccd1 _13577_/S sky130_fd_sc_hd__buf_6
X_10776_ _19307_/Q _18719_/Q _18756_/Q _18330_/Q _10785_/S _09506_/A vssd1 vssd1 vccd1
+ vccd1 _10776_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10332__S0 _10286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15303_ _14601_/X _19065_/Q _15311_/S vssd1 vssd1 vccd1 vccd1 _15304_/A sky130_fd_sc_hd__mux2_1
X_12515_ _13005_/A vssd1 vssd1 vccd1 vccd1 _12515_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19071_ _19071_/CLK _19071_/D vssd1 vssd1 vccd1 vccd1 _19071_/Q sky130_fd_sc_hd__dfxtp_1
X_16283_ _16283_/A vssd1 vssd1 vccd1 vccd1 _19409_/D sky130_fd_sc_hd__clkbuf_1
X_13495_ _13274_/X _18346_/Q _13503_/S vssd1 vssd1 vccd1 vccd1 _13496_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16292__A _19414_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15400__S _15400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18022_ _18022_/A vssd1 vssd1 vccd1 vccd1 _19782_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16723__C _16750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12446_ _12446_/A vssd1 vssd1 vccd1 vccd1 _12446_/X sky130_fd_sc_hd__clkbuf_1
X_15234_ _15234_/A vssd1 vssd1 vccd1 vccd1 _19034_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12377_ _17125_/A _11516_/X _12302_/X vssd1 vssd1 vccd1 vccd1 _12377_/Y sky130_fd_sc_hd__o21ai_1
X_15165_ _19004_/Q _15089_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11328_ _10639_/X _11327_/X _09484_/A vssd1 vssd1 vccd1 vccd1 _11328_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_output83_A _12175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14116_ _13931_/X _18573_/Q _14118_/S vssd1 vssd1 vccd1 vccd1 _14117_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15096_ _18974_/Q _15095_/X _15099_/S vssd1 vssd1 vccd1 vccd1 _15097_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ _19086_/CLK _18924_/D vssd1 vssd1 vccd1 vccd1 _18924_/Q sky130_fd_sc_hd__dfxtp_1
X_11259_ _10943_/X _11252_/X _11254_/X _11258_/X _09464_/A vssd1 vssd1 vccd1 vccd1
+ _11259_/X sky130_fd_sc_hd__a311o_1
X_14047_ _14047_/A vssd1 vssd1 vccd1 vccd1 _18543_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16231__S _16235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09634__A _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18855_ _19365_/CLK _18855_/D vssd1 vssd1 vccd1 vccd1 _18855_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16979__A1 _15542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17806_ _17733_/A _17675_/X _17805_/Y _17386_/A vssd1 vssd1 vccd1 vccd1 _17806_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18786_ _19202_/CLK _18786_/D vssd1 vssd1 vccd1 vccd1 _18786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15998_ _15998_/A _19136_/Q vssd1 vssd1 vccd1 vccd1 _15998_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_83_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17737_ _17737_/A vssd1 vssd1 vccd1 vccd1 _17737_/X sky130_fd_sc_hd__buf_2
X_14949_ _14949_/A vssd1 vssd1 vccd1 vccd1 _18920_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_161_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19361_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13590__S _13593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17668_ _17419_/X _17658_/X _17666_/Y _17852_/A vssd1 vssd1 vccd1 vccd1 _17668_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_165_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19407_ _19838_/CLK _19407_/D vssd1 vssd1 vccd1 vccd1 _19407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16619_ _19832_/Q _16619_/B _19817_/Q _16619_/D vssd1 vssd1 vccd1 vccd1 _16625_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_126_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12217__A1 _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17599_ _17392_/X _17622_/A _17402_/X vssd1 vssd1 vccd1 vccd1 _17599_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19338_ _19356_/CLK _19338_/D vssd1 vssd1 vccd1 vccd1 _19338_/Q sky130_fd_sc_hd__dfxtp_2
Xclkbuf_leaf_176_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19369_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17156__A1 _17174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19269_ _19301_/CLK _19269_/D vssd1 vssd1 vccd1 vccd1 _19269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14715__A _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10626__S1 _10567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_114_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19645_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_132_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09924_ _19732_/Q vssd1 vssd1 vccd1 vccd1 _09924_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17616__C1 _17716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09855_ _18410_/Q _18671_/Q _18570_/Q _18905_/Q _09854_/X _09676_/A vssd1 vssd1 vccd1
+ vccd1 _09856_/B sky130_fd_sc_hd__mux4_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input7_A io_dbus_rdata[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09786_ _09786_/A vssd1 vssd1 vccd1 vccd1 _11387_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_129_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19796_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14596__S _14599_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13513__B _16000_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10622_/Y _10625_/Y _10627_/Y _10629_/Y _09572_/A vssd1 vssd1 vccd1 vccd1
+ _10630_/X sky130_fd_sc_hd__o221a_4
XFILLER_81_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10561_ _19280_/Q _19118_/Q _18527_/Q _18297_/Q _10542_/A _09443_/A vssd1 vssd1 vccd1
+ vccd1 _10562_/B sky130_fd_sc_hd__mux4_1
XFILLER_10_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15220__S _15228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12300_ _19417_/Q _12093_/X _12296_/X _12299_/Y vssd1 vssd1 vccd1 vccd1 _16298_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_139_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09719__A _10509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13280_ _19765_/Q vssd1 vssd1 vccd1 vccd1 _16142_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_155_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ _09761_/A _10478_/X _10490_/X _09834_/A _10491_/Y vssd1 vssd1 vccd1 vccd1
+ _12464_/B sky130_fd_sc_hd__o32a_4
XANTENNA__11968__B _11968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12231_ _19350_/Q _12274_/B _12230_/X vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_163_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16840__A _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12162_ _12162_/A vssd1 vssd1 vccd1 vccd1 _17802_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_146_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13675__S _13675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ _19300_/Q _18712_/Q _18749_/Q _18323_/Q _11112_/X _11075_/A vssd1 vssd1 vccd1
+ vccd1 _11113_/X sky130_fd_sc_hd__mux4_1
X_16970_ _16970_/A vssd1 vssd1 vccd1 vccd1 _16970_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12093_ _12093_/A vssd1 vssd1 vccd1 vccd1 _12093_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17607__C1 _17532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ _11044_/A _11044_/B _11044_/C vssd1 vssd1 vccd1 vccd1 _11044_/Y sky130_fd_sc_hd__nor3_1
X_15921_ _15921_/A vssd1 vssd1 vccd1 vccd1 _19295_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_104_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12695__A1 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10155__C1 _09754_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12695__B2 _12694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15890__S _15898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18640_ _19297_/CLK _18640_/D vssd1 vssd1 vccd1 vccd1 _18640_/Q sky130_fd_sc_hd__dfxtp_1
X_15852_ _13614_/X _19265_/Q _15852_/S vssd1 vssd1 vccd1 vccd1 _15853_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14803_ _14803_/A vssd1 vssd1 vccd1 vccd1 _18853_/D sky130_fd_sc_hd__clkbuf_1
X_18571_ _18990_/CLK _18571_/D vssd1 vssd1 vccd1 vccd1 _18571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15783_ _15839_/A vssd1 vssd1 vccd1 vccd1 _15852_/S sky130_fd_sc_hd__buf_6
XFILLER_149_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12995_ _12994_/A _13019_/C _12832_/A vssd1 vssd1 vccd1 vccd1 _12995_/X sky130_fd_sc_hd__o21a_1
XFILLER_73_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _17210_/X _17255_/X _17524_/S vssd1 vssd1 vccd1 vccd1 _17522_/X sky130_fd_sc_hd__mux2_1
X_14734_ _14734_/A vssd1 vssd1 vccd1 vccd1 _18823_/D sky130_fd_sc_hd__clkbuf_1
X_11946_ _11487_/S _12021_/A _12022_/A vssd1 vssd1 vccd1 vccd1 _11946_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_93_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19550_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13423__B _13423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17453_ _17535_/B vssd1 vssd1 vccd1 vccd1 _17625_/S sky130_fd_sc_hd__clkbuf_2
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14665_ _14550_/X _18793_/Q _14665_/S vssd1 vssd1 vccd1 vccd1 _14666_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _11877_/A vssd1 vssd1 vccd1 vccd1 _11877_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16404_ _19450_/Q _16406_/C _16403_/Y vssd1 vssd1 vccd1 vccd1 _19450_/D sky130_fd_sc_hd__o21a_1
X_13616_ _13616_/A vssd1 vssd1 vccd1 vccd1 _18384_/D sky130_fd_sc_hd__clkbuf_1
X_17384_ _17360_/X _17381_/X _17648_/S vssd1 vssd1 vccd1 vccd1 _17384_/X sky130_fd_sc_hd__mux2_1
X_10828_ _18585_/Q _18856_/Q _19080_/Q _18824_/Q _09598_/A _10802_/X vssd1 vssd1 vccd1
+ vccd1 _10828_/X sky130_fd_sc_hd__mux4_1
X_14596_ _14595_/X _18770_/Q _14599_/S vssd1 vssd1 vccd1 vccd1 _14597_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19123_ _19285_/CLK _19123_/D vssd1 vssd1 vccd1 vccd1 _19123_/Q sky130_fd_sc_hd__dfxtp_1
X_16335_ _16344_/A _16340_/C vssd1 vssd1 vccd1 vccd1 _16335_/Y sky130_fd_sc_hd__nor2_1
X_13547_ _15031_/A vssd1 vssd1 vccd1 vccd1 _13547_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10759_ _09597_/X _10756_/X _10758_/X _09602_/X vssd1 vssd1 vccd1 vccd1 _10759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18007__A _18029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19054_ _19054_/CLK _19054_/D vssd1 vssd1 vccd1 vccd1 _19054_/Q sky130_fd_sc_hd__dfxtp_1
X_16266_ _16266_/A _16266_/B vssd1 vssd1 vccd1 vccd1 _16267_/A sky130_fd_sc_hd__or2_1
X_13478_ _13478_/A vssd1 vssd1 vccd1 vccd1 _18338_/D sky130_fd_sc_hd__clkbuf_1
X_18005_ _19775_/Q _19396_/Q _18005_/S vssd1 vssd1 vccd1 vccd1 _18006_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15217_ _19027_/Q _15060_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__mux2_1
X_12429_ _12429_/A _12429_/B vssd1 vssd1 vccd1 vccd1 _12430_/C sky130_fd_sc_hd__xor2_2
XANTENNA__16750__A _19551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16197_ _16197_/A vssd1 vssd1 vccd1 vccd1 _19371_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_31_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19127_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12922__A2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15148_ _18996_/Q _15063_/X _15156_/S vssd1 vssd1 vccd1 vccd1 _15149_/A sky130_fd_sc_hd__mux2_1
XFILLER_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15079_ _15079_/A vssd1 vssd1 vccd1 vccd1 _15079_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18907_ _19390_/CLK _18907_/D vssd1 vssd1 vccd1 vccd1 _18907_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10146__C1 _09859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_46_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19089_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_42_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09640_ _10073_/A vssd1 vssd1 vccd1 vccd1 _09640_/X sky130_fd_sc_hd__buf_4
XFILLER_56_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18838_ _19320_/CLK _18838_/D vssd1 vssd1 vccd1 vccd1 _18838_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10303__A _10303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__S0 _10579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ _09571_/A vssd1 vssd1 vccd1 vccd1 _09572_/A sky130_fd_sc_hd__buf_4
X_18769_ _19320_/CLK _18769_/D vssd1 vssd1 vccd1 vccd1 _18769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15305__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16925__A input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11134__A _18782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12610__A1 _19331_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15975__S _15981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13495__S _13503_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09907_ _09952_/S vssd1 vssd1 vccd1 vccd1 _10112_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_76_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17491__A _17504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11309__A _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09838_ _18634_/Q _18969_/Q _09840_/S vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__mux2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15615__A1 _15612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09769_ _09769_/A vssd1 vssd1 vccd1 vccd1 _10270_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15215__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11800_ _19637_/Q _11801_/B vssd1 vssd1 vccd1 vccd1 _11802_/A sky130_fd_sc_hd__and2_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__A1 _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12780_ _12975_/A _12779_/Y _18744_/Q _09235_/B vssd1 vssd1 vccd1 vccd1 _12781_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_162_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _11683_/A _11683_/B _11730_/X vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__a21o_2
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14450_ _13845_/X _18711_/Q _14456_/S vssd1 vssd1 vccd1 vccd1 _14451_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11696_/B _11810_/S _19633_/Q vssd1 vssd1 vccd1 vccd1 _11662_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_42_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13401_ _15629_/A vssd1 vssd1 vccd1 vccd1 _15494_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_168_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10613_ _19310_/Q _18722_/Q _18759_/Q _18333_/Q _10546_/S _09419_/A vssd1 vssd1 vccd1
+ vccd1 _10614_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10883__A _18782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14381_ _14381_/A vssd1 vssd1 vccd1 vccd1 _18680_/D sky130_fd_sc_hd__clkbuf_1
X_11593_ _11579_/X _11580_/Y _11593_/S vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__mux2_4
XFILLER_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16120_ _16118_/X _19350_/Q _16140_/S vssd1 vssd1 vccd1 vccd1 _16121_/A sky130_fd_sc_hd__mux2_1
XFILLER_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10544_ _10612_/A _10544_/B vssd1 vssd1 vccd1 vccd1 _10544_/X sky130_fd_sc_hd__or2_1
X_13332_ _13332_/A vssd1 vssd1 vccd1 vccd1 _18311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15885__S _15887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10094__S _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16051_ _16055_/A _16055_/C vssd1 vssd1 vccd1 vccd1 _16051_/Y sky130_fd_sc_hd__xnor2_2
X_13263_ _19689_/Q _12529_/A _13009_/X _19656_/Q vssd1 vssd1 vccd1 vccd1 _13263_/X
+ sky130_fd_sc_hd__a22o_1
X_10475_ _10485_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10475_/Y sky130_fd_sc_hd__nor2_1
XFILLER_109_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15002_ _15002_/A vssd1 vssd1 vccd1 vccd1 _18944_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_68_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12214_ _17820_/B _12214_/B vssd1 vssd1 vccd1 vccd1 _12215_/B sky130_fd_sc_hd__and2_1
X_13194_ _13194_/A vssd1 vssd1 vccd1 vccd1 _18303_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19810_ _19866_/CLK _19810_/D vssd1 vssd1 vccd1 vccd1 _19810_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12025__D _17722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15186__A _15243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12145_ _12170_/A _17222_/A vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__or2_1
XFILLER_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16953_ _16953_/A _16970_/A vssd1 vssd1 vccd1 vccd1 _16953_/Y sky130_fd_sc_hd__nand2_1
X_12076_ _19647_/Q _12105_/C vssd1 vssd1 vccd1 vccd1 _12076_/Y sky130_fd_sc_hd__nor2_1
XFILLER_111_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19741_ _19779_/CLK _19741_/D vssd1 vssd1 vccd1 vccd1 _19741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13418__B _13418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13865__A0 _13864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15904_ _15904_/A vssd1 vssd1 vccd1 vccd1 _19287_/D sky130_fd_sc_hd__clkbuf_1
X_11027_ _19271_/Q _19109_/Q _18518_/Q _18288_/Q _11149_/A _09512_/A vssd1 vssd1 vccd1
+ vccd1 _11027_/X sky130_fd_sc_hd__mux4_1
X_19672_ _19694_/CLK _19672_/D vssd1 vssd1 vccd1 vccd1 _19672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16884_ _19606_/Q _16881_/B _16883_/Y vssd1 vssd1 vccd1 vccd1 _19606_/D sky130_fd_sc_hd__o21a_1
XFILLER_65_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10774__S0 _10633_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18623_ _19086_/CLK _18623_/D vssd1 vssd1 vccd1 vccd1 _18623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15835_ _13589_/X _19257_/Q _15837_/S vssd1 vssd1 vccd1 vccd1 _15836_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11891__A2 _12455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13434__A _14197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18554_ _18824_/CLK _18554_/D vssd1 vssd1 vccd1 vccd1 _18554_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15766_ _15766_/A vssd1 vssd1 vccd1 vccd1 _19226_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13093__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12978_ input31/X _12974_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _12978_/X sky130_fd_sc_hd__a21o_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17505_/A vssd1 vssd1 vccd1 vccd1 _17505_/Y sky130_fd_sc_hd__inv_2
X_14717_ _14785_/S vssd1 vssd1 vccd1 vccd1 _14726_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_61_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09350__C _18122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__A3 _10444_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _11929_/A _11929_/B vssd1 vssd1 vccd1 vccd1 _11931_/A sky130_fd_sc_hd__nor2_1
X_18485_ _19012_/CLK _18485_/D vssd1 vssd1 vccd1 vccd1 _18485_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15697_ _15697_/A vssd1 vssd1 vccd1 vccd1 _19195_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17436_ _17511_/S _17242_/X _17435_/X vssd1 vssd1 vccd1 vccd1 _17436_/Y sky130_fd_sc_hd__o21ai_1
X_14648_ _14525_/X _18785_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14649_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17367_ _17276_/X _17264_/X _17367_/S vssd1 vssd1 vccd1 vccd1 _17368_/A sky130_fd_sc_hd__mux2_1
X_14579_ _14579_/A vssd1 vssd1 vccd1 vccd1 _14579_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10829__S1 _10817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19106_ _19268_/CLK _19106_/D vssd1 vssd1 vccd1 vccd1 _19106_/Q sky130_fd_sc_hd__dfxtp_1
X_16318_ _19485_/Q _19484_/Q _19486_/Q _16496_/A vssd1 vssd1 vccd1 vccd1 _16324_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__09359__A _17795_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17298_ _17288_/X _17296_/X _17615_/A vssd1 vssd1 vccd1 vccd1 _17298_/X sky130_fd_sc_hd__mux2_1
XFILLER_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19037_ _19389_/CLK _19037_/D vssd1 vssd1 vccd1 vccd1 _19037_/Q sky130_fd_sc_hd__dfxtp_1
X_16249_ _16255_/A _16249_/B vssd1 vssd1 vccd1 vccd1 _16250_/A sky130_fd_sc_hd__or2_1
XFILLER_161_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 _11877_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[9] sky130_fd_sc_hd__buf_2
XFILLER_127_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput113 _12460_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[13] sky130_fd_sc_hd__buf_2
XFILLER_126_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput124 _12472_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[23] sky130_fd_sc_hd__buf_2
XFILLER_142_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput135 _12447_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[4] sky130_fd_sc_hd__buf_2
Xoutput146 _16272_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[13] sky130_fd_sc_hd__buf_2
XFILLER_99_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput157 _16295_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[23] sky130_fd_sc_hd__buf_2
Xoutput168 _16251_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[4] sky130_fd_sc_hd__buf_2
XANTENNA__12513__A _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11006__S1 _11005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17598__A1 _17731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09822__A _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ _10969_/A vssd1 vssd1 vccd1 vccd1 _09624_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16270__A1 _11969_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ _09658_/A vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__buf_4
XFILLER_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11095__B1 _11070_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14874__S _14882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09485_ _09485_/A vssd1 vssd1 vccd1 vccd1 _10296_/A sky130_fd_sc_hd__buf_2
XFILLER_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_164_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ _10260_/A vssd1 vssd1 vccd1 vccd1 _10260_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_118_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12898__A1 _19557_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16089__A1 _19345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17286__A0 _12309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ _10200_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10191_/X sky130_fd_sc_hd__or2_1
XFILLER_121_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14114__S _14118_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15734__A _15780_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11039__A _11219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13950_ _14049_/S vssd1 vssd1 vccd1 vccd1 _13963_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18110__A _18136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11322__A1 _09651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10756__S0 _10660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09610__S1 _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ _19593_/Q _12560_/X _12562_/X _19461_/Q _12900_/X vssd1 vssd1 vccd1 vccd1
+ _15485_/B sky130_fd_sc_hd__a221o_2
XFILLER_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13881_ _13880_/X _18493_/Q _13887_/S vssd1 vssd1 vccd1 vccd1 _13882_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10676__A3 _10675_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__A _10878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ _15612_/X _18279_/Q _09234_/X _13398_/X _15619_/X vssd1 vssd1 vccd1 vccd1
+ _15620_/X sky130_fd_sc_hd__a32o_2
XFILLER_28_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13254__A _13254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12832_ _12832_/A vssd1 vssd1 vccd1 vccd1 _13113_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09279__B1 _12606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10597__B _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15601_/A vssd1 vssd1 vccd1 vccd1 _15569_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _18271_/Q _12759_/X _10303_/A _12762_/X vssd1 vssd1 vccd1 vccd1 _18271_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11625__A2 _11612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14502_/A vssd1 vssd1 vccd1 vccd1 _14511_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18270_ _19162_/CLK _18270_/D vssd1 vssd1 vccd1 vccd1 _18270_/Q sky130_fd_sc_hd__dfxtp_1
X_11714_ _11723_/S _12444_/B _11632_/Y vssd1 vssd1 vccd1 vccd1 _17256_/A sky130_fd_sc_hd__o21a_1
XFILLER_42_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15482_ _19711_/Q _15481_/X _15482_/S vssd1 vssd1 vccd1 vccd1 _15482_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _18142_/B vssd1 vssd1 vccd1 vccd1 _12694_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17221_ _17221_/A vssd1 vssd1 vccd1 vccd1 _17696_/B sky130_fd_sc_hd__clkbuf_4
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _13925_/X _18704_/Q _14439_/S vssd1 vssd1 vccd1 vccd1 _14434_/A sky130_fd_sc_hd__mux2_1
X_11645_ _12100_/A vssd1 vssd1 vccd1 vccd1 _12372_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17152_ _17152_/A vssd1 vssd1 vccd1 vccd1 _19702_/D sky130_fd_sc_hd__clkbuf_1
Xinput15 io_dbus_rdata[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_4
X_14364_ _14364_/A vssd1 vssd1 vccd1 vccd1 _18674_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput26 io_dbus_rdata[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_4
XFILLER_11_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11576_ _09171_/B _09124_/A _09124_/B vssd1 vssd1 vccd1 vccd1 _11577_/C sky130_fd_sc_hd__o21ai_1
XFILLER_156_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput37 io_ibus_inst[12] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 io_ibus_inst[22] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16103_ _16107_/A _16107_/C vssd1 vssd1 vccd1 vccd1 _16103_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__15524__A0 _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput59 io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_1
X_13315_ _19766_/Q _19767_/Q _13315_/C vssd1 vssd1 vccd1 vccd1 _13336_/B sky130_fd_sc_hd__and3_1
X_17083_ _19688_/Q _12715_/X _17083_/S vssd1 vssd1 vccd1 vccd1 _17084_/A sky130_fd_sc_hd__mux2_1
X_10527_ _18592_/Q _18863_/Q _19087_/Q _18831_/Q _10481_/S _10262_/A vssd1 vssd1 vccd1
+ vccd1 _10527_/X sky130_fd_sc_hd__mux4_1
XFILLER_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14295_ _14635_/A _18224_/B vssd1 vssd1 vccd1 vccd1 _14296_/A sky130_fd_sc_hd__and2_1
XFILLER_109_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12338__B1 _19419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16034_ _16034_/A vssd1 vssd1 vccd1 vccd1 _19335_/D sky130_fd_sc_hd__clkbuf_1
X_10458_ _10250_/A _10455_/X _10457_/X _10243_/A vssd1 vssd1 vccd1 vccd1 _10458_/X
+ sky130_fd_sc_hd__o211a_1
X_13246_ _13245_/A _13256_/C _12832_/A vssd1 vssd1 vccd1 vccd1 _13246_/X sky130_fd_sc_hd__o21a_1
XFILLER_170_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17816__A2 _17658_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10389_ _19188_/Q _18802_/Q _19252_/Q _18371_/Q _10274_/X _10263_/X vssd1 vssd1 vccd1
+ vccd1 _10390_/B sky130_fd_sc_hd__mux4_1
XANTENNA__14024__S _14027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ _13234_/A _13177_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13177_/X sky130_fd_sc_hd__or3_1
XFILLER_111_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11561__A1 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12128_ _12369_/A _12123_/Y _12127_/X _11686_/X vssd1 vssd1 vccd1 vccd1 _12128_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_2_0_clock_A clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17985_ _17985_/A vssd1 vssd1 vccd1 vccd1 _19765_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16936_ _19630_/Q _16931_/X _16935_/X _16933_/X vssd1 vssd1 vccd1 vccd1 _19630_/D
+ sky130_fd_sc_hd__o211a_1
X_19724_ _19724_/CLK _19724_/D vssd1 vssd1 vccd1 vccd1 _19724_/Q sky130_fd_sc_hd__dfxtp_4
X_12059_ _12059_/A _12059_/B vssd1 vssd1 vccd1 vccd1 _12060_/A sky130_fd_sc_hd__xnor2_1
XFILLER_42_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09601__S1 _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19655_ _19660_/CLK _19655_/D vssd1 vssd1 vccd1 vccd1 _19655_/Q sky130_fd_sc_hd__dfxtp_1
X_16867_ _19600_/Q _16864_/B _16866_/Y vssd1 vssd1 vccd1 vccd1 _19600_/D sky130_fd_sc_hd__o21a_1
XFILLER_92_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15818_ _13563_/X _19249_/Q _15826_/S vssd1 vssd1 vccd1 vccd1 _15819_/A sky130_fd_sc_hd__mux2_1
XFILLER_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18606_ _19389_/CLK _18606_/D vssd1 vssd1 vccd1 vccd1 _18606_/Q sky130_fd_sc_hd__dfxtp_1
X_19586_ _19586_/CLK _19586_/D vssd1 vssd1 vccd1 vccd1 _19586_/Q sky130_fd_sc_hd__dfxtp_1
X_16798_ _19573_/Q _16800_/B _19571_/Q _16798_/D vssd1 vssd1 vccd1 vccd1 _16807_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_92_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18537_ _19290_/CLK _18537_/D vssd1 vssd1 vccd1 vccd1 _18537_/Q sky130_fd_sc_hd__dfxtp_1
X_15749_ _15749_/A vssd1 vssd1 vccd1 vccd1 _19218_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14694__S _14698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16004__A1 _19330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09270_ _09270_/A _09270_/B vssd1 vssd1 vccd1 vccd1 _09271_/D sky130_fd_sc_hd__or2_1
X_18468_ _19124_/CLK _18468_/D vssd1 vssd1 vccd1 vccd1 _18468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17419_ _17419_/A vssd1 vssd1 vccd1 vccd1 _17419_/X sky130_fd_sc_hd__clkbuf_2
X_18399_ _18894_/CLK _18399_/D vssd1 vssd1 vccd1 vccd1 _18399_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_159_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11227__S1 _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14869__S _14871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__C1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10738__S0 _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09606_ _09717_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _09606_/X sky130_fd_sc_hd__or2_1
XFILLER_83_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__B _13391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13057__B2 _19341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09537_ _10631_/S vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11163__S0 _10904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09468_ _09468_/A vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__buf_2
XFILLER_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_164_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ _10603_/S vssd1 vssd1 vccd1 vccd1 _10602_/S sky130_fd_sc_hd__buf_2
XFILLER_8_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _11433_/A _11431_/C _11431_/A vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__a21o_1
XFILLER_138_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09984__A1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11361_ _11361_/A _11361_/B vssd1 vssd1 vccd1 vccd1 _11415_/A sky130_fd_sc_hd__nand2_1
XFILLER_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12852__S _12887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14633__A _14633_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13100_ _19439_/Q _13005_/A _13099_/X vssd1 vssd1 vccd1 vccd1 _13100_/X sky130_fd_sc_hd__o21a_1
XFILLER_152_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ _10312_/A vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__buf_2
XFILLER_4_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09727__A _09727_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14080_ _14080_/A vssd1 vssd1 vccd1 vccd1 _18556_/D sky130_fd_sc_hd__clkbuf_1
X_11292_ _11461_/A _11292_/B vssd1 vssd1 vccd1 vccd1 _11463_/C sky130_fd_sc_hd__nand2_1
XFILLER_106_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10243_ _10243_/A vssd1 vssd1 vccd1 vccd1 _10243_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_106_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13031_ _19750_/Q _13031_/B vssd1 vssd1 vccd1 vccd1 _13064_/C sky130_fd_sc_hd__and2_1
XFILLER_106_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input45_A io_ibus_inst[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10174_ _10174_/A _10174_/B vssd1 vssd1 vccd1 vccd1 _10174_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14779__S _14781_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15464__A _15603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17770_ _17673_/A _17733_/B _17767_/Y _17769_/X vssd1 vssd1 vccd1 vccd1 _17771_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_120_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14982_ _18937_/Q vssd1 vssd1 vccd1 vccd1 _14983_/A sky130_fd_sc_hd__clkbuf_1
X_16721_ _16724_/C _16724_/D _19550_/Q vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_89_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13933_ _13933_/A vssd1 vssd1 vccd1 vccd1 _18509_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_93_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12600__B _12600_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19440_ _19583_/CLK _19440_/D vssd1 vssd1 vccd1 vccd1 _19440_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17431__B1 _09315_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16652_ _19528_/Q _16663_/D vssd1 vssd1 vccd1 vccd1 _16655_/B sky130_fd_sc_hd__and2_1
XFILLER_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13864_ _14544_/A vssd1 vssd1 vccd1 vccd1 _13864_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10401__A _10401_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15603_ _15603_/A vssd1 vssd1 vccd1 vccd1 _15627_/S sky130_fd_sc_hd__clkbuf_2
X_12815_ _19589_/Q vssd1 vssd1 vccd1 vccd1 _16836_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19371_ _19373_/CLK _19371_/D vssd1 vssd1 vccd1 vccd1 _19371_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16583_ _19508_/Q _16584_/C _19509_/Q vssd1 vssd1 vccd1 vccd1 _16585_/B sky130_fd_sc_hd__a21oi_1
X_13795_ _13795_/A vssd1 vssd1 vccd1 vccd1 _18461_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11154__S0 _10904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18322_ _19235_/CLK _18322_/D vssd1 vssd1 vccd1 vccd1 _18322_/Q sky130_fd_sc_hd__dfxtp_1
X_15534_ hold11/A _15534_/B vssd1 vssd1 vccd1 vccd1 _15534_/X sky130_fd_sc_hd__or2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ hold18/A _12744_/X _10798_/A _12740_/X vssd1 vssd1 vccd1 vccd1 _18260_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17734__B2 _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18253_ _19720_/CLK _18253_/D vssd1 vssd1 vccd1 vccd1 _18253_/Q sky130_fd_sc_hd__dfxtp_2
X_15465_ _15636_/S vssd1 vssd1 vccd1 vccd1 _15483_/S sky130_fd_sc_hd__buf_2
XANTENNA__16942__C1 _16833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12677_ _12677_/A vssd1 vssd1 vccd1 vccd1 _12677_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17204_ _17680_/B _17802_/B _17263_/A vssd1 vssd1 vccd1 vccd1 _17204_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11232__A _11232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14416_ _14416_/A vssd1 vssd1 vccd1 vccd1 _18696_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18184_ _18184_/A vssd1 vssd1 vccd1 vccd1 _19844_/D sky130_fd_sc_hd__clkbuf_1
X_11628_ _17225_/A _17207_/A _11840_/A vssd1 vssd1 vccd1 vccd1 _11634_/A sky130_fd_sc_hd__o21ai_1
X_15396_ _19106_/Q _15006_/X _15400_/S vssd1 vssd1 vccd1 vccd1 _15397_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17135_ _17142_/A _17135_/B vssd1 vssd1 vccd1 vccd1 _17136_/A sky130_fd_sc_hd__and2_1
X_14347_ _14347_/A vssd1 vssd1 vccd1 vccd1 _18666_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15639__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11559_ _11559_/A vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_171_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_155_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17066_ _19680_/Q _12550_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17067_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14278_ _14623_/A vssd1 vssd1 vccd1 vccd1 _14278_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16017_ _16021_/A _16021_/C vssd1 vssd1 vccd1 vccd1 _16017_/Y sky130_fd_sc_hd__xnor2_2
X_13229_ _13228_/X _18305_/Q _13252_/S vssd1 vssd1 vccd1 vccd1 _13230_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17854__A _17856_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12731__B1 _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_151_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12998__A _15028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13593__S _13593_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17968_ _19758_/Q _19790_/Q _17968_/S vssd1 vssd1 vccd1 vccd1 _17969_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09372__A _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19707_ _19724_/CLK _19707_/D vssd1 vssd1 vccd1 vccd1 _19707_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09586__S0 _10030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16919_ _16919_/A vssd1 vssd1 vccd1 vccd1 _16932_/A sky130_fd_sc_hd__buf_2
X_17899_ _17899_/A _17899_/B vssd1 vssd1 vccd1 vccd1 _17899_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10196__S1 _09676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19638_ _19669_/CLK _19638_/D vssd1 vssd1 vccd1 vccd1 _19638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19569_ _19668_/CLK _19569_/D vssd1 vssd1 vccd1 vccd1 _19569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15313__S _15315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13622__A _13690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ _17994_/S vssd1 vssd1 vccd1 vccd1 _09322_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__09889__S1 _09888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10273__A1 _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09253_ _16623_/A _16623_/B _09253_/C _09253_/D vssd1 vssd1 vccd1 vccd1 _09270_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_167_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09184_ _18077_/A _18075_/A _09236_/C _09236_/D vssd1 vssd1 vccd1 vccd1 _11560_/B
+ sky130_fd_sc_hd__nand4b_4
XFILLER_105_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10025__A1 _09557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09966__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13768__S _13776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09547__A _09547_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13069__A _15041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17764__A _17768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12722__A0 hold21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__S _09981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14599__S _14599_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13278__A1 input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_90_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_112_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10930_ _10919_/Y _10924_/Y _10926_/Y _10928_/Y _11044_/A vssd1 vssd1 vccd1 vccd1
+ _10930_/X sky130_fd_sc_hd__o221a_1
XFILLER_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17964__A1 _19788_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_95_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ _11263_/S vssd1 vssd1 vccd1 vccd1 _11071_/S sky130_fd_sc_hd__buf_4
XFILLER_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12600_ _12602_/B _12600_/B vssd1 vssd1 vccd1 vccd1 _12600_/Y sky130_fd_sc_hd__nor2_1
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13532__A _13615_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13596_/A vssd1 vssd1 vccd1 vccd1 _13593_/S sky130_fd_sc_hd__buf_6
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10792_ _18586_/Q _18857_/Q _19081_/Q _18825_/Q _10579_/X _10060_/A vssd1 vssd1 vccd1
+ vccd1 _10792_/X sky130_fd_sc_hd__mux4_1
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12677_/A vssd1 vssd1 vccd1 vccd1 _12958_/A sky130_fd_sc_hd__clkbuf_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10367__S _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15250_ _14525_/X _19041_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15251_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12462_ _12462_/A _12462_/B vssd1 vssd1 vccd1 vccd1 _12462_/Y sky130_fd_sc_hd__nor2_1
XFILLER_173_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14201_ _18609_/Q _13943_/X _14209_/S vssd1 vssd1 vccd1 vccd1 _14202_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13678__S _13686_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09957__A1 _09905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11413_ _11413_/A _12480_/B vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__or2_1
XFILLER_172_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15181_ _15181_/A vssd1 vssd1 vccd1 vccd1 _19010_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12393_ _19357_/Q _12069_/X _11686_/X _12392_/X _12071_/X vssd1 vssd1 vccd1 vccd1
+ _12393_/X sky130_fd_sc_hd__o221a_1
XFILLER_153_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14132_ _18579_/Q _13956_/X _14136_/S vssd1 vssd1 vccd1 vccd1 _14133_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09457__A _10046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _11344_/A vssd1 vssd1 vccd1 vccd1 _11344_/Y sky130_fd_sc_hd__inv_2
XFILLER_126_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14063_ _13854_/X _18549_/Q _14063_/S vssd1 vssd1 vccd1 vccd1 _14064_/A sky130_fd_sc_hd__mux2_1
X_18940_ _19388_/CLK _18940_/D vssd1 vssd1 vccd1 vccd1 _18940_/Q sky130_fd_sc_hd__dfxtp_1
X_11275_ _19298_/Q _18710_/Q _18747_/Q _18321_/Q _11071_/S _11220_/A vssd1 vssd1 vccd1
+ vccd1 _11275_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13014_ _19434_/Q _13005_/X _13013_/X vssd1 vssd1 vccd1 vccd1 _13014_/X sky130_fd_sc_hd__o21a_1
X_10226_ _09762_/A _10212_/X _10224_/X _09835_/A _10225_/Y vssd1 vssd1 vccd1 vccd1
+ _12470_/B sky130_fd_sc_hd__o32a_4
XANTENNA_output151_A _12136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18871_ _19291_/CLK _18871_/D vssd1 vssd1 vccd1 vccd1 _18871_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10157_ _18471_/Q _19062_/Q _19224_/Q _18439_/Q _10114_/S _09888_/X vssd1 vssd1 vccd1
+ vccd1 _10158_/B sky130_fd_sc_hd__mux4_1
X_17822_ _17710_/S _17823_/B _17821_/X _17466_/X vssd1 vssd1 vccd1 vccd1 _17822_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14302__S _14310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14965_ _14965_/A vssd1 vssd1 vccd1 vccd1 _18928_/D sky130_fd_sc_hd__clkbuf_1
X_17753_ _17753_/A _17756_/B vssd1 vssd1 vccd1 vccd1 _17753_/Y sky130_fd_sc_hd__nand2_1
X_10088_ _10088_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__and2_1
XFILLER_63_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16704_ _19544_/Q _19543_/Q _19542_/Q _16704_/D vssd1 vssd1 vccd1 vccd1 _16712_/D
+ sky130_fd_sc_hd__and4_1
X_13916_ _13915_/X _18504_/Q _13919_/S vssd1 vssd1 vccd1 vccd1 _13917_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17684_ _17684_/A vssd1 vssd1 vccd1 vccd1 _17684_/Y sky130_fd_sc_hd__clkinv_2
X_14896_ _18895_/Q _13997_/X _14904_/S vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17955__A1 _19784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16635_ _16666_/A _16635_/B vssd1 vssd1 vccd1 vccd1 _16635_/Y sky130_fd_sc_hd__nor2_1
X_19423_ _19423_/CLK _19423_/D vssd1 vssd1 vccd1 vccd1 _19423_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09920__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _13847_/A vssd1 vssd1 vccd1 vccd1 _18482_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16229__S _16235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14538__A _14621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16566_ hold1/X _16567_/C _19503_/Q vssd1 vssd1 vccd1 vccd1 _16568_/B sky130_fd_sc_hd__a21oi_1
X_19354_ _19357_/CLK _19354_/D vssd1 vssd1 vccd1 vccd1 _19354_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13778_ _13835_/S vssd1 vssd1 vccd1 vccd1 _13787_/S sky130_fd_sc_hd__buf_2
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18305_ _18902_/CLK _18305_/D vssd1 vssd1 vccd1 vccd1 _18305_/Q sky130_fd_sc_hd__dfxtp_1
X_15517_ _15516_/X _19147_/Q _15517_/S vssd1 vssd1 vccd1 vccd1 _15518_/A sky130_fd_sc_hd__mux2_1
X_19285_ _19285_/CLK _19285_/D vssd1 vssd1 vccd1 vccd1 _19285_/Q sky130_fd_sc_hd__dfxtp_1
X_12729_ _12769_/A vssd1 vssd1 vccd1 vccd1 _12747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_149_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16497_ _16524_/A _16501_/C vssd1 vssd1 vccd1 vccd1 _16497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18236_ _18248_/A _18236_/B vssd1 vssd1 vccd1 vccd1 _18237_/A sky130_fd_sc_hd__and2_1
X_15448_ _15448_/A vssd1 vssd1 vccd1 vccd1 _19129_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16930__A2 _12674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__A1 _10289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09948__A1 _09844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18167_ _18167_/A vssd1 vssd1 vccd1 vccd1 _19840_/D sky130_fd_sc_hd__clkbuf_1
X_15379_ _19099_/Q _15086_/X _15383_/S vssd1 vssd1 vccd1 vccd1 _15380_/A sky130_fd_sc_hd__mux2_1
X_17118_ _18100_/A _09210_/X _17115_/X _17175_/B vssd1 vssd1 vccd1 vccd1 _17118_/X
+ sky130_fd_sc_hd__a31o_1
X_18098_ _19846_/Q _12694_/X _18096_/Y _18097_/X vssd1 vssd1 vccd1 vccd1 _19814_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_172_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_172_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17049_ _17049_/A vssd1 vssd1 vccd1 vccd1 _19672_/D sky130_fd_sc_hd__clkbuf_1
X_09940_ _19322_/Q _18734_/Q _18771_/Q _18345_/Q _10137_/S _10090_/A vssd1 vssd1 vccd1
+ vccd1 _09941_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09871_ _09871_/A vssd1 vssd1 vccd1 vccd1 _09871_/X sky130_fd_sc_hd__clkbuf_4
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_112_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12180__A1 _19348_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13617__A _14297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12521__A _12521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09830__A _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ _09305_/A _09305_/B vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__nor2_1
XFILLER_142_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14882__S _14882_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09236_ _18077_/A _18075_/A _09236_/C _09236_/D vssd1 vssd1 vccd1 vccd1 _11569_/B
+ sky130_fd_sc_hd__and4_2
XANTENNA_clkbuf_leaf_37_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09939__A1 _09844_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13196__B1 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09167_ _09167_/A _09167_/B _09167_/C vssd1 vssd1 vccd1 vccd1 _17165_/B sky130_fd_sc_hd__or3_1
XFILLER_119_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09098_ _19837_/Q vssd1 vssd1 vccd1 vccd1 _18075_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_108_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11060_ _11208_/A vssd1 vssd1 vccd1 vccd1 _11188_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10011_ _10289_/A _10010_/X _09485_/A vssd1 vssd1 vccd1 vccd1 _10011_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14448__A0 _13837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14122__S _14122_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16838__A _16838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14750_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14759_/S sky130_fd_sc_hd__buf_6
XFILLER_85_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11962_ _11962_/A vssd1 vssd1 vccd1 vccd1 _16278_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_57_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ _12865_/X _18420_/Q _13703_/S vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15948__A0 _13544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _18584_/Q _18855_/Q _19079_/Q _18823_/Q _10852_/S _10837_/A vssd1 vssd1 vccd1
+ vccd1 _10913_/X sky130_fd_sc_hd__mux4_1
X_14681_ _14573_/X _18800_/Q _14687_/S vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11893_ _11893_/A _17642_/A vssd1 vssd1 vccd1 vccd1 _11950_/C sky130_fd_sc_hd__or2_1
XFILLER_72_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16420_ _16423_/A _16833_/A vssd1 vssd1 vccd1 vccd1 _19456_/D sky130_fd_sc_hd__nor2_1
XANTENNA__10580__S1 _10060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13632_ _13632_/A vssd1 vssd1 vccd1 vccd1 _18389_/D sky130_fd_sc_hd__clkbuf_1
X_10844_ _19306_/Q _18718_/Q _18755_/Q _18329_/Q _10854_/S _10837_/X vssd1 vssd1 vccd1
+ vccd1 _10844_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16351_ _19433_/Q _16351_/B _16351_/C vssd1 vssd1 vccd1 vccd1 _16352_/C sky130_fd_sc_hd__and3_1
X_13563_ _15047_/A vssd1 vssd1 vccd1 vccd1 _13563_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10775_ _10779_/A _10775_/B vssd1 vssd1 vccd1 vccd1 _10775_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10332__S1 _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ _15302_/A vssd1 vssd1 vccd1 vccd1 _15311_/S sky130_fd_sc_hd__buf_4
X_12514_ _12962_/A vssd1 vssd1 vccd1 vccd1 _13005_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__15176__A1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19070_ _19264_/CLK _19070_/D vssd1 vssd1 vccd1 vccd1 _19070_/Q sky130_fd_sc_hd__dfxtp_1
X_16282_ _16282_/A _16282_/B vssd1 vssd1 vccd1 vccd1 _16283_/A sky130_fd_sc_hd__and2_1
X_13494_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13503_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_173_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18021_ _19782_/Q _11969_/B _18027_/S vssd1 vssd1 vccd1 vccd1 _18022_/A sky130_fd_sc_hd__mux2_1
X_15233_ _19034_/Q _15083_/X _15239_/S vssd1 vssd1 vccd1 vccd1 _15234_/A sky130_fd_sc_hd__mux2_1
XFILLER_138_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12445_ _12450_/A _12445_/B vssd1 vssd1 vccd1 vccd1 _12446_/A sky130_fd_sc_hd__and2b_1
XFILLER_139_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10825__S _10872_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11510__A _17166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ _15164_/A vssd1 vssd1 vccd1 vccd1 _19003_/D sky130_fd_sc_hd__clkbuf_1
X_12376_ _12366_/Y _12134_/X _12375_/X vssd1 vssd1 vccd1 vccd1 _12376_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_125_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17873__A0 _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ _14115_/A vssd1 vssd1 vccd1 vccd1 _18572_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ _18590_/Q _18861_/Q _19085_/Q _18829_/Q _10579_/X _10705_/A vssd1 vssd1 vccd1
+ vccd1 _11327_/X sky130_fd_sc_hd__mux4_1
XFILLER_114_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15095_ _15095_/A vssd1 vssd1 vccd1 vccd1 _15095_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_140_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_107_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18923_ _19085_/CLK _18923_/D vssd1 vssd1 vccd1 vccd1 _18923_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output76_A _12009_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ _18543_/Q _14045_/X _14049_/S vssd1 vssd1 vccd1 vccd1 _14047_/A sky130_fd_sc_hd__mux2_1
X_11258_ _11252_/A _11255_/X _11257_/X _11134_/X vssd1 vssd1 vccd1 vccd1 _11258_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10209_/Y sky130_fd_sc_hd__nor2_1
X_18854_ _19367_/CLK _18854_/D vssd1 vssd1 vccd1 vccd1 _18854_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11189_ _19269_/Q _19107_/Q _18516_/Q _18286_/Q _10873_/S _11177_/X vssd1 vssd1 vccd1
+ vccd1 _11189_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17805_ _17597_/X _17687_/B _17804_/X vssd1 vssd1 vccd1 vccd1 _17805_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_95_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18785_ _19235_/CLK _18785_/D vssd1 vssd1 vccd1 vccd1 _18785_/Q sky130_fd_sc_hd__dfxtp_1
X_15997_ _15997_/A vssd1 vssd1 vccd1 vccd1 _19329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13871__S _13871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14948_ _18920_/Q vssd1 vssd1 vccd1 vccd1 _14949_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17736_ _17736_/A vssd1 vssd1 vccd1 vccd1 _19721_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11673__A0 _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ _17871_/A vssd1 vssd1 vccd1 vccd1 _17852_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_14879_ _14879_/A vssd1 vssd1 vccd1 vccd1 _18887_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19406_ _19807_/CLK _19406_/D vssd1 vssd1 vccd1 vccd1 _19406_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_62_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16618_ _09301_/A _09301_/B _11551_/B _11702_/C vssd1 vssd1 vccd1 vccd1 _16626_/C
+ sky130_fd_sc_hd__o31ai_1
X_17598_ _17731_/S _17257_/X _17457_/X vssd1 vssd1 vccd1 vccd1 _17622_/A sky130_fd_sc_hd__o21ai_2
XFILLER_51_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16549_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16585_/A sky130_fd_sc_hd__clkbuf_2
X_19337_ _19356_/CLK _19337_/D vssd1 vssd1 vccd1 vccd1 _19337_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_148_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19268_ _19268_/CLK _19268_/D vssd1 vssd1 vccd1 vccd1 _19268_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14715__B _14860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18219_ _18219_/A vssd1 vssd1 vccd1 vccd1 _19856_/D sky130_fd_sc_hd__clkbuf_1
X_19199_ _19249_/CLK _19199_/D vssd1 vssd1 vccd1 vccd1 _19199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_129_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14207__S _14209_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11420__A _11420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_144_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_160_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09923_ _09914_/Y _09917_/Y _09920_/Y _09922_/Y _09831_/X vssd1 vssd1 vccd1 vccd1
+ _09923_/X sky130_fd_sc_hd__o221a_1
XANTENNA__15546__B _15546_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_160_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09854_ _10367_/S vssd1 vssd1 vccd1 vccd1 _09854_/X sky130_fd_sc_hd__buf_4
XFILLER_105_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10164__B1 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17092__A1 _15620_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09785_ _09785_/A vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__buf_2
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__A1 _12230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09609__B1 _09995_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10560_ _18463_/Q _19054_/Q _19216_/Q _18431_/Q _09415_/A _09443_/X vssd1 vssd1 vccd1
+ vccd1 _10560_/X sky130_fd_sc_hd__mux4_2
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14625__B _18205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _19814_/Q vssd1 vssd1 vccd1 vccd1 _13619_/A sky130_fd_sc_hd__inv_4
XFILLER_154_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _19723_/Q vssd1 vssd1 vccd1 vccd1 _10491_/Y sky130_fd_sc_hd__inv_2
XFILLER_154_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _12230_/A vssd1 vssd1 vccd1 vccd1 _12230_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_136_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12145__B _17222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12392__A1 _12389_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12161_ _12208_/A _12468_/B _12160_/Y vssd1 vssd1 vccd1 vccd1 _12162_/A sky130_fd_sc_hd__o21ai_1
XFILLER_122_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14641__A _14641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11112_ _11219_/S vssd1 vssd1 vccd1 vccd1 _11112_/X sky130_fd_sc_hd__buf_2
XFILLER_150_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12092_ _12092_/A vssd1 vssd1 vccd1 vccd1 _12092_/Y sky130_fd_sc_hd__inv_2
XFILLER_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13341__B1 _13340_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11043_ _11026_/A _11038_/X _11041_/X _11042_/X vssd1 vssd1 vccd1 vccd1 _11044_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15920_ _19295_/Q _14614_/A _15920_/S vssd1 vssd1 vccd1 vccd1 _15921_/A sky130_fd_sc_hd__mux2_1
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17083__A1 _12715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ _15851_/A vssd1 vssd1 vccd1 vccd1 _19264_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_162_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14802_ _18853_/Q _13965_/X _14810_/S vssd1 vssd1 vccd1 vccd1 _14803_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15782_ _16169_/A _15782_/B vssd1 vssd1 vccd1 vccd1 _15839_/A sky130_fd_sc_hd__nand2_4
X_18570_ _19385_/CLK _18570_/D vssd1 vssd1 vccd1 vccd1 _18570_/Q sky130_fd_sc_hd__dfxtp_1
X_12994_ _12994_/A _13019_/C vssd1 vssd1 vccd1 vccd1 _12994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ _14544_/X _18823_/Q _14737_/S vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__mux2_1
X_17521_ _17521_/A vssd1 vssd1 vccd1 vccd1 _19710_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09312__A2 _09311_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ _11944_/A _12159_/B _12208_/A vssd1 vssd1 vccd1 vccd1 _12022_/A sky130_fd_sc_hd__o21ai_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17654_/B _17451_/X _17577_/S vssd1 vssd1 vccd1 vccd1 _17452_/X sky130_fd_sc_hd__mux2_1
XFILLER_45_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14664_ _14664_/A vssd1 vssd1 vccd1 vccd1 _18792_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _11876_/A _11876_/B vssd1 vssd1 vccd1 vccd1 _11877_/A sky130_fd_sc_hd__xor2_2
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _19450_/Q _16406_/C _16402_/X vssd1 vssd1 vccd1 vccd1 _16403_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13615_ _18384_/Q _13614_/X _13615_/S vssd1 vssd1 vccd1 vccd1 _13616_/A sky130_fd_sc_hd__mux2_1
X_17383_ _17732_/S vssd1 vssd1 vccd1 vccd1 _17648_/S sky130_fd_sc_hd__clkbuf_2
X_10827_ _09600_/A _10824_/X _10826_/X vssd1 vssd1 vccd1 vccd1 _10827_/X sky130_fd_sc_hd__a21o_1
X_14595_ _14595_/A vssd1 vssd1 vccd1 vccd1 _14595_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16334_ _16342_/D vssd1 vssd1 vccd1 vccd1 _16340_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_19122_ _19284_/CLK _19122_/D vssd1 vssd1 vccd1 vccd1 _19122_/Q sky130_fd_sc_hd__dfxtp_1
X_13546_ _13546_/A vssd1 vssd1 vccd1 vccd1 _18362_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16346__B1 _16293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10758_ _11305_/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10758_/X sky130_fd_sc_hd__or2_1
XFILLER_158_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19053_ _19245_/CLK _19053_/D vssd1 vssd1 vccd1 vccd1 _19053_/Q sky130_fd_sc_hd__dfxtp_1
X_16265_ _16265_/A vssd1 vssd1 vccd1 vccd1 _19402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13477_ _13138_/X _18338_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _13478_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14027__S _14027_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10689_ _10689_/A _10689_/B vssd1 vssd1 vccd1 vccd1 _10689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_139_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15216_ _15216_/A vssd1 vssd1 vccd1 vccd1 _19026_/D sky130_fd_sc_hd__clkbuf_1
X_18004_ _18004_/A vssd1 vssd1 vccd1 vccd1 _19774_/D sky130_fd_sc_hd__clkbuf_1
X_12428_ _12401_/Y _12381_/B _12427_/Y _17387_/B vssd1 vssd1 vccd1 vccd1 _12429_/B
+ sky130_fd_sc_hd__a31o_1
X_16196_ _13551_/X _19371_/Q _16202_/S vssd1 vssd1 vccd1 vccd1 _16197_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16750__B _16750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15147_ _15158_/A vssd1 vssd1 vccd1 vccd1 _15156_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_142_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _12360_/A _17885_/B vssd1 vssd1 vccd1 vccd1 _12388_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ _15078_/A vssd1 vssd1 vccd1 vccd1 _18968_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18906_ _19386_/CLK _18906_/D vssd1 vssd1 vccd1 vccd1 _18906_/Q sky130_fd_sc_hd__dfxtp_1
X_14029_ _14601_/A vssd1 vssd1 vccd1 vccd1 _14029_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12071__A _15632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10241__S0 _10450_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10697__A1 _10639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18837_ _19223_/CLK _18837_/D vssd1 vssd1 vccd1 vccd1 _18837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_132_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold16_A hold16/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10303__B _12468_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10792__S1 _10060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09570_ _10929_/A vssd1 vssd1 vccd1 vccd1 _09571_/A sky130_fd_sc_hd__clkbuf_2
X_18768_ _19319_/CLK _18768_/D vssd1 vssd1 vccd1 vccd1 _18768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18023__A0 _19783_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09380__A _09380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17719_ _11988_/A _17737_/A _17714_/X _17718_/Y _11539_/S vssd1 vssd1 vccd1 vccd1
+ _17719_/X sky130_fd_sc_hd__o221a_2
XFILLER_24_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18699_ _19319_/CLK _18699_/D vssd1 vssd1 vccd1 vccd1 _18699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16925__B _16929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17129__A2 _09096_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16337__B1 _16293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13776__S _13776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clock_A clock vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09906_ _18410_/Q _18671_/Q _18570_/Q _18905_/Q _09904_/X _09905_/X vssd1 vssd1 vccd1
+ vccd1 _09906_/X sky130_fd_sc_hd__mux4_1
XFILLER_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _09762_/X _09814_/X _09832_/X _09835_/X _09836_/Y vssd1 vssd1 vccd1 vccd1
+ _12478_/B sky130_fd_sc_hd__o32a_4
XFILLER_101_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_100_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09768_ _09768_/A vssd1 vssd1 vccd1 vccd1 _09769_/A sky130_fd_sc_hd__buf_2
XANTENNA__14400__S _14406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09699_ _10450_/S vssd1 vssd1 vccd1 vccd1 _09700_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A _17237_/A vssd1 vssd1 vccd1 vccd1 _11730_/X sky130_fd_sc_hd__and2_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11661_ _11708_/A vssd1 vssd1 vccd1 vccd1 _11810_/S sky130_fd_sc_hd__clkbuf_2
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13400_ _13400_/A vssd1 vssd1 vccd1 vccd1 _15629_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15231__S _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10612_ _10612_/A _10612_/B vssd1 vssd1 vccd1 vccd1 _10612_/X sky130_fd_sc_hd__or2_1
XANTENNA__16328__B1 _16293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14380_ _13848_/X _18680_/Q _14384_/S vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__mux2_1
X_11592_ _09171_/B _09211_/A _09211_/B _11586_/Y _11591_/X vssd1 vssd1 vccd1 vccd1
+ _11593_/S sky130_fd_sc_hd__a311o_1
XFILLER_168_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13330_/X _18311_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _13332_/A sky130_fd_sc_hd__mux2_1
X_10543_ _18926_/Q _18692_/Q _19374_/Q _19022_/Q _10763_/S _09590_/X vssd1 vssd1 vccd1
+ vccd1 _10544_/B sky130_fd_sc_hd__mux4_1
XFILLER_167_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11060__A _11208_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16050_ _16050_/A vssd1 vssd1 vccd1 vccd1 _19338_/D sky130_fd_sc_hd__clkbuf_1
X_13262_ _19481_/Q vssd1 vssd1 vccd1 vccd1 _16493_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_143_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ _19186_/Q _18800_/Q _19250_/Q _18369_/Q _10274_/A _10521_/A vssd1 vssd1 vccd1
+ vccd1 _10475_/B sky130_fd_sc_hd__mux4_1
XFILLER_109_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_160_clock clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 _19074_/CLK sky130_fd_sc_hd__clkbuf_16
X_15001_ _18944_/Q _14996_/X _15013_/S vssd1 vssd1 vccd1 vccd1 _15002_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12213_ _17820_/B _12214_/B vssd1 vssd1 vccd1 vccd1 _12242_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13686__S _13686_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ _13191_/X _18303_/Q _13252_/S vssd1 vssd1 vccd1 vccd1 _13194_/A sky130_fd_sc_hd__mux2_1
XFILLER_108_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09465__A _09465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12144_ _12170_/A _17222_/A vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_3_2_0_clock_A clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19740_ _19740_/CLK _19740_/D vssd1 vssd1 vccd1 vccd1 _19740_/Q sky130_fd_sc_hd__dfxtp_1
X_16952_ _15481_/X _16943_/X _16951_/X _16933_/X vssd1 vssd1 vccd1 vccd1 _19635_/D
+ sky130_fd_sc_hd__o211a_1
X_12075_ _13418_/A vssd1 vssd1 vccd1 vccd1 _12075_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_6_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_175_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19081_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_159_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15903_ _19287_/Q _14589_/A _15909_/S vssd1 vssd1 vccd1 vccd1 _15904_/A sky130_fd_sc_hd__mux2_1
X_11026_ _11026_/A _11026_/B vssd1 vssd1 vccd1 vccd1 _11026_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19671_ _19671_/CLK _19671_/D vssd1 vssd1 vccd1 vccd1 _19671_/Q sky130_fd_sc_hd__dfxtp_1
X_16883_ _16883_/A _16887_/C vssd1 vssd1 vccd1 vccd1 _16883_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11340__A2 _11329_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10774__S1 _10060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18622_ _19085_/CLK _18622_/D vssd1 vssd1 vccd1 vccd1 _18622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15834_ _15834_/A vssd1 vssd1 vccd1 vccd1 _19256_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14310__S _14310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11628__B1 _11840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18553_ _18824_/CLK _18553_/D vssd1 vssd1 vccd1 vccd1 _18553_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09916__S0 _10114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15765_ _13592_/X _19226_/Q _15765_/S vssd1 vssd1 vccd1 vccd1 _15766_/A sky130_fd_sc_hd__mux2_1
X_12977_ _12977_/A vssd1 vssd1 vccd1 vccd1 _12977_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13093__A2 _12974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17500_/X _17503_/X _17504_/S vssd1 vssd1 vccd1 vccd1 _17505_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ _11928_/A _17201_/A vssd1 vssd1 vccd1 vccd1 _11929_/B sky130_fd_sc_hd__and2_1
X_14716_ _14772_/A vssd1 vssd1 vccd1 vccd1 _14785_/S sky130_fd_sc_hd__buf_6
XFILLER_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18484_ _19012_/CLK _18484_/D vssd1 vssd1 vccd1 vccd1 _18484_/Q sky130_fd_sc_hd__dfxtp_1
X_15696_ _14601_/X _19195_/Q _15704_/S vssd1 vssd1 vccd1 vccd1 _15697_/A sky130_fd_sc_hd__mux2_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17435_ _17446_/S _17435_/B vssd1 vssd1 vccd1 vccd1 _17435_/X sky130_fd_sc_hd__or2_1
X_14647_ _14647_/A vssd1 vssd1 vccd1 vccd1 _18784_/D sky130_fd_sc_hd__clkbuf_1
X_11859_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11859_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_61_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16237__S _16239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15141__S _15145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18018__A _18029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13450__A _13507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14578_ _14578_/A vssd1 vssd1 vccd1 vccd1 _18764_/D sky130_fd_sc_hd__clkbuf_1
X_17366_ _17294_/S _17275_/X _17365_/X vssd1 vssd1 vccd1 vccd1 _17506_/B sky130_fd_sc_hd__a21oi_1
XFILLER_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19105_ _19267_/CLK _19105_/D vssd1 vssd1 vccd1 vccd1 _19105_/Q sky130_fd_sc_hd__dfxtp_1
X_16317_ _19481_/Q _19483_/Q _19482_/Q _16486_/A vssd1 vssd1 vccd1 vccd1 _16496_/A
+ sky130_fd_sc_hd__and4_1
X_13529_ _18357_/Q _13528_/X _13529_/S vssd1 vssd1 vccd1 vccd1 _13530_/A sky130_fd_sc_hd__mux2_1
XFILLER_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17297_ _17456_/S vssd1 vssd1 vccd1 vccd1 _17615_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16761__A _19562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12066__A _12066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16248_ _16248_/A vssd1 vssd1 vccd1 vccd1 _19394_/D sky130_fd_sc_hd__clkbuf_1
X_19036_ _19388_/CLK _19036_/D vssd1 vssd1 vccd1 vccd1 _19036_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_128_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19356_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_127_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput103 _09096_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[0] sky130_fd_sc_hd__buf_2
X_16179_ _16179_/A vssd1 vssd1 vccd1 vccd1 _19363_/D sky130_fd_sc_hd__clkbuf_1
Xoutput114 _12461_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[14] sky130_fd_sc_hd__buf_2
XANTENNA__14281__A _14281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput125 _12473_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[24] sky130_fd_sc_hd__buf_2
Xoutput136 _12448_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[5] sky130_fd_sc_hd__buf_2
Xoutput147 _16274_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[14] sky130_fd_sc_hd__buf_2
XFILLER_115_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09375__A _18780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput158 _12279_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[24] sky130_fd_sc_hd__buf_2
XANTENNA__10462__S0 _10499_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput169 _16253_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[5] sky130_fd_sc_hd__buf_2
XFILLER_114_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12513__B _12536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12108__A1 _18114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11316__C1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09622_ _18641_/Q vssd1 vssd1 vccd1 vccd1 _10969_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09553_ _09553_/A vssd1 vssd1 vccd1 vccd1 _09658_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11095__B2 _12447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09484_ _09484_/A vssd1 vssd1 vccd1 vccd1 _09485_/A sky130_fd_sc_hd__buf_2
XFILLER_52_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15986__S _15992_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16671__A _16714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16730__B1 _19553_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_139_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12704__A _13009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11555__C1 _18104_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19549_/CLK sky130_fd_sc_hd__clkbuf_16
X_10190_ _18406_/Q _18667_/Q _18566_/Q _18901_/Q _09868_/A _09927_/A vssd1 vssd1 vccd1
+ vccd1 _10191_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14639__A3 _18029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_160_clock_A clkbuf_4_8_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12900_ _19525_/Q _12782_/X _12699_/X _16540_/B _12899_/X vssd1 vssd1 vccd1 vccd1
+ _12900_/X sky130_fd_sc_hd__a221o_1
XANTENNA__15226__S _15228_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10756__S1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_101_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13535__A _15019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13880_ _14560_/A vssd1 vssd1 vccd1 vccd1 _13880_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14130__S _14136_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12831_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12831_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10508__S1 _09710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11055__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15550_ _15519_/X _15546_/X _15548_/Y _15549_/X hold10/X vssd1 vssd1 vccd1 vccd1
+ _15550_/X sky130_fd_sc_hd__a32o_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12769_/A vssd1 vssd1 vccd1 vccd1 _12762_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_30_clock clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19291_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14501_ _14501_/A vssd1 vssd1 vccd1 vccd1 _18734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _17183_/A _11713_/B _17177_/A _11566_/X vssd1 vssd1 vccd1 vccd1 _12050_/A
+ sky130_fd_sc_hd__or4b_4
X_15481_ _15478_/X _15479_/X _15480_/Y _13403_/X _18255_/Q vssd1 vssd1 vccd1 vccd1
+ _15481_/X sky130_fd_sc_hd__a32o_4
XANTENNA__10833__B2 _19715_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _18121_/A vssd1 vssd1 vccd1 vccd1 _18142_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_15_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17220_ _17709_/B _17779_/B _17263_/A vssd1 vssd1 vccd1 vccd1 _17220_/X sky130_fd_sc_hd__mux2_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14432_ _14432_/A vssd1 vssd1 vccd1 vccd1 _18703_/D sky130_fd_sc_hd__clkbuf_1
X_11644_ _12392_/S _11644_/B vssd1 vssd1 vccd1 vccd1 _11644_/Y sky130_fd_sc_hd__nand2_1
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15896__S _15898_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17151_ _17160_/A _17151_/B vssd1 vssd1 vccd1 vccd1 _17152_/A sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_45_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19120_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17677__A _17917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14363_ _13931_/X _18674_/Q _14365_/S vssd1 vssd1 vccd1 vccd1 _14364_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_155_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_85_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _11575_/A _11575_/B _17183_/C _17174_/B vssd1 vssd1 vccd1 vccd1 _11575_/X
+ sky130_fd_sc_hd__or4_1
Xinput16 io_dbus_rdata[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_2
Xinput27 io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_2
XFILLER_128_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16102_ _16102_/A vssd1 vssd1 vccd1 vccd1 _19347_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput38 io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09894__S _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13314_ input21/X _13134_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _13314_/X sky130_fd_sc_hd__a21o_1
Xinput49 io_ibus_inst[23] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_2
X_17082_ _17082_/A vssd1 vssd1 vccd1 vccd1 _19687_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15524__A1 _15522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10526_ _10531_/A _10526_/B vssd1 vssd1 vccd1 vccd1 _10526_/Y sky130_fd_sc_hd__nor2_1
XFILLER_156_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14294_ input50/X _14282_/X _14293_/X _14278_/X _18130_/A vssd1 vssd1 vccd1 vccd1
+ _18224_/B sky130_fd_sc_hd__a32o_2
XFILLER_109_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_143_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16033_ _16031_/X _19335_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15197__A _15243_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13245_ _13245_/A _13256_/C vssd1 vssd1 vccd1 vccd1 _13245_/Y sky130_fd_sc_hd__nand2_1
X_10457_ _10514_/A _10457_/B vssd1 vssd1 vccd1 vccd1 _10457_/X sky130_fd_sc_hd__or2_1
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12614__A _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09195__A _19811_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13429__B _17023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ _19759_/Q _13176_/B vssd1 vssd1 vccd1 vccd1 _13213_/C sky130_fd_sc_hd__and2_1
X_10388_ _10297_/X _10378_/Y _10383_/X _10387_/Y _09812_/A vssd1 vssd1 vccd1 vccd1
+ _10388_/X sky130_fd_sc_hd__o311a_4
XFILLER_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11561__A2 _18102_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12127_ _12322_/A _12322_/B _12127_/C _12127_/D vssd1 vssd1 vccd1 vccd1 _12127_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_97_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17984_ _16142_/A _19797_/Q _17990_/S vssd1 vssd1 vccd1 vccd1 _17985_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19723_ _19725_/CLK _19723_/D vssd1 vssd1 vccd1 vccd1 _19723_/Q sky130_fd_sc_hd__dfxtp_2
X_16935_ _16935_/A _16931_/X vssd1 vssd1 vccd1 vccd1 _16935_/X sky130_fd_sc_hd__or2b_1
X_12058_ _12008_/A _12008_/B _12034_/A _12057_/Y vssd1 vssd1 vccd1 vccd1 _12059_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11009_ _18454_/Q _19045_/Q _19207_/Q _18422_/Q _10940_/S _11005_/X vssd1 vssd1 vccd1
+ vccd1 _11010_/B sky130_fd_sc_hd__mux4_1
XFILLER_42_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19654_ _19660_/CLK _19654_/D vssd1 vssd1 vccd1 vccd1 _19654_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14040__S _14043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16866_ _16883_/A _16871_/C vssd1 vssd1 vccd1 vccd1 _16866_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18605_ _19264_/CLK _18605_/D vssd1 vssd1 vccd1 vccd1 _18605_/Q sky130_fd_sc_hd__dfxtp_1
X_15817_ _15839_/A vssd1 vssd1 vccd1 vccd1 _15826_/S sky130_fd_sc_hd__buf_6
XFILLER_19_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19585_ _19671_/CLK _19585_/D vssd1 vssd1 vccd1 vccd1 _19585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16797_ _16800_/B _16800_/C _19573_/Q vssd1 vssd1 vccd1 vccd1 _16799_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18536_ _19291_/CLK _18536_/D vssd1 vssd1 vccd1 vccd1 _18536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ _13567_/X _19218_/Q _15754_/S vssd1 vssd1 vccd1 vccd1 _15749_/A sky130_fd_sc_hd__mux2_1
XFILLER_80_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18467_ _19058_/CLK _18467_/D vssd1 vssd1 vccd1 vccd1 _18467_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15679_ _15679_/A vssd1 vssd1 vccd1 vccd1 _19187_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17418_ _17468_/A _17418_/B vssd1 vssd1 vccd1 vccd1 _17418_/Y sky130_fd_sc_hd__nand2_1
X_18398_ _19309_/CLK _18398_/D vssd1 vssd1 vccd1 vccd1 _18398_/Q sky130_fd_sc_hd__dfxtp_1
X_17349_ _17345_/Y _17347_/Y _17497_/S vssd1 vssd1 vccd1 vccd1 _17350_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10588__B1 _09630_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10683__S0 _10576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15515__B2 hold18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12329__A1 _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19019_ _19278_/CLK _19019_/D vssd1 vssd1 vccd1 vccd1 _19019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_162_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12524__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09833__A _09833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_84_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09605_ _19200_/Q _18814_/Q _19264_/Q _18383_/Q _10603_/S _10669_/A vssd1 vssd1 vccd1
+ vccd1 _09606_/B sky130_fd_sc_hd__mux4_1
XFILLER_84_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__C _12956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14885__S _14893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16666__A _16666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11068__A1 _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _10579_/A vssd1 vssd1 vccd1 vccd1 _10631_/S sky130_fd_sc_hd__buf_4
XFILLER_24_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11163__S1 _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ _09726_/A _09454_/X _09456_/X _09462_/X _09752_/A vssd1 vssd1 vccd1 vccd1
+ _09467_/X sky130_fd_sc_hd__a311o_4
XFILLER_24_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13090__A _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09398_ _11299_/S vssd1 vssd1 vccd1 vccd1 _10603_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__12568__A1 _19627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11360_ _11423_/A _11360_/B _11422_/A _11431_/C vssd1 vssd1 vccd1 vccd1 _11361_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10311_ _10311_/A vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__buf_4
XFILLER_138_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11291_ _11291_/A _12453_/A vssd1 vssd1 vccd1 vccd1 _11292_/B sky130_fd_sc_hd__or2_1
XFILLER_138_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13030_ _16055_/A _13031_/B _13113_/C vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__10426__S0 _10339_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10242_ _10406_/A _10242_/B vssd1 vssd1 vccd1 vccd1 _10242_/X sky130_fd_sc_hd__or2_1
XFILLER_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15745__A _15767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10173_ _18407_/Q _18668_/Q _18567_/Q _18902_/Q _09904_/X _09905_/X vssd1 vssd1 vccd1
+ vccd1 _10174_/B sky130_fd_sc_hd__mux4_1
XFILLER_105_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input38_A io_ibus_inst[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14981_ _14981_/A vssd1 vssd1 vccd1 vccd1 _18936_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_5_0_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_5_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
X_16720_ _16724_/C _16724_/D _16719_/Y vssd1 vssd1 vccd1 vccd1 _19549_/D sky130_fd_sc_hd__o21a_1
X_13932_ _13931_/X _18509_/Q _13935_/S vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16651_ _16660_/A _16651_/B _16663_/D vssd1 vssd1 vccd1 vccd1 _19527_/D sky130_fd_sc_hd__nor3_1
X_13863_ _13863_/A vssd1 vssd1 vccd1 vccd1 _18487_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17431__B2 _17430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14795__S _14799_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10401__B _12466_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15602_ _19732_/Q _15600_/X _15626_/S vssd1 vssd1 vccd1 vccd1 _15602_/X sky130_fd_sc_hd__mux2_1
X_12814_ _12814_/A vssd1 vssd1 vccd1 vccd1 _18283_/D sky130_fd_sc_hd__clkbuf_1
X_19370_ _19370_/CLK _19370_/D vssd1 vssd1 vccd1 vccd1 _19370_/Q sky130_fd_sc_hd__dfxtp_1
X_16582_ _19508_/Q _16584_/C _16581_/Y vssd1 vssd1 vccd1 vccd1 _19508_/D sky130_fd_sc_hd__o21a_1
X_13794_ _13048_/X _18461_/Q _13798_/S vssd1 vssd1 vccd1 vccd1 _13795_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17719__C1 _11539_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16295__B _16295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11154__S1 _11033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18321_ _19202_/CLK _18321_/D vssd1 vssd1 vccd1 vccd1 _18321_/Q sky130_fd_sc_hd__dfxtp_1
X_15533_ _15533_/A vssd1 vssd1 vccd1 vccd1 _19150_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ hold12/A _12744_/X _11291_/A _12740_/X vssd1 vssd1 vccd1 vccd1 _18259_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _15603_/A vssd1 vssd1 vccd1 vccd1 _15636_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18252_ _19799_/CLK _18252_/D vssd1 vssd1 vccd1 vccd1 _18252_/Q sky130_fd_sc_hd__dfxtp_2
X_12676_ _19543_/Q vssd1 vssd1 vccd1 vccd1 _16706_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14415_ _13899_/X _18696_/Q _14417_/S vssd1 vssd1 vccd1 vccd1 _14416_/A sky130_fd_sc_hd__mux2_1
X_17203_ _17203_/A vssd1 vssd1 vccd1 vccd1 _17263_/A sky130_fd_sc_hd__clkbuf_2
X_11627_ _11670_/A _12443_/B _11600_/Y vssd1 vssd1 vccd1 vccd1 _17225_/A sky130_fd_sc_hd__o21ai_1
XFILLER_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18183_ _18190_/A _18183_/B vssd1 vssd1 vccd1 vccd1 _18184_/A sky130_fd_sc_hd__and2_1
X_15395_ _15395_/A vssd1 vssd1 vccd1 vccd1 _19105_/D sky130_fd_sc_hd__clkbuf_1
X_14346_ _13905_/X _18666_/Q _14354_/S vssd1 vssd1 vccd1 vccd1 _14347_/A sky130_fd_sc_hd__mux2_1
X_17134_ _17114_/A _17115_/X _17149_/A _17140_/A _15612_/X vssd1 vssd1 vccd1 vccd1
+ _17135_/B sky130_fd_sc_hd__a32o_1
XANTENNA__09918__A _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11558_ _17174_/A _17166_/C vssd1 vssd1 vccd1 vccd1 _11562_/C sky130_fd_sc_hd__or2_1
XFILLER_156_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17065_ _17065_/A vssd1 vssd1 vccd1 vccd1 _19679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10509_ _10509_/A _10509_/B vssd1 vssd1 vccd1 vccd1 _10509_/X sky130_fd_sc_hd__or2_1
X_14277_ _18229_/A vssd1 vssd1 vccd1 vccd1 _14277_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_144_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11489_ _11491_/B _11489_/B _11489_/C vssd1 vssd1 vccd1 vccd1 _11495_/B sky130_fd_sc_hd__or3_1
XFILLER_170_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16016_ _16016_/A vssd1 vssd1 vccd1 vccd1 _19332_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13228_ _14592_/A vssd1 vssd1 vccd1 vccd1 _13228_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_171_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17854__B _17856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__B _12063_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_97_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12731__A1 _18253_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _19571_/Q _12518_/X _13158_/X _12538_/X vssd1 vssd1 vccd1 vccd1 _13159_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_124_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11090__S0 _10969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17670__A1 _11904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17967_ _17967_/A vssd1 vssd1 vccd1 vccd1 _19757_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10799__A _18780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19706_ _19706_/CLK _19706_/D vssd1 vssd1 vccd1 vccd1 _19706_/Q sky130_fd_sc_hd__dfxtp_1
X_16918_ _16520_/B _16915_/B _16917_/Y vssd1 vssd1 vccd1 vccd1 _19619_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09586__S1 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17898_ _17896_/X _17897_/Y _17898_/S vssd1 vssd1 vccd1 vccd1 _17898_/X sky130_fd_sc_hd__mux2_1
XFILLER_168_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19637_ _19669_/CLK _19637_/D vssd1 vssd1 vccd1 vccd1 _19637_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16849_ _16849_/A vssd1 vssd1 vccd1 vccd1 _16854_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15390__A _15446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19568_ _19668_/CLK _19568_/D vssd1 vssd1 vccd1 vccd1 _19568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09321_ _12720_/A vssd1 vssd1 vccd1 vccd1 _17994_/S sky130_fd_sc_hd__clkbuf_2
X_18519_ _19367_/CLK _18519_/D vssd1 vssd1 vccd1 vccd1 _18519_/Q sky130_fd_sc_hd__dfxtp_1
X_19499_ _19502_/CLK _19499_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__09663__A1 _11418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ _19830_/Q _19828_/Q _19827_/Q _19829_/Q vssd1 vssd1 vccd1 vccd1 _09253_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09183_ _19849_/Q _19848_/Q _09186_/A vssd1 vssd1 vccd1 vccd1 _11574_/A sky130_fd_sc_hd__or3_2
XANTENNA__10656__S0 _10729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_107_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11081__S0 _10969_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17661__A1 _17662_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11289__A1 _10895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11289__B2 _12448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10860_ _18585_/Q _18856_/Q _19080_/Q _18824_/Q _09626_/A _10855_/A vssd1 vssd1 vccd1
+ vccd1 _10860_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09519_ _09519_/A vssd1 vssd1 vccd1 vccd1 _10017_/S sky130_fd_sc_hd__buf_4
XFILLER_17_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _11331_/A _10791_/B vssd1 vssd1 vccd1 vccd1 _10791_/Y sky130_fd_sc_hd__nor2_1
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _13391_/A _13391_/B vssd1 vssd1 vccd1 vccd1 _12677_/A sky130_fd_sc_hd__nor2_1
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ _12461_/A _12461_/B vssd1 vssd1 vccd1 vccd1 _12461_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14644__A _14700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18116__A _18116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ _14268_/S vssd1 vssd1 vccd1 vccd1 _14209_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_166_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11213__A1 _11007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11412_ _11412_/A _11492_/C vssd1 vssd1 vccd1 vccd1 _11420_/A sky130_fd_sc_hd__and2_2
X_15180_ _19010_/Q _15006_/X _15184_/S vssd1 vssd1 vccd1 vccd1 _15181_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12392_ _12391_/X _12389_/Y _12392_/S vssd1 vssd1 vccd1 vccd1 _12392_/X sky130_fd_sc_hd__mux2_1
XFILLER_165_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12961__A1 _16760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ _14131_/A vssd1 vssd1 vccd1 vccd1 _18578_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12961__B2 _16963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ _11343_/A _11342_/Y vssd1 vssd1 vccd1 vccd1 _11344_/A sky130_fd_sc_hd__or2b_1
XFILLER_153_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14062_ _14062_/A vssd1 vssd1 vccd1 vccd1 _18548_/D sky130_fd_sc_hd__clkbuf_1
X_11274_ _11278_/A _11274_/B vssd1 vssd1 vccd1 vccd1 _11274_/Y sky130_fd_sc_hd__nor2_1
XFILLER_140_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13013_ _19562_/Q _13006_/X _13011_/X _13012_/X vssd1 vssd1 vccd1 vccd1 _13013_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_152_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13910__A0 _13909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10225_ _19728_/Q vssd1 vssd1 vccd1 vccd1 _10225_/Y sky130_fd_sc_hd__inv_2
X_18870_ _19088_/CLK _18870_/D vssd1 vssd1 vccd1 vccd1 _18870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17821_ _17765_/A _17819_/B _17800_/A _17820_/X vssd1 vssd1 vccd1 vccd1 _17821_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10156_ _09667_/X _10146_/X _10155_/X _09758_/X _19729_/Q vssd1 vssd1 vccd1 vccd1
+ _10181_/A sky130_fd_sc_hd__a32o_4
XFILLER_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17752_ _17756_/B _12089_/X vssd1 vssd1 vccd1 vccd1 _17752_/X sky130_fd_sc_hd__or2b_1
XFILLER_48_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14964_ _18928_/Q vssd1 vssd1 vccd1 vccd1 _14965_/A sky130_fd_sc_hd__clkbuf_1
X_10087_ _10087_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _10088_/B sky130_fd_sc_hd__or2_1
XFILLER_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16703_ _16706_/C _16706_/D _19544_/Q vssd1 vssd1 vccd1 vccd1 _16705_/B sky130_fd_sc_hd__a21oi_1
X_13915_ _14595_/A vssd1 vssd1 vccd1 vccd1 _13915_/X sky130_fd_sc_hd__clkbuf_2
X_17683_ _17673_/X _17675_/X _17682_/Y vssd1 vssd1 vccd1 vccd1 _17683_/Y sky130_fd_sc_hd__o21ai_1
X_14895_ _14917_/A vssd1 vssd1 vccd1 vccd1 _14904_/S sky130_fd_sc_hd__buf_4
XFILLER_75_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19422_ _19423_/CLK _19422_/D vssd1 vssd1 vccd1 vccd1 _19422_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__15414__S _15422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16634_ _19522_/Q _16634_/B _16659_/B vssd1 vssd1 vccd1 vccd1 _16635_/B sky130_fd_sc_hd__and3_1
X_13846_ _13845_/X _18482_/Q _13855_/S vssd1 vssd1 vccd1 vccd1 _13847_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19353_ _19357_/CLK _19353_/D vssd1 vssd1 vccd1 vccd1 _19353_/Q sky130_fd_sc_hd__dfxtp_1
X_16565_ hold1/A _16567_/C _16564_/Y vssd1 vssd1 vccd1 vccd1 _19502_/D sky130_fd_sc_hd__o21a_1
X_13777_ _13777_/A vssd1 vssd1 vccd1 vccd1 _18453_/D sky130_fd_sc_hd__clkbuf_1
X_10989_ _18614_/Q _18949_/Q _11241_/S vssd1 vssd1 vccd1 vccd1 _10990_/B sky130_fd_sc_hd__mux2_1
XFILLER_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18304_ _19287_/CLK _18304_/D vssd1 vssd1 vccd1 vccd1 _18304_/Q sky130_fd_sc_hd__dfxtp_1
X_15516_ _19716_/Q _15515_/X _15516_/S vssd1 vssd1 vccd1 vccd1 _15516_/X sky130_fd_sc_hd__mux2_1
X_19284_ _19284_/CLK _19284_/D vssd1 vssd1 vccd1 vccd1 _19284_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10886__S0 _11172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12728_ _12751_/A _12730_/C vssd1 vssd1 vccd1 vccd1 _12769_/A sky130_fd_sc_hd__nor2_4
X_16496_ _16496_/A vssd1 vssd1 vccd1 vccd1 _16501_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18235_ input53/X _18197_/X _18229_/X _18234_/X _18138_/A vssd1 vssd1 vccd1 vccd1
+ _18236_/B sky130_fd_sc_hd__a32o_1
X_12659_ _13008_/A vssd1 vssd1 vccd1 vccd1 _12659_/X sky130_fd_sc_hd__clkbuf_2
X_15447_ _19129_/Q _15079_/X _15455_/S vssd1 vssd1 vccd1 vccd1 _15448_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14554__A _14621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11204__A1 _11007_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09648__A _10586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18166_ _18170_/A _18166_/B vssd1 vssd1 vccd1 vccd1 _18167_/A sky130_fd_sc_hd__and2_1
XFILLER_8_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10638__S0 _10576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15378_ _15378_/A vssd1 vssd1 vccd1 vccd1 _19098_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17117_ _17117_/A _17117_/B vssd1 vssd1 vccd1 vccd1 _17175_/B sky130_fd_sc_hd__nor2_1
XFILLER_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14329_ _14329_/A vssd1 vssd1 vccd1 vccd1 _18658_/D sky130_fd_sc_hd__clkbuf_1
X_18097_ _18097_/A vssd1 vssd1 vccd1 vccd1 _18097_/X sky130_fd_sc_hd__buf_2
X_17048_ _19672_/Q _15509_/X _17050_/S vssd1 vssd1 vccd1 vccd1 _17049_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_143_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ _09927_/A vssd1 vssd1 vccd1 vccd1 _09871_/A sky130_fd_sc_hd__clkbuf_4
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11063__S0 _11011_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10715__B1 _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__B1 _09833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__S0 _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18999_ _19127_/CLK _18999_/D vssd1 vssd1 vccd1 vccd1 _18999_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15654__A0 _14541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13109__S _13172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11418__A _11418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15324__S _15328_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13633__A _13690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17159__B1 _17140_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09304_ _19702_/Q vssd1 vssd1 vccd1 vccd1 _09305_/A sky130_fd_sc_hd__inv_2
XFILLER_55_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09235_ _13400_/A _09235_/B _09234_/X vssd1 vssd1 vccd1 vccd1 _09235_/X sky130_fd_sc_hd__or3b_1
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18108__C1 _18097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _09166_/A _09166_/B _09176_/B vssd1 vssd1 vccd1 vccd1 _09208_/A sky130_fd_sc_hd__or3b_2
XFILLER_163_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12943__A1 input30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15994__S _15996_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ _19838_/Q vssd1 vssd1 vccd1 vccd1 _18077_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_162_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11054__S0 _11241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10010_ _18475_/Q _19066_/Q _19228_/Q _18443_/Q _09539_/A _09543_/A vssd1 vssd1 vccd1
+ vccd1 _10010_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09999_ _19292_/Q _19130_/Q _18539_/Q _18309_/Q _09850_/A _09671_/A vssd1 vssd1 vccd1
+ vccd1 _09999_/X sky130_fd_sc_hd__mux4_1
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11961_ _19404_/Q vssd1 vssd1 vccd1 vccd1 _11969_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_151_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13700_ _13700_/A vssd1 vssd1 vccd1 vccd1 _18419_/D sky130_fd_sc_hd__clkbuf_1
X_10912_ _10961_/A _10912_/B vssd1 vssd1 vccd1 vccd1 _10912_/Y sky130_fd_sc_hd__nor2_1
X_14680_ _14680_/A vssd1 vssd1 vccd1 vccd1 _18799_/D sky130_fd_sc_hd__clkbuf_1
X_11892_ _11892_/A vssd1 vssd1 vccd1 vccd1 _17662_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16070__A0 _15542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13631_ _12886_/X _18389_/Q _13631_/S vssd1 vssd1 vccd1 vccd1 _13632_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10843_ _10848_/A _10843_/B vssd1 vssd1 vccd1 vccd1 _10843_/Y sky130_fd_sc_hd__nor2_1
XFILLER_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16350_ _16351_/B _16351_/C _19433_/Q vssd1 vssd1 vccd1 vccd1 _16352_/B sky130_fd_sc_hd__a21oi_1
X_13562_ _13562_/A vssd1 vssd1 vccd1 vccd1 _18367_/D sky130_fd_sc_hd__clkbuf_1
X_10774_ _19179_/Q _18793_/Q _19243_/Q _18362_/Q _10633_/S _10060_/A vssd1 vssd1 vccd1
+ vccd1 _10775_/B sky130_fd_sc_hd__mux4_1
XFILLER_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12513_ _12600_/B _12536_/B vssd1 vssd1 vccd1 vccd1 _12962_/A sky130_fd_sc_hd__or2_1
X_15301_ _15301_/A vssd1 vssd1 vccd1 vccd1 _19064_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16281_ _12066_/B _16278_/X _12073_/Y _12079_/Y _16280_/X vssd1 vssd1 vccd1 vccd1
+ _19408_/D sky130_fd_sc_hd__o221a_1
XFILLER_13_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13493_ _13493_/A vssd1 vssd1 vccd1 vccd1 _18345_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14384__A0 _13854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18020_ _18020_/A vssd1 vssd1 vccd1 vccd1 _19781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_173_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12444_ _12447_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _12444_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09468__A _09468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15232_ _15232_/A vssd1 vssd1 vccd1 vccd1 _19033_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12606__B _12606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_154_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12934__A1 _19335_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12934__B2 _19145_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ _19003_/Q _15086_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15164_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12375_ _12233_/X _12367_/Y _12368_/X _12078_/A _12374_/X vssd1 vssd1 vccd1 vccd1
+ _12375_/X sky130_fd_sc_hd__o311a_1
XFILLER_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14114_ _13928_/X _18572_/Q _14118_/S vssd1 vssd1 vccd1 vccd1 _14115_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11326_ _11331_/A _11326_/B vssd1 vssd1 vccd1 vccd1 _11326_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17873__A1 _17872_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15094_ _15094_/A vssd1 vssd1 vccd1 vccd1 _18973_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18922_ _19370_/CLK _18922_/D vssd1 vssd1 vccd1 vccd1 _18922_/Q sky130_fd_sc_hd__dfxtp_1
X_14045_ _14617_/A vssd1 vssd1 vccd1 vccd1 _14045_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11257_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11257_/X sky130_fd_sc_hd__or2_1
X_10208_ _18470_/Q _19061_/Q _19223_/Q _18438_/Q _09955_/S _09905_/A vssd1 vssd1 vccd1
+ vccd1 _10209_/B sky130_fd_sc_hd__mux4_1
XFILLER_68_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18853_ _19365_/CLK _18853_/D vssd1 vssd1 vccd1 vccd1 _18853_/Q sky130_fd_sc_hd__dfxtp_1
X_11188_ _11188_/A _11188_/B vssd1 vssd1 vccd1 vccd1 _11188_/X sky130_fd_sc_hd__or2_1
XFILLER_68_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11370__B1 _09740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17804_ _17673_/A _17801_/X _17803_/X _17633_/A vssd1 vssd1 vccd1 vccd1 _17804_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10139_ _18631_/Q _18966_/Q _10185_/S vssd1 vssd1 vccd1 vccd1 _10139_/X sky130_fd_sc_hd__mux2_1
X_18784_ _19203_/CLK _18784_/D vssd1 vssd1 vccd1 vccd1 _18784_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15996_ _13614_/X _19329_/Q _15996_/S vssd1 vssd1 vccd1 vccd1 _15997_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17735_ _19721_/Q _17734_/X _17873_/S vssd1 vssd1 vccd1 vccd1 _17736_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14947_ _14947_/A vssd1 vssd1 vccd1 vccd1 _18919_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18050__A1 _19416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17666_ _17659_/X _17663_/X _17665_/X vssd1 vssd1 vccd1 vccd1 _17666_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14878_ _18887_/Q _13972_/X _14882_/S vssd1 vssd1 vccd1 vccd1 _14879_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19405_ _19807_/CLK _19405_/D vssd1 vssd1 vccd1 vccd1 _19405_/Q sky130_fd_sc_hd__dfxtp_1
X_16617_ _19519_/Q _16614_/B _16616_/Y vssd1 vssd1 vccd1 vccd1 _19519_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ _13330_/X _18477_/Q _13831_/S vssd1 vssd1 vccd1 vccd1 _13830_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17597_ _17597_/A vssd1 vssd1 vccd1 vccd1 _17597_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16764__A _16812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19336_ _19356_/CLK _19336_/D vssd1 vssd1 vccd1 vccd1 _19336_/Q sky130_fd_sc_hd__dfxtp_2
X_16548_ _16551_/B _16551_/C _16547_/Y vssd1 vssd1 vccd1 vccd1 _19496_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19267_ _19267_/CLK _19267_/D vssd1 vssd1 vccd1 vccd1 _19267_/Q sky130_fd_sc_hd__dfxtp_1
X_16479_ _16524_/A _16483_/C vssd1 vssd1 vccd1 vccd1 _16479_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14284__A _14290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18218_ _18224_/A _18218_/B vssd1 vssd1 vccd1 vccd1 _18219_/A sky130_fd_sc_hd__and2_1
XANTENNA__09378__A _09416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19198_ _19388_/CLK _19198_/D vssd1 vssd1 vccd1 vccd1 _19198_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18105__A2 _18086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12516__B _12536_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18149_ _09236_/D _12674_/A _18148_/Y input34/X vssd1 vssd1 vccd1 vccd1 _18150_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_144_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_160_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09922_ _09890_/A _09921_/X _09767_/A vssd1 vssd1 vccd1 vccd1 _09922_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11036__S0 _11149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14223__S _14231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09853_ _10368_/S vssd1 vssd1 vccd1 vccd1 _10367_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_113_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10164__A1 _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10052__A _10684_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ _09784_/A vssd1 vssd1 vccd1 vccd1 _09784_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09841__A _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16052__A0 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14893__S _14893_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09609__A1 _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13405__A2 _13404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09218_ _19859_/Q _09347_/B vssd1 vssd1 vccd1 vccd1 _09223_/B sky130_fd_sc_hd__nor2_1
XFILLER_127_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _09764_/A _10483_/X _10485_/Y _10489_/Y _09812_/A vssd1 vssd1 vccd1 vccd1
+ _10490_/X sky130_fd_sc_hd__o311a_4
XFILLER_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12916__A1 _16752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09149_ _11530_/A _11587_/A vssd1 vssd1 vccd1 vccd1 _11577_/B sky130_fd_sc_hd__nor2_1
XFILLER_136_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11275__S0 _11071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__A _11354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12160_ _09351_/A _11507_/A _12209_/A vssd1 vssd1 vccd1 vccd1 _12160_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_162_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11111_ _11111_/A _11111_/B vssd1 vssd1 vccd1 vccd1 _11111_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_2_2_0_clock_A clkbuf_2_3_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11027__S0 _11149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13538__A _15022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12091_ _12091_/A _12091_/B vssd1 vssd1 vccd1 vccd1 _12092_/A sky130_fd_sc_hd__xnor2_1
XFILLER_146_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11042_ _11042_/A vssd1 vssd1 vccd1 vccd1 _11042_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_104_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15850_ _13611_/X _19264_/Q _15852_/S vssd1 vssd1 vccd1 vccd1 _15851_/A sky130_fd_sc_hd__mux2_1
X_14801_ _14858_/S vssd1 vssd1 vccd1 vccd1 _14810_/S sky130_fd_sc_hd__buf_2
XFILLER_58_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input20_A io_dbus_rdata[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15781_ _15781_/A vssd1 vssd1 vccd1 vccd1 _19233_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12993_ _19748_/Q vssd1 vssd1 vccd1 vccd1 _12994_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_92_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17520_ _19710_/Q _17519_/X _17520_/S vssd1 vssd1 vccd1 vccd1 _17521_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18032__A1 _12066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13273__A _15079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__A1 _19330_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14732_ _14732_/A vssd1 vssd1 vccd1 vccd1 _18822_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11944_ _11944_/A vssd1 vssd1 vccd1 vccd1 _12021_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17448_/X _17449_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17451_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14663_ _14547_/X _18792_/Q _14665_/S vssd1 vssd1 vccd1 vccd1 _14664_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11875_ _11854_/A _11854_/B _11848_/A vssd1 vssd1 vccd1 vccd1 _11876_/B sky130_fd_sc_hd__a21oi_1
XFILLER_72_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output107_A _12482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16402_ _16546_/A vssd1 vssd1 vccd1 vccd1 _16402_/X sky130_fd_sc_hd__buf_2
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10826_ _09394_/A _10825_/X _10953_/A vssd1 vssd1 vccd1 vccd1 _10826_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11407__A1 _09823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13614_ _15098_/A vssd1 vssd1 vccd1 vccd1 _13614_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__12604__B1 _12603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17382_ _17391_/A vssd1 vssd1 vccd1 vccd1 _17732_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14594_ _14594_/A vssd1 vssd1 vccd1 vccd1 _18769_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19121_ _19377_/CLK _19121_/D vssd1 vssd1 vccd1 vccd1 _19121_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_2_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16333_ _19428_/Q _19427_/Q _19426_/Q _16333_/D vssd1 vssd1 vccd1 vccd1 _16342_/D
+ sky130_fd_sc_hd__and4_1
XANTENNA__12080__A1 _12066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13545_ _18362_/Q _13544_/X _13545_/S vssd1 vssd1 vccd1 vccd1 _13546_/A sky130_fd_sc_hd__mux2_1
X_10757_ _19275_/Q _19113_/Q _18522_/Q _18292_/Q _10654_/A _10655_/A vssd1 vssd1 vccd1
+ vccd1 _10758_/B sky130_fd_sc_hd__mux4_1
XFILLER_158_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14308__S _14310_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_155_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19052_ _19054_/CLK _19052_/D vssd1 vssd1 vccd1 vccd1 _19052_/Q sky130_fd_sc_hd__dfxtp_1
X_16264_ _16266_/A _16264_/B vssd1 vssd1 vccd1 vccd1 _16265_/A sky130_fd_sc_hd__or2_1
X_13476_ _13476_/A vssd1 vssd1 vccd1 vccd1 _18337_/D sky130_fd_sc_hd__clkbuf_1
X_10688_ _18923_/Q _18689_/Q _19371_/Q _19019_/Q _10566_/X _10586_/X vssd1 vssd1 vccd1
+ vccd1 _10689_/B sky130_fd_sc_hd__mux4_1
XANTENNA__09459__S0 _09980_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18003_ _19774_/Q _19395_/Q _18005_/S vssd1 vssd1 vccd1 vccd1 _18004_/A sky130_fd_sc_hd__mux2_1
X_15215_ _19026_/Q _15057_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15216_/A sky130_fd_sc_hd__mux2_1
X_12427_ _17907_/B vssd1 vssd1 vccd1 vccd1 _12427_/Y sky130_fd_sc_hd__inv_2
XFILLER_173_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15928__A _15996_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16195_ _16195_/A vssd1 vssd1 vccd1 vccd1 _19370_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17846__A1 _17910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15146_ _15146_/A vssd1 vssd1 vccd1 vccd1 _18995_/D sky130_fd_sc_hd__clkbuf_1
X_12358_ _12358_/A vssd1 vssd1 vccd1 vccd1 _17885_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__09926__A _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15139__S _15145_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11309_ _11309_/A _11309_/B vssd1 vssd1 vccd1 vccd1 _11309_/X sky130_fd_sc_hd__or2_1
X_15077_ _18968_/Q _15076_/X _15077_/S vssd1 vssd1 vccd1 vccd1 _15078_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11018__S0 _11149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12289_ _12289_/A vssd1 vssd1 vccd1 vccd1 _17845_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__14043__S _14043_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ _14028_/A vssd1 vssd1 vccd1 vccd1 _18537_/D sky130_fd_sc_hd__clkbuf_1
X_18905_ _19197_/CLK _18905_/D vssd1 vssd1 vccd1 vccd1 _18905_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15609__A0 _19733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18836_ _19286_/CLK _18836_/D vssd1 vssd1 vccd1 vccd1 _18836_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10241__S1 _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11894__A1 _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18767_ _19319_/CLK _18767_/D vssd1 vssd1 vccd1 vccd1 _18767_/Q sky130_fd_sc_hd__dfxtp_1
X_15979_ _13589_/X _19321_/Q _15981_/S vssd1 vssd1 vccd1 vccd1 _15980_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18023__A1 _11969_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17718_ _17434_/X _17717_/X _17473_/X vssd1 vssd1 vccd1 vccd1 _17718_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_36_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18698_ _19124_/CLK _18698_/D vssd1 vssd1 vccd1 vccd1 _18698_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17649_ _17646_/X _17648_/X _17386_/A vssd1 vssd1 vccd1 vccd1 _17649_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11415__B _11420_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19319_ _19319_/CLK _19319_/D vssd1 vssd1 vccd1 vccd1 _19319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17102__B _17102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14348__A0 _13909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16941__B _17010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09836__A _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__S0 _10940_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09905_ _09905_/A vssd1 vssd1 vccd1 vccd1 _09905_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_101_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13792__S _13798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11885__A1 _16963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09836_ _19735_/Q vssd1 vssd1 vccd1 vccd1 _09836_/Y sky130_fd_sc_hd__inv_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15615__A3 _09234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09767_ _09767_/A vssd1 vssd1 vccd1 vccd1 _09767_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_132_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18014__A1 _11879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _10451_/S vssd1 vssd1 vccd1 vccd1 _10450_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_159_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11660_ _19631_/Q _13430_/A vssd1 vssd1 vccd1 vccd1 _11708_/A sky130_fd_sc_hd__and2_1
XFILLER_14_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _19182_/Q _18796_/Q _19246_/Q _18365_/Q _10546_/S _09419_/A vssd1 vssd1 vccd1
+ vccd1 _10612_/B sky130_fd_sc_hd__mux4_1
XFILLER_23_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11591_ _17184_/C _11591_/B _11591_/C _11591_/D vssd1 vssd1 vccd1 vccd1 _11591_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__14128__S _14136_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__A _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ _14611_/A vssd1 vssd1 vccd1 vccd1 _13330_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_168_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10542_ _10542_/A vssd1 vssd1 vccd1 vccd1 _10763_/S sky130_fd_sc_hd__buf_4
XFILLER_155_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13261_ _13261_/A vssd1 vssd1 vccd1 vccd1 _13261_/X sky130_fd_sc_hd__clkbuf_2
X_10473_ _10531_/A _10472_/X _10297_/A vssd1 vssd1 vccd1 vccd1 _10473_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15000_ _15099_/S vssd1 vssd1 vccd1 vccd1 _15013_/S sky130_fd_sc_hd__buf_4
X_12212_ _12162_/A _12164_/B _17810_/A _12305_/A vssd1 vssd1 vccd1 vccd1 _12214_/B
+ sky130_fd_sc_hd__o31a_1
X_13192_ _13275_/A vssd1 vssd1 vccd1 vccd1 _13252_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__17828__B2 _12225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input68_A io_irq_spi_irq vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10376__B2 _19725_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_123_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12143_ _19790_/Q _11351_/A _12143_/S vssd1 vssd1 vccd1 vccd1 _17222_/A sky130_fd_sc_hd__mux2_2
XFILLER_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13314__A1 input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16951_ _16951_/A _16957_/B vssd1 vssd1 vccd1 vccd1 _16951_/X sky130_fd_sc_hd__or2_1
XFILLER_150_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12074_ _12074_/A vssd1 vssd1 vccd1 vccd1 _13418_/A sky130_fd_sc_hd__buf_4
XFILLER_96_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15902_ _15902_/A vssd1 vssd1 vccd1 vccd1 _19286_/D sky130_fd_sc_hd__clkbuf_1
X_11025_ _18454_/Q _19045_/Q _19207_/Q _18422_/Q _10969_/X _11266_/A vssd1 vssd1 vccd1
+ vccd1 _11026_/B sky130_fd_sc_hd__mux4_1
X_19670_ _19695_/CLK _19670_/D vssd1 vssd1 vccd1 vccd1 _19670_/Q sky130_fd_sc_hd__dfxtp_1
X_16882_ _16882_/A vssd1 vssd1 vccd1 vccd1 _16887_/C sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_3_6_0_clock_A clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16298__B _16298_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__A _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__A3 _11338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18621_ _19098_/CLK _18621_/D vssd1 vssd1 vccd1 vccd1 _18621_/Q sky130_fd_sc_hd__dfxtp_1
X_15833_ _13586_/X _19256_/Q _15837_/S vssd1 vssd1 vccd1 vccd1 _15834_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18005__A1 _19396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18552_ _19305_/CLK _18552_/D vssd1 vssd1 vccd1 vccd1 _18552_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15764_ _15764_/A vssd1 vssd1 vccd1 vccd1 _19225_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09916__S1 _09888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12976_ _12976_/A _12976_/B vssd1 vssd1 vccd1 vccd1 _12977_/A sky130_fd_sc_hd__or2_2
XFILLER_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17524_/S _17609_/B _17502_/X _17337_/Y vssd1 vssd1 vccd1 vccd1 _17503_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_45_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _18096_/A _14860_/B _14715_/C _14860_/D vssd1 vssd1 vccd1 vccd1 _14772_/A
+ sky130_fd_sc_hd__nand4_4
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _19736_/CLK _18483_/D vssd1 vssd1 vccd1 vccd1 _18483_/Q sky130_fd_sc_hd__dfxtp_1
X_11927_ _11927_/A vssd1 vssd1 vccd1 vccd1 _11929_/A sky130_fd_sc_hd__inv_2
XFILLER_61_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15695_ _15695_/A vssd1 vssd1 vccd1 vccd1 _15704_/S sky130_fd_sc_hd__buf_6
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15422__S _15422_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17203__A _17203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17434_ _17571_/A vssd1 vssd1 vccd1 vccd1 _17434_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_162_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14646_ _14519_/X _18784_/Q _14654_/S vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11858_ _11857_/Y _11855_/A _11858_/S vssd1 vssd1 vccd1 vccd1 _11858_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17365_ _17375_/S _17365_/B vssd1 vssd1 vccd1 vccd1 _17365_/X sky130_fd_sc_hd__and2b_1
X_10809_ _10953_/A _10809_/B vssd1 vssd1 vccd1 vccd1 _10809_/X sky130_fd_sc_hd__or2_1
X_14577_ _14576_/X _18764_/Q _14583_/S vssd1 vssd1 vccd1 vccd1 _14578_/A sky130_fd_sc_hd__mux2_1
X_11789_ _11729_/A _11762_/A _11762_/B vssd1 vssd1 vccd1 vccd1 _11790_/B sky130_fd_sc_hd__a21boi_1
XFILLER_159_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19104_ _19268_/CLK _19104_/D vssd1 vssd1 vccd1 vccd1 _19104_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16316_ _19479_/Q _19478_/Q _19480_/Q _16478_/A vssd1 vssd1 vccd1 vccd1 _16486_/A
+ sky130_fd_sc_hd__and4_1
X_13528_ _15012_/A vssd1 vssd1 vccd1 vccd1 _13528_/X sky130_fd_sc_hd__clkbuf_2
X_17296_ _17291_/X _17294_/X _17509_/S vssd1 vssd1 vccd1 vccd1 _17296_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12066__B _12066_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19035_ _19035_/CLK _19035_/D vssd1 vssd1 vccd1 vccd1 _19035_/Q sky130_fd_sc_hd__dfxtp_1
X_16247_ _16255_/A _16247_/B vssd1 vssd1 vccd1 vccd1 _16248_/A sky130_fd_sc_hd__or2_1
XFILLER_127_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13459_ _12999_/X _18330_/Q _13459_/S vssd1 vssd1 vccd1 vccd1 _13460_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput104 _17122_/A vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[1] sky130_fd_sc_hd__buf_2
X_16178_ _13525_/X _19363_/Q _16180_/S vssd1 vssd1 vccd1 vccd1 _16179_/A sky130_fd_sc_hd__mux2_1
Xoutput115 _12462_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[15] sky130_fd_sc_hd__buf_2
XFILLER_115_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput126 _12474_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[25] sky130_fd_sc_hd__buf_2
XFILLER_99_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput137 _12449_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[6] sky130_fd_sc_hd__buf_2
Xoutput148 _16276_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[15] sky130_fd_sc_hd__buf_2
XFILLER_141_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _15129_/A vssd1 vssd1 vccd1 vccd1 _18987_/D sky130_fd_sc_hd__clkbuf_1
Xoutput159 _16298_/B vssd1 vssd1 vccd1 vccd1 io_ibus_addr[25] sky130_fd_sc_hd__buf_2
XFILLER_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16489__A _16546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18244__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18244__B2 _18144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15058__A1 _15057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09391__A _18780_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09621_ _10719_/A vssd1 vssd1 vccd1 vccd1 _11335_/A sky130_fd_sc_hd__clkbuf_4
X_18819_ _19237_/CLK _18819_/D vssd1 vssd1 vccd1 vccd1 _18819_/Q sky130_fd_sc_hd__dfxtp_1
X_19799_ _19799_/CLK _19799_/D vssd1 vssd1 vccd1 vccd1 _19799_/Q sky130_fd_sc_hd__dfxtp_1
X_09552_ _09552_/A vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__buf_2
XFILLER_71_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11095__A2 _12448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _10073_/A vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13241__A0 _13240_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09996__B1 _09995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17259__S _17504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16730__A1 _16731_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__A _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09843__S0 _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_103_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18235__A1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18235__B2 _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11858__A1 _11855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14411__S _14417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12720__A _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09819_ _19326_/Q _18738_/Q _18775_/Q _18349_/Q _11385_/S _09785_/A vssd1 vssd1 vccd1
+ vccd1 _09819_/X sky130_fd_sc_hd__mux4_1
XANTENNA__17994__A0 _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13027__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12830_ _12830_/A vssd1 vssd1 vccd1 vccd1 _18284_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10240__A _10509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _18270_/Q _12759_/X _11351_/A _12755_/X vssd1 vssd1 vccd1 vccd1 _18270_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12866__S _12887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _13918_/X _18734_/Q _14500_/S vssd1 vssd1 vccd1 vccd1 _14501_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13551__A _15035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17023__A _17023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11712_ _19395_/Q _11640_/X _11692_/X _11711_/X vssd1 vssd1 vccd1 vccd1 _16249_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _18071_/S vssd1 vssd1 vccd1 vccd1 _18121_/A sky130_fd_sc_hd__clkbuf_2
X_15480_ _15494_/A _18255_/Q vssd1 vssd1 vccd1 vccd1 _15480_/Y sky130_fd_sc_hd__nand2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10833__A2 _10821_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11858_/S vssd1 vssd1 vccd1 vccd1 _12392_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14431_ _13921_/X _18703_/Q _14439_/S vssd1 vssd1 vccd1 vccd1 _14432_/A sky130_fd_sc_hd__mux2_1
XFILLER_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17150_ _09096_/Y _17149_/X _17140_/X _19702_/Q vssd1 vssd1 vccd1 vccd1 _17151_/B
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_opt_1_0_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_1_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_156_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14362_ _14362_/A vssd1 vssd1 vccd1 vccd1 _18673_/D sky130_fd_sc_hd__clkbuf_1
X_11574_ _11574_/A _11574_/B vssd1 vssd1 vccd1 vccd1 _17183_/C sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_28_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_13_0_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 io_dbus_rdata[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
XFILLER_168_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16101_ _16100_/X _19347_/Q _16112_/S vssd1 vssd1 vccd1 vccd1 _16102_/A sky130_fd_sc_hd__mux2_1
Xinput28 io_dbus_rdata[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__13697__S _13703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput39 io_ibus_inst[14] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10525_ _18400_/Q _18661_/Q _18560_/Q _18895_/Q _10433_/S _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10526_/B sky130_fd_sc_hd__mux4_1
X_13313_ _13313_/A vssd1 vssd1 vccd1 vccd1 _18310_/D sky130_fd_sc_hd__clkbuf_1
X_17081_ _19687_/Q _12689_/X _17083_/S vssd1 vssd1 vccd1 vccd1 _17082_/A sky130_fd_sc_hd__mux2_1
X_14293_ _18229_/A vssd1 vssd1 vccd1 vccd1 _14293_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16032_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16053_/S sky130_fd_sc_hd__clkbuf_2
XANTENNA__09476__A _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13244_ _19763_/Q vssd1 vssd1 vccd1 vccd1 _13245_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10456_ _18401_/Q _18662_/Q _18561_/Q _18896_/Q _10500_/S _09672_/A vssd1 vssd1 vccd1
+ vccd1 _10457_/B sky130_fd_sc_hd__mux4_1
XFILLER_124_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_108_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12614__B _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13175_ _16107_/A _13176_/B vssd1 vssd1 vccd1 vccd1 _13177_/B sky130_fd_sc_hd__nor2_1
XFILLER_151_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10387_ _10390_/A _10384_/X _10386_/X vssd1 vssd1 vccd1 vccd1 _10387_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12126_ _12126_/A _12151_/C vssd1 vssd1 vccd1 vccd1 _12127_/D sky130_fd_sc_hd__nand2_1
XFILLER_151_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17983_ _17983_/A vssd1 vssd1 vccd1 vccd1 _19764_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18226__A1 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19722_ _19725_/CLK _19722_/D vssd1 vssd1 vccd1 vccd1 _19722_/Q sky130_fd_sc_hd__dfxtp_2
X_16934_ _19629_/Q _16931_/X _16932_/X _16933_/X vssd1 vssd1 vccd1 vccd1 _19629_/D
+ sky130_fd_sc_hd__o211a_1
X_12057_ _12005_/A _12030_/A _12032_/B vssd1 vssd1 vccd1 vccd1 _12057_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_77_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12630__A _16890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18226__B2 _18132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11008_ _11064_/A _11006_/X _11007_/X vssd1 vssd1 vccd1 vccd1 _11008_/X sky130_fd_sc_hd__o21a_1
XFILLER_42_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19653_ _19693_/CLK _19653_/D vssd1 vssd1 vccd1 vccd1 _19653_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16865_ _16865_/A vssd1 vssd1 vccd1 vccd1 _16871_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18604_ _19390_/CLK _18604_/D vssd1 vssd1 vccd1 vccd1 _18604_/Q sky130_fd_sc_hd__dfxtp_1
X_15816_ _15816_/A vssd1 vssd1 vccd1 vccd1 _19248_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19584_ _19845_/CLK _19584_/D vssd1 vssd1 vccd1 vccd1 _19584_/Q sky130_fd_sc_hd__dfxtp_2
X_16796_ _16800_/B _16800_/C _16795_/Y vssd1 vssd1 vccd1 vccd1 _19572_/D sky130_fd_sc_hd__o21a_1
XFILLER_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18535_ _18902_/CLK _18535_/D vssd1 vssd1 vccd1 vccd1 _18535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _15747_/A vssd1 vssd1 vccd1 vccd1 _19217_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ _19672_/Q _17028_/A _12958_/X _19336_/Q vssd1 vssd1 vccd1 vccd1 _12959_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18029__A _18029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15152__S _15156_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13461__A _13507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18466_ _19284_/CLK _18466_/D vssd1 vssd1 vccd1 vccd1 _18466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15678_ _14576_/X _19187_/Q _15682_/S vssd1 vssd1 vccd1 vccd1 _15679_/A sky130_fd_sc_hd__mux2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13223__A0 _19729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17417_ _17920_/B vssd1 vssd1 vccd1 vccd1 _17468_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14629_ _14635_/A _18207_/B vssd1 vssd1 vccd1 vccd1 _14630_/A sky130_fd_sc_hd__and2_1
X_18397_ _18894_/CLK _18397_/D vssd1 vssd1 vccd1 vccd1 _18397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16772__A _19565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _17396_/A vssd1 vssd1 vccd1 vccd1 _17497_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_158_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10588__A1 _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17279_ _17273_/X _17277_/X _17407_/A vssd1 vssd1 vccd1 vccd1 _17279_/X sky130_fd_sc_hd__mux2_1
XANTENNA__14292__A _16301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10683__S1 _10577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13526__A1 _13525_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09386__A _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19018_ _19085_/CLK _19018_/D vssd1 vssd1 vccd1 vccd1 _19018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_114_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10760__A1 _09434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18211__B _18211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14231__S _14231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09604_ _09434_/A _09593_/X _09595_/X _09603_/X _09374_/A vssd1 vssd1 vccd1 vccd1
+ _09604_/X sky130_fd_sc_hd__a221o_2
XFILLER_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10060__A _10060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09535_ _10590_/A vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__buf_2
XFILLER_37_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09466_ _09614_/A vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_25_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10371__S0 _09700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09397_ _10824_/S vssd1 vssd1 vccd1 vccd1 _11299_/S sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_174_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19113_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10028__B1 _09833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14406__S _14406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _10310_/A vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__buf_2
XANTENNA__13517__A1 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11290_ _11096_/Y _11287_/X _11467_/A _11467_/B vssd1 vssd1 vccd1 vccd1 _11463_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_164_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_189_clock clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 _19370_/CLK sky130_fd_sc_hd__clkbuf_16
X_10241_ _18405_/Q _18666_/Q _18565_/Q _18900_/Q _10450_/S _10238_/A vssd1 vssd1 vccd1
+ vccd1 _10242_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10426__S1 _10270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10172_ _09890_/A _10171_/X _09823_/A vssd1 vssd1 vccd1 vccd1 _10172_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_160_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15237__S _15239_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19807_/CLK sky130_fd_sc_hd__clkbuf_16
X_14980_ _18936_/Q vssd1 vssd1 vccd1 vccd1 _14981_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13931_ _14611_/A vssd1 vssd1 vccd1 vccd1 _13931_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_75_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11066__A _11128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16650_ _19525_/Q _16650_/B _16650_/C _16656_/C vssd1 vssd1 vccd1 vccd1 _16663_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13862_ _13861_/X _18487_/Q _13871_/S vssd1 vssd1 vccd1 vccd1 _13863_/A sky130_fd_sc_hd__mux2_1
XFILLER_75_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15601_ _15601_/A vssd1 vssd1 vccd1 vccd1 _15626_/S sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_127_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19357_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15480__B _18255_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ _12801_/X _18283_/Q _12887_/S vssd1 vssd1 vccd1 vccd1 _12814_/A sky130_fd_sc_hd__mux2_1
X_16581_ _19508_/Q _16584_/C _16546_/X vssd1 vssd1 vccd1 vccd1 _16581_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13793_ _13793_/A vssd1 vssd1 vccd1 vccd1 _18460_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18320_ _19645_/CLK _18320_/D vssd1 vssd1 vccd1 vccd1 _18320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15532_ _15531_/X _19150_/Q _15544_/S vssd1 vssd1 vccd1 vccd1 _15533_/A sky130_fd_sc_hd__mux2_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12744_/A vssd1 vssd1 vccd1 vccd1 _12744_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10362__S0 _10247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _19799_/CLK _18251_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_2
X_15463_ _15463_/A _15463_/B vssd1 vssd1 vccd1 vccd1 _15603_/A sky130_fd_sc_hd__or2_4
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16942__A1 _13404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12675_ _19584_/Q input70/X vssd1 vssd1 vccd1 vccd1 _12675_/X sky130_fd_sc_hd__or2_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17202_ _17202_/A vssd1 vssd1 vccd1 vccd1 _17802_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__15700__S _15704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12559__A2 _12507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14414_ _14414_/A vssd1 vssd1 vccd1 vccd1 _18695_/D sky130_fd_sc_hd__clkbuf_1
X_18182_ input65/X _18178_/X _18168_/X _18174_/X _19844_/Q vssd1 vssd1 vccd1 vccd1
+ _18183_/B sky130_fd_sc_hd__a32o_1
XFILLER_129_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11626_ _11723_/S vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__clkbuf_2
X_15394_ _19105_/Q _15003_/X _15400_/S vssd1 vssd1 vccd1 vccd1 _15395_/A sky130_fd_sc_hd__mux2_1
X_17133_ _17133_/A _17133_/B vssd1 vssd1 vccd1 vccd1 _17140_/A sky130_fd_sc_hd__nor2_2
XFILLER_128_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14345_ _14356_/A vssd1 vssd1 vccd1 vccd1 _14354_/S sky130_fd_sc_hd__clkbuf_4
X_11557_ _17175_/A _17917_/A _11557_/C _11557_/D vssd1 vssd1 vccd1 vccd1 _11562_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_156_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12625__A _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_156_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17064_ _19679_/Q _15550_/X _17072_/S vssd1 vssd1 vccd1 vccd1 _17065_/A sky130_fd_sc_hd__mux2_1
X_10508_ _19185_/Q _18799_/Q _19249_/Q _18368_/Q _10496_/X _09710_/A vssd1 vssd1 vccd1
+ vccd1 _10509_/B sky130_fd_sc_hd__mux4_1
X_14276_ _18040_/A vssd1 vssd1 vccd1 vccd1 _18229_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_output99_A _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11488_ _11485_/X _11492_/C _11492_/D _11487_/X vssd1 vssd1 vccd1 vccd1 _11489_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_143_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16015_ _16014_/X _19332_/Q _16025_/S vssd1 vssd1 vccd1 vccd1 _16016_/A sky130_fd_sc_hd__mux2_1
X_10439_ _10439_/A _10439_/B vssd1 vssd1 vccd1 vccd1 _10439_/Y sky130_fd_sc_hd__nor2_1
X_13227_ _15070_/A vssd1 vssd1 vccd1 vccd1 _14592_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12731__A2 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ _19157_/Q _12526_/X _12958_/X _19347_/Q _13157_/X vssd1 vssd1 vccd1 vccd1
+ _13158_/X sky130_fd_sc_hd__a221o_1
XFILLER_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11090__S1 _11100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12020_/X _12466_/B _12108_/Y vssd1 vssd1 vccd1 vccd1 _17779_/A sky130_fd_sc_hd__a21oi_4
X_13089_ _15044_/A vssd1 vssd1 vccd1 vccd1 _14566_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17670__A2 _17328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17966_ _16091_/B _19789_/Q _17968_/S vssd1 vssd1 vccd1 vccd1 _17967_/A sky130_fd_sc_hd__mux2_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16917_ _16520_/B _16915_/B _16344_/A vssd1 vssd1 vccd1 vccd1 _16917_/Y sky130_fd_sc_hd__a21oi_1
X_19705_ _19706_/CLK _19705_/D vssd1 vssd1 vccd1 vccd1 _19705_/Q sky130_fd_sc_hd__dfxtp_1
X_17897_ _17899_/A _17899_/B vssd1 vssd1 vccd1 vccd1 _17897_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09360__A1 _11512_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19636_ _19669_/CLK _19636_/D vssd1 vssd1 vccd1 vccd1 _19636_/Q sky130_fd_sc_hd__dfxtp_1
X_16848_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16883_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_93_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19567_ _19667_/CLK _19567_/D vssd1 vssd1 vccd1 vccd1 _19567_/Q sky130_fd_sc_hd__dfxtp_2
X_16779_ _19567_/Q _19566_/Q vssd1 vssd1 vccd1 vccd1 _16780_/D sky130_fd_sc_hd__and2_1
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14287__A _14290_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _16245_/A _18071_/S vssd1 vssd1 vccd1 vccd1 _12720_/A sky130_fd_sc_hd__nor2_4
XFILLER_80_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18518_ _19365_/CLK _18518_/D vssd1 vssd1 vccd1 vccd1 _18518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19498_ _19540_/CLK _19498_/D vssd1 vssd1 vccd1 vccd1 _19498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09663__A2 _12479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19543_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09251_ _16622_/A _12605_/A vssd1 vssd1 vccd1 vccd1 _12660_/B sky130_fd_sc_hd__nor2_2
X_18449_ _19202_/CLK _18449_/D vssd1 vssd1 vccd1 vccd1 _18449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _09113_/A _09182_/B _09182_/C vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__nand3b_1
XFILLER_119_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10656__S1 _10655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_174_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14750__A _14772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09844__A _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_115_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11081__S1 _11266_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13366__A _15095_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11289__A2 _12450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14896__S _14904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19376_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_84_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12238__A1 _11618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09518_ _11318_/S vssd1 vssd1 vccd1 vccd1 _09519_/A sky130_fd_sc_hd__clkbuf_8
Xclkbuf_leaf_59_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19287_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10790_ _18394_/Q _18655_/Q _18554_/Q _18889_/Q _10692_/S _09628_/X vssd1 vssd1 vccd1
+ vccd1 _10791_/B sky130_fd_sc_hd__mux4_1
XFILLER_71_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10344__S0 _10215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09989_/A vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__clkbuf_4
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12460_/A _12461_/B vssd1 vssd1 vccd1 vccd1 _12460_/Y sky130_fd_sc_hd__nor2_1
XFILLER_166_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11411_ _12422_/A _12482_/C vssd1 vssd1 vccd1 vccd1 _11492_/C sky130_fd_sc_hd__nand2_1
X_12391_ _12391_/A _12410_/C vssd1 vssd1 vccd1 vccd1 _12391_/X sky130_fd_sc_hd__xor2_1
XANTENNA__14136__S _14136_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14130_ _18578_/Q _13953_/X _14136_/S vssd1 vssd1 vccd1 vccd1 _14131_/A sky130_fd_sc_hd__mux2_1
X_11342_ _11342_/A _12460_/A vssd1 vssd1 vccd1 vccd1 _11342_/Y sky130_fd_sc_hd__nand2_1
XFILLER_152_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16152__A2 _15620_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15756__A _15767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14061_ _13851_/X _18548_/Q _14063_/S vssd1 vssd1 vccd1 vccd1 _14062_/A sky130_fd_sc_hd__mux2_1
X_11273_ _19170_/Q _18784_/Q _19234_/Q _18353_/Q _11112_/X _10910_/A vssd1 vssd1 vccd1
+ vccd1 _11274_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18132__A _18132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ _13012_/A vssd1 vssd1 vccd1 vccd1 _13012_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input50_A io_ibus_inst[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _09909_/A _10214_/Y _10219_/X _10223_/Y _09813_/A vssd1 vssd1 vccd1 vccd1
+ _10224_/X sky130_fd_sc_hd__o311a_2
XANTENNA__09754__A _09754_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11921__A0 _19855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17820_ _17917_/A _17820_/B vssd1 vssd1 vccd1 vccd1 _17820_/X sky130_fd_sc_hd__or2_1
XFILLER_95_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10155_ _09730_/A _10148_/X _10150_/X _10154_/X _09754_/X vssd1 vssd1 vccd1 vccd1
+ _10155_/X sky130_fd_sc_hd__a311o_1
XFILLER_48_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_95_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16860__B1 _16812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17751_ _10539_/Y _17652_/X _17750_/X vssd1 vssd1 vccd1 vccd1 _19722_/D sky130_fd_sc_hd__a21oi_1
XFILLER_88_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14963_ _14963_/A vssd1 vssd1 vccd1 vccd1 _18927_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_48_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_10086_ _10086_/A _09926_/Y vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__or2b_1
XFILLER_75_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16702_ _16806_/A vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__buf_4
X_13914_ _13914_/A vssd1 vssd1 vccd1 vccd1 _18503_/D sky130_fd_sc_hd__clkbuf_1
X_17682_ _17679_/X _17681_/Y _17646_/A vssd1 vssd1 vccd1 vccd1 _17682_/Y sky130_fd_sc_hd__a21oi_1
X_14894_ _14894_/A vssd1 vssd1 vccd1 vccd1 _18894_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19421_ _19421_/CLK _19421_/D vssd1 vssd1 vccd1 vccd1 _19421_/Q sky130_fd_sc_hd__dfxtp_1
X_16633_ _16660_/A _16633_/B _16633_/C vssd1 vssd1 vccd1 vccd1 _19521_/D sky130_fd_sc_hd__nor3_1
XFILLER_63_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13845_ _14525_/A vssd1 vssd1 vccd1 vccd1 _13845_/X sky130_fd_sc_hd__buf_2
XFILLER_35_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19352_ _19357_/CLK _19352_/D vssd1 vssd1 vccd1 vccd1 _19352_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16564_ hold1/A _16567_/C _16546_/X vssd1 vssd1 vccd1 vccd1 _16564_/Y sky130_fd_sc_hd__a21oi_1
X_13776_ _12886_/X _18453_/Q _13776_/S vssd1 vssd1 vccd1 vccd1 _13777_/A sky130_fd_sc_hd__mux2_1
X_10988_ _10895_/X _12450_/B _10987_/Y vssd1 vssd1 vccd1 vccd1 _11463_/A sky130_fd_sc_hd__o21bai_1
X_18303_ _19027_/CLK _18303_/D vssd1 vssd1 vccd1 vccd1 _18303_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12339__B _19419_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15515_ _15478_/X _15513_/X _15514_/Y _15508_/X hold18/X vssd1 vssd1 vccd1 vccd1
+ _15515_/X sky130_fd_sc_hd__a32o_4
X_19283_ _19377_/CLK _19283_/D vssd1 vssd1 vccd1 vccd1 _19283_/Q sky130_fd_sc_hd__dfxtp_1
X_12727_ _17795_/A vssd1 vssd1 vccd1 vccd1 _12727_/X sky130_fd_sc_hd__buf_4
X_16495_ _16541_/A _16495_/B _16495_/C vssd1 vssd1 vccd1 vccd1 _19482_/D sky130_fd_sc_hd__nor3_1
XFILLER_148_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10886__S1 _10817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18234_ _18234_/A vssd1 vssd1 vccd1 vccd1 _18234_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17211__A _17211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09929__A _10197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15446_ _15446_/A vssd1 vssd1 vccd1 vccd1 _15455_/S sky130_fd_sc_hd__buf_4
X_12658_ _19564_/Q vssd1 vssd1 vccd1 vccd1 _16778_/C sky130_fd_sc_hd__clkbuf_2
X_18165_ input61/X _18155_/X _18066_/S _12657_/X _18081_/A vssd1 vssd1 vccd1 vccd1
+ _18166_/B sky130_fd_sc_hd__a32o_1
X_11609_ _19771_/Q _11260_/X _11678_/A vssd1 vssd1 vccd1 vccd1 _12487_/B sky130_fd_sc_hd__mux2_8
XANTENNA__10638__S1 _09651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14046__S _14049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15377_ _19098_/Q _15083_/X _15383_/S vssd1 vssd1 vccd1 vccd1 _15378_/A sky130_fd_sc_hd__mux2_1
X_12589_ _12589_/A _12589_/B vssd1 vssd1 vccd1 vccd1 _12590_/B sky130_fd_sc_hd__or2_2
XFILLER_156_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17116_ _17917_/A vssd1 vssd1 vccd1 vccd1 _17907_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_117_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14328_ _13880_/X _18658_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14329_/A sky130_fd_sc_hd__mux2_1
X_18096_ _18096_/A _18142_/B vssd1 vssd1 vccd1 vccd1 _18096_/Y sky130_fd_sc_hd__nand2_1
X_17047_ _17047_/A vssd1 vssd1 vccd1 vccd1 _19671_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14259_ _14259_/A vssd1 vssd1 vccd1 vccd1 _18635_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14570__A _14602_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12165__A0 _19791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11063__S1 _11012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09581__A1 _09760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16300__C1 _16280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__S1 _10802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18998_ _19127_/CLK _18998_/D vssd1 vssd1 vccd1 vccd1 _18998_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11418__B _12479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17949_ _19749_/Q _19781_/Q _17957_/S vssd1 vssd1 vccd1 vccd1 _17950_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19619_ _19619_/CLK _19619_/D vssd1 vssd1 vccd1 vccd1 _19619_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13125__S _13172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17159__A1 _12482_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_110_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09303_ _19704_/Q _12975_/B _19702_/Q vssd1 vssd1 vccd1 vccd1 _09303_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_55_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _09289_/B vssd1 vssd1 vccd1 vccd1 _09234_/X sky130_fd_sc_hd__buf_4
X_09165_ _09167_/C _09175_/C vssd1 vssd1 vccd1 vccd1 _11566_/C sky130_fd_sc_hd__or2_1
XFILLER_163_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_108_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12943__A2 _12781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _09124_/A vssd1 vssd1 vccd1 vccd1 _09096_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_174_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14480__A _14502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11054__S1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12712__B _12712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09998_ _09998_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09998_/X sky130_fd_sc_hd__or2_1
XFILLER_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16842__B1 _16812_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11960_ _11960_/A vssd1 vssd1 vccd1 vccd1 _11968_/B sky130_fd_sc_hd__clkinv_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10911_ _18392_/Q _18653_/Q _18552_/Q _18887_/Q _09625_/A _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10912_/B sky130_fd_sc_hd__mux4_1
X_11891_ _11942_/A _12455_/B _11890_/X vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__a21o_1
XFILLER_151_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _13630_/A vssd1 vssd1 vccd1 vccd1 _18388_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10842_ _19178_/Q _18792_/Q _19242_/Q _18361_/Q _09626_/A _10837_/X vssd1 vssd1 vccd1
+ vccd1 _10843_/B sky130_fd_sc_hd__mux4_1
XFILLER_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10317__S0 _10367_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13561_ _18367_/Q _13560_/X _13561_/S vssd1 vssd1 vccd1 vccd1 _13562_/A sky130_fd_sc_hd__mux2_1
XFILLER_13_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10773_ _10773_/A vssd1 vssd1 vccd1 vccd1 _10779_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18127__A _18127_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15300_ _14598_/X _19064_/Q _15300_/S vssd1 vssd1 vccd1 vccd1 _15301_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15250__S _15256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12512_ _12584_/A vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__buf_2
XFILLER_40_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16280_ _18136_/A vssd1 vssd1 vccd1 vccd1 _16280_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_139_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13492_ _13251_/X _18345_/Q _13492_/S vssd1 vssd1 vccd1 vccd1 _13493_/A sky130_fd_sc_hd__mux2_1
X_15231_ _19033_/Q _15079_/X _15239_/S vssd1 vssd1 vccd1 vccd1 _15232_/A sky130_fd_sc_hd__mux2_1
X_12443_ _12447_/A _12443_/B vssd1 vssd1 vccd1 vccd1 _12443_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_126_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15162_ _15162_/A vssd1 vssd1 vccd1 vccd1 _19002_/D sky130_fd_sc_hd__clkbuf_1
X_12374_ _11794_/X _12369_/Y _12372_/X _12373_/Y vssd1 vssd1 vccd1 vccd1 _12374_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_60_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_154_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14113_ _14113_/A vssd1 vssd1 vccd1 vccd1 _18571_/D sky130_fd_sc_hd__clkbuf_1
X_11325_ _18398_/Q _18659_/Q _18558_/Q _18893_/Q _10692_/S _09628_/X vssd1 vssd1 vccd1
+ vccd1 _11326_/B sky130_fd_sc_hd__mux4_1
XFILLER_125_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15093_ _18973_/Q _15092_/X _15093_/S vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__mux2_1
XFILLER_107_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09484__A _09484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11256_ _18449_/Q _19040_/Q _19202_/Q _18417_/Q _11123_/A _11124_/A vssd1 vssd1 vccd1
+ vccd1 _11257_/B sky130_fd_sc_hd__mux4_2
X_18921_ _19369_/CLK _18921_/D vssd1 vssd1 vccd1 vccd1 _18921_/Q sky130_fd_sc_hd__dfxtp_1
X_14044_ _14044_/A vssd1 vssd1 vccd1 vccd1 _18542_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10207_ _10209_/A _10206_/X _09822_/A vssd1 vssd1 vccd1 vccd1 _10207_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11519__A _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11187_ _18452_/Q _19043_/Q _19205_/Q _18420_/Q _11127_/S _11177_/X vssd1 vssd1 vccd1
+ vccd1 _11188_/B sky130_fd_sc_hd__mux4_1
X_18852_ _19076_/CLK _18852_/D vssd1 vssd1 vccd1 vccd1 _18852_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_151_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _10138_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _10138_/X sky130_fd_sc_hd__and2_1
X_17803_ _17726_/A _17726_/B _17800_/B _17802_/X vssd1 vssd1 vccd1 vccd1 _17803_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18783_ _19724_/CLK _18783_/D vssd1 vssd1 vccd1 vccd1 _18783_/Q sky130_fd_sc_hd__dfxtp_1
X_15995_ _15995_/A vssd1 vssd1 vccd1 vccd1 _19328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_83_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15425__S _15433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17734_ _17592_/A _17729_/X _17733_/Y _17518_/X _12009_/B vssd1 vssd1 vccd1 vccd1
+ _17734_/X sky130_fd_sc_hd__a32o_2
XFILLER_76_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14946_ _18919_/Q vssd1 vssd1 vccd1 vccd1 _14947_/A sky130_fd_sc_hd__clkbuf_1
X_10069_ _10590_/A _10068_/X _09820_/A vssd1 vssd1 vccd1 vccd1 _10069_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_85_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10556__S0 _09415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17665_ _17662_/A _17662_/B _17419_/A _17664_/Y vssd1 vssd1 vccd1 vccd1 _17665_/X
+ sky130_fd_sc_hd__o211a_1
X_14877_ _14877_/A vssd1 vssd1 vccd1 vccd1 _18886_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_78_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16061__A1 _19340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16616_ _19519_/Q _16614_/B _16590_/X vssd1 vssd1 vccd1 vccd1 _16616_/Y sky130_fd_sc_hd__a21oi_1
X_19404_ _19699_/CLK _19404_/D vssd1 vssd1 vccd1 vccd1 _19404_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11254__A _11254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13828_ _13828_/A vssd1 vssd1 vccd1 vccd1 _18476_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17596_ _17596_/A vssd1 vssd1 vccd1 vccd1 _17786_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10308__S0 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16547_ _16551_/B _16551_/C _16546_/X vssd1 vssd1 vccd1 vccd1 _16547_/Y sky130_fd_sc_hd__a21oi_1
X_19335_ _19356_/CLK _19335_/D vssd1 vssd1 vccd1 vccd1 _19335_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_50_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ _13759_/A vssd1 vssd1 vccd1 vccd1 _18446_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19266_ _19298_/CLK _19266_/D vssd1 vssd1 vccd1 vccd1 _19266_/Q sky130_fd_sc_hd__dfxtp_1
X_16478_ _16478_/A vssd1 vssd1 vccd1 vccd1 _16483_/C sky130_fd_sc_hd__clkbuf_1
XANTENNA__14284__B _18218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18217_ _18217_/A vssd1 vssd1 vccd1 vccd1 _19855_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11701__B _12621_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15429_ _19121_/Q _15054_/X _15433_/S vssd1 vssd1 vccd1 vccd1 _15430_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17876__A _17878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19197_ _19197_/CLK _19197_/D vssd1 vssd1 vccd1 vccd1 _19197_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16780__A _19565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18148_ _18148_/A _18188_/A vssd1 vssd1 vccd1 vccd1 _18148_/Y sky130_fd_sc_hd__nand2_1
XFILLER_144_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10397__C1 _09830_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18079_ _19807_/Q _18079_/B _18099_/A vssd1 vssd1 vccd1 vccd1 _18079_/X sky130_fd_sc_hd__or3_1
XFILLER_171_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09921_ _19291_/Q _19129_/Q _18538_/Q _18308_/Q _09904_/X _09888_/X vssd1 vssd1 vccd1
+ vccd1 _09921_/X sky130_fd_sc_hd__mux4_1
XANTENNA__09394__A _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11036__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09852_ _10413_/S vssd1 vssd1 vccd1 vccd1 _10368_/S sky130_fd_sc_hd__buf_2
XFILLER_112_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16939__B _18071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _18509_/Q _19004_/Q _09786_/A vssd1 vssd1 vccd1 vccd1 _09784_/A sky130_fd_sc_hd__mux2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13644__A _13690_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17116__A _17917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10479__S _10479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11164__A _11164_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14063__A0 _13854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ _19858_/Q _19857_/Q _19856_/Q _19855_/Q vssd1 vssd1 vccd1 vccd1 _09347_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_136_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09148_ _11585_/C _09338_/C _09175_/C vssd1 vssd1 vccd1 vccd1 _11587_/A sky130_fd_sc_hd__or3_1
XFILLER_147_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10388__C1 _09812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11275__S1 _11220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10927__A1 _19111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__B _12470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16626__A_N _09241_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09079_ _09166_/B vssd1 vssd1 vccd1 vccd1 _09186_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11110_ _19172_/Q _18786_/Q _19236_/Q _18355_/Q _09624_/A _11020_/X vssd1 vssd1 vccd1
+ vccd1 _11111_/B sky130_fd_sc_hd__mux4_1
XFILLER_151_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ _12056_/A _12089_/X _12059_/A _12059_/B vssd1 vssd1 vccd1 vccd1 _12091_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_162_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11027__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12442__B _12442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _11232_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11041_/X sky130_fd_sc_hd__or2_1
XANTENNA__11339__A _19720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14800_ _14800_/A vssd1 vssd1 vccd1 vccd1 _18852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13554__A _15038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15780_ _13614_/X _19233_/Q _15780_/S vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ _19716_/Q _15513_/B _13247_/S vssd1 vssd1 vccd1 vccd1 _12992_/X sky130_fd_sc_hd__mux2_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16006__A_N _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ _14541_/X _18822_/Q _14737_/S vssd1 vssd1 vccd1 vccd1 _14732_/A sky130_fd_sc_hd__mux2_1
XANTENNA_input13_A io_dbus_rdata[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11943_ _11943_/A _12159_/A vssd1 vssd1 vccd1 vccd1 _11944_/A sky130_fd_sc_hd__nand2_1
XFILLER_73_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16043__A1 _19337_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17450_ _17456_/S vssd1 vssd1 vccd1 vccd1 _17576_/S sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _14662_/A vssd1 vssd1 vccd1 vccd1 _18791_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_73_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11874_ _11872_/X _11874_/B vssd1 vssd1 vccd1 vccd1 _11876_/A sky130_fd_sc_hd__and2b_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16401_ _19449_/Q _16399_/B _16400_/Y vssd1 vssd1 vccd1 vccd1 _19449_/D sky130_fd_sc_hd__o21a_1
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13613_ _13613_/A vssd1 vssd1 vccd1 vccd1 _18383_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _17370_/X _17379_/Y _17654_/A vssd1 vssd1 vccd1 vccd1 _17381_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10825_ _18489_/Q _18984_/Q _10872_/S vssd1 vssd1 vccd1 vccd1 _10825_/X sky130_fd_sc_hd__mux2_1
XFILLER_60_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14593_ _14592_/X _18769_/Q _14599_/S vssd1 vssd1 vccd1 vccd1 _14594_/A sky130_fd_sc_hd__mux2_1
XFILLER_158_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19120_ _19120_/CLK _19120_/D vssd1 vssd1 vccd1 vccd1 _19120_/Q sky130_fd_sc_hd__dfxtp_1
X_16332_ _16341_/A _16332_/B _16332_/C vssd1 vssd1 vccd1 vccd1 _19427_/D sky130_fd_sc_hd__nor3_1
XFILLER_158_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13544_ _15028_/A vssd1 vssd1 vccd1 vccd1 _13544_/X sky130_fd_sc_hd__buf_2
X_10756_ _18458_/Q _19049_/Q _19211_/Q _18426_/Q _10660_/X _09707_/A vssd1 vssd1 vccd1
+ vccd1 _10756_/X sky130_fd_sc_hd__mux4_1
XFILLER_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17543__A1 _17532_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19051_ _19245_/CLK _19051_/D vssd1 vssd1 vccd1 vccd1 _19051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16263_ _16263_/A vssd1 vssd1 vccd1 vccd1 _19401_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17696__A _17696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ _13124_/X _18337_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _13476_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10687_ _09820_/A _10680_/Y _10682_/Y _10684_/Y _10686_/Y vssd1 vssd1 vccd1 vccd1
+ _10687_/X sky130_fd_sc_hd__o32a_1
XFILLER_145_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18002_ _18002_/A vssd1 vssd1 vccd1 vccd1 _19773_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09459__S1 _09390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15214_ _15214_/A vssd1 vssd1 vccd1 vccd1 _19025_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_139_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12426_ _17920_/A _12426_/B vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__nand2_2
X_16194_ _13547_/X _19370_/Q _16202_/S vssd1 vssd1 vccd1 vccd1 _16195_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15145_ _18995_/Q _15060_/X _15145_/S vssd1 vssd1 vccd1 vccd1 _15146_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14324__S _14332_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ _19799_/Q _11416_/A _12357_/S vssd1 vssd1 vccd1 vccd1 _12358_/A sky130_fd_sc_hd__mux2_8
XANTENNA__09926__B _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output81_A _12149_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11308_ _19183_/Q _18797_/Q _19247_/Q _18366_/Q _10729_/S _10655_/X vssd1 vssd1 vccd1
+ vccd1 _11309_/B sky130_fd_sc_hd__mux4_1
X_15076_ _15076_/A vssd1 vssd1 vccd1 vccd1 _15076_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__11018__S1 _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12288_ _12288_/A _12314_/A vssd1 vssd1 vccd1 vccd1 _12312_/B sky130_fd_sc_hd__or2_2
XFILLER_84_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18904_ _19096_/CLK _18904_/D vssd1 vssd1 vccd1 vccd1 _18904_/Q sky130_fd_sc_hd__dfxtp_1
X_14027_ _18537_/Q _14026_/X _14027_/S vssd1 vssd1 vccd1 vccd1 _14028_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10153__A _10197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ _11239_/A _12443_/B vssd1 vssd1 vccd1 vccd1 _11239_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18835_ _19378_/CLK _18835_/D vssd1 vssd1 vccd1 vccd1 _18835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18766_ _19378_/CLK _18766_/D vssd1 vssd1 vccd1 vccd1 _18766_/Q sky130_fd_sc_hd__dfxtp_1
X_15978_ _15978_/A vssd1 vssd1 vccd1 vccd1 _19320_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17717_ _17715_/Y _17716_/X _17717_/S vssd1 vssd1 vccd1 vccd1 _17717_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14929_ _14929_/A vssd1 vssd1 vccd1 vccd1 _18910_/D sky130_fd_sc_hd__clkbuf_1
X_18697_ _19124_/CLK _18697_/D vssd1 vssd1 vccd1 vccd1 _18697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09235__C_N _09234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17648_ _17579_/X _17647_/X _17648_/S vssd1 vssd1 vccd1 vccd1 _17648_/X sky130_fd_sc_hd__mux2_2
XFILLER_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15793__A0 _13528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17579_ _17654_/A _17351_/Y _17399_/Y vssd1 vssd1 vccd1 vccd1 _17579_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12808__A _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19318_ _19319_/CLK _19318_/D vssd1 vssd1 vccd1 vccd1 _19318_/Q sky130_fd_sc_hd__dfxtp_1
X_19249_ _19249_/CLK _19249_/D vssd1 vssd1 vccd1 vccd1 _19249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14234__S _14242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11009__S1 _11005_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09904_ _10217_/S vssd1 vssd1 vccd1 vccd1 _09904_/X sky130_fd_sc_hd__buf_4
XFILLER_116_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10768__S0 _11297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input5_A io_dbus_rdata[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09835_ _09835_/A vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__buf_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15065__S _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09766_ _09909_/A vssd1 vssd1 vccd1 vccd1 _09767_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11637__A2 _17317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09697_ _10138_/A _09691_/X _09732_/A vssd1 vssd1 vccd1 vccd1 _09697_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16025__A1 _19334_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17773__A1 _12092_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14409__S _14417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ _09995_/X _10601_/X _10605_/X _10609_/X _09374_/A vssd1 vssd1 vccd1 vccd1
+ _10610_/X sky130_fd_sc_hd__a311o_4
XFILLER_168_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11590_ _09210_/X _09211_/A _09211_/B _17109_/A _11557_/C vssd1 vssd1 vccd1 vccd1
+ _11591_/D sky130_fd_sc_hd__a311o_1
XFILLER_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11341__B _12460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ _11347_/A _12462_/A vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__or2_1
XFILLER_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10238__A _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13260_ _13260_/A vssd1 vssd1 vccd1 vccd1 _13260_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10472_ _19282_/Q _19120_/Q _18529_/Q _18299_/Q _10260_/A _09769_/A vssd1 vssd1 vccd1
+ vccd1 _10472_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13011__B2 _19338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17289__A0 _12383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12211_ _12301_/A _12471_/B _12210_/Y vssd1 vssd1 vccd1 vccd1 _17820_/B sky130_fd_sc_hd__o21ai_4
XFILLER_170_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13191_ _14585_/A vssd1 vssd1 vccd1 vccd1 _13191_/X sky130_fd_sc_hd__buf_2
XFILLER_109_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12453__A _12453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10376__A2 _10364_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12770__B1 _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12142_ _12142_/A _12142_/B vssd1 vssd1 vccd1 vccd1 _12170_/A sky130_fd_sc_hd__xnor2_1
XFILLER_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13983__S _13995_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16950_ _19634_/Q _16943_/X _16949_/X vssd1 vssd1 vccd1 vccd1 _19634_/D sky130_fd_sc_hd__a21o_1
X_12073_ _11794_/X _12063_/Y _12067_/X _12072_/Y vssd1 vssd1 vccd1 vccd1 _12073_/Y
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__18140__A _18140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15901_ _19286_/Q _14585_/A _15909_/S vssd1 vssd1 vccd1 vccd1 _15902_/A sky130_fd_sc_hd__mux2_1
X_11024_ _11024_/A vssd1 vssd1 vccd1 vccd1 _11026_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16881_ _16881_/A _16881_/B _16881_/C vssd1 vssd1 vccd1 vccd1 _19605_/D sky130_fd_sc_hd__nor3_1
XFILLER_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_24_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ _15832_/A vssd1 vssd1 vccd1 vccd1 _19255_/D sky130_fd_sc_hd__clkbuf_1
X_18620_ _18987_/CLK _18620_/D vssd1 vssd1 vccd1 vccd1 _18620_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15763_ _13589_/X _19225_/Q _15765_/S vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__mux2_1
X_18551_ _19272_/CLK _18551_/D vssd1 vssd1 vccd1 vccd1 _18551_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12975_ _12975_/A _12975_/B _19702_/Q input30/X vssd1 vssd1 vccd1 vccd1 _12976_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17213__A0 _17743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17502_ _17511_/S _17396_/B _17500_/S vssd1 vssd1 vccd1 vccd1 _17502_/X sky130_fd_sc_hd__o21a_1
X_14714_ _14714_/A vssd1 vssd1 vccd1 vccd1 _18815_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _19361_/CLK _18482_/D vssd1 vssd1 vccd1 vccd1 _18482_/Q sky130_fd_sc_hd__dfxtp_1
X_11926_ _11928_/A _17201_/A vssd1 vssd1 vccd1 vccd1 _11927_/A sky130_fd_sc_hd__or2_1
X_15694_ _15694_/A vssd1 vssd1 vccd1 vccd1 _19194_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ _17871_/A vssd1 vssd1 vccd1 vccd1 _17571_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645_ _14713_/S vssd1 vssd1 vccd1 vccd1 _14654_/S sky130_fd_sc_hd__clkbuf_4
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11857_ _11879_/A _11879_/C vssd1 vssd1 vccd1 vccd1 _11857_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10808_ _19306_/Q _18718_/Q _18755_/Q _18329_/Q _10872_/S _10802_/X vssd1 vssd1 vccd1
+ vccd1 _10809_/B sky130_fd_sc_hd__mux4_1
X_17364_ _17364_/A vssd1 vssd1 vccd1 vccd1 _17364_/Y sky130_fd_sc_hd__clkinv_2
X_14576_ _14576_/A vssd1 vssd1 vccd1 vccd1 _14576_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11788_ _11788_/A _11788_/B _11788_/C vssd1 vssd1 vccd1 vccd1 _11790_/A sky130_fd_sc_hd__and3_1
X_16315_ _19475_/Q _19477_/Q _19476_/Q _16469_/A vssd1 vssd1 vccd1 vccd1 _16478_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10064__A1 _10289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19103_ _19297_/CLK _19103_/D vssd1 vssd1 vccd1 vccd1 _19103_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15939__A _15996_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13527_ _13527_/A vssd1 vssd1 vccd1 vccd1 _18356_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_158_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17295_ _17501_/S vssd1 vssd1 vccd1 vccd1 _17509_/S sky130_fd_sc_hd__clkbuf_2
X_10739_ _10769_/A _10739_/B vssd1 vssd1 vccd1 vccd1 _10739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_174_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_159_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19034_ _19386_/CLK _19034_/D vssd1 vssd1 vccd1 vccd1 _19034_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09937__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16246_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16255_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_173_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ _13458_/A vssd1 vssd1 vccd1 vccd1 _18329_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12409_ _12391_/A _12410_/C _19422_/Q vssd1 vssd1 vccd1 vccd1 _12409_/Y sky130_fd_sc_hd__a21oi_1
X_16177_ _16177_/A vssd1 vssd1 vccd1 vccd1 _19362_/D sky130_fd_sc_hd__clkbuf_1
X_13389_ _17028_/A _13389_/B _16937_/B _16939_/A vssd1 vssd1 vccd1 vccd1 _13391_/D
+ sky130_fd_sc_hd__or4_2
Xoutput105 _17174_/A vssd1 vssd1 vccd1 vccd1 io_dbus_ld_type[2] sky130_fd_sc_hd__buf_2
XFILLER_126_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput116 _12464_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[16] sky130_fd_sc_hd__buf_2
XANTENNA__12761__B1 _11351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput127 _12476_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[26] sky130_fd_sc_hd__buf_2
XFILLER_5_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput138 _12450_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[7] sky130_fd_sc_hd__buf_2
X_15128_ _18987_/Q _15035_/X _15134_/S vssd1 vssd1 vccd1 vccd1 _15129_/A sky130_fd_sc_hd__mux2_1
XFILLER_142_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput149 _12080_/X vssd1 vssd1 vccd1 vccd1 io_ibus_addr[16] sky130_fd_sc_hd__buf_2
XFILLER_99_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15059_ _15059_/A vssd1 vssd1 vccd1 vccd1 _18962_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09672__A _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold21_A hold21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_95_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09620_ _10839_/A vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__clkbuf_2
X_18818_ _19202_/CLK _18818_/D vssd1 vssd1 vccd1 vccd1 _18818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19798_ _19800_/CLK _19798_/D vssd1 vssd1 vccd1 vccd1 _19798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09551_ _18645_/Q vssd1 vssd1 vccd1 vccd1 _09552_/A sky130_fd_sc_hd__inv_2
X_18749_ _19202_/CLK _18749_/D vssd1 vssd1 vccd1 vccd1 _18749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17204__A0 _17680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09482_ _09482_/A vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18209__B _18209_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14229__S _14231_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16191__A0 _13544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09843__S1 _09714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09582__A _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_115_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09818_ _10129_/A vssd1 vssd1 vccd1 vccd1 _11402_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10521__A _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09749_ _19294_/Q _19132_/Q _18541_/Q _18311_/Q _09743_/A _09715_/X vssd1 vssd1 vccd1
+ vccd1 _09750_/B sky130_fd_sc_hd__mux4_1
XFILLER_27_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ _18269_/Q _12759_/X _10401_/A _12755_/X vssd1 vssd1 vccd1 vccd1 _18269_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _16162_/S _11710_/X _11623_/X vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__a21o_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _19586_/Q _12690_/X _14518_/B vssd1 vssd1 vccd1 vccd1 _12691_/X sky130_fd_sc_hd__mux2_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10833__A3 _10832_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A vssd1 vssd1 vccd1 vccd1 _14439_/S sky130_fd_sc_hd__buf_4
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ _12100_/A vssd1 vssd1 vccd1 vccd1 _11858_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12167__B _17202_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14361_ _13928_/X _18673_/Q _14365_/S vssd1 vssd1 vccd1 vccd1 _14362_/A sky130_fd_sc_hd__mux2_1
XFILLER_168_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_128_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11573_ _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11575_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18135__A _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16100_ _12233_/X _15568_/X _16099_/Y vssd1 vssd1 vccd1 vccd1 _16100_/X sky130_fd_sc_hd__a21o_1
Xinput18 io_dbus_rdata[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_2
X_13312_ _13311_/X _18310_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _13313_/A sky130_fd_sc_hd__mux2_1
X_17080_ _17080_/A vssd1 vssd1 vccd1 vccd1 _19686_/D sky130_fd_sc_hd__clkbuf_1
X_10524_ _10277_/A _10523_/X _09821_/A vssd1 vssd1 vccd1 vccd1 _10524_/Y sky130_fd_sc_hd__o21ai_1
Xinput29 io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_4
XFILLER_168_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14292_ _16301_/A vssd1 vssd1 vccd1 vccd1 _14635_/A sky130_fd_sc_hd__clkbuf_1
X_16031_ _16919_/A _16029_/Y _16052_/S vssd1 vssd1 vccd1 vccd1 _16031_/X sky130_fd_sc_hd__mux2_1
X_13243_ input17/X _13134_/X _13167_/A vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__a21o_1
XFILLER_136_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10455_ _18593_/Q _18864_/Q _19088_/Q _18832_/Q _10499_/S _10229_/A vssd1 vssd1 vccd1
+ vccd1 _10455_/X sky130_fd_sc_hd__mux4_1
XFILLER_109_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12743__B1 _10895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13174_ _19759_/Q vssd1 vssd1 vccd1 vccd1 _16107_/A sky130_fd_sc_hd__clkbuf_2
X_10386_ _10471_/A _10385_/X _09764_/A vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__o21a_1
X_12125_ _19410_/Q _12151_/C vssd1 vssd1 vccd1 vccd1 _12127_/C sky130_fd_sc_hd__or2_1
XFILLER_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14496__A0 _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17982_ _19764_/Q _19796_/Q _17990_/S vssd1 vssd1 vccd1 vccd1 _17983_/A sky130_fd_sc_hd__mux2_1
X_19721_ _19736_/CLK _19721_/D vssd1 vssd1 vccd1 vccd1 _19721_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__09492__A _09644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16933_ _16981_/A vssd1 vssd1 vccd1 vccd1 _16933_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12056_ _12056_/A _12089_/A vssd1 vssd1 vccd1 vccd1 _12059_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10506__C1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09911__A1 _10174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11007_ _11007_/A vssd1 vssd1 vccd1 vccd1 _11007_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19652_ _19693_/CLK _19652_/D vssd1 vssd1 vccd1 vccd1 _19652_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16864_ _16881_/A _16864_/B _16864_/C vssd1 vssd1 vccd1 vccd1 _19599_/D sky130_fd_sc_hd__nor3_1
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18603_ _19098_/CLK _18603_/D vssd1 vssd1 vccd1 vccd1 _18603_/Q sky130_fd_sc_hd__dfxtp_1
X_15815_ _13560_/X _19248_/Q _15815_/S vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15996__A0 _13614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16795_ _16800_/B _16800_/C _16764_/X vssd1 vssd1 vccd1 vccd1 _16795_/Y sky130_fd_sc_hd__a21oi_1
X_19583_ _19583_/CLK _19583_/D vssd1 vssd1 vccd1 vccd1 _19583_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15433__S _15433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18534_ _19287_/CLK _18534_/D vssd1 vssd1 vccd1 vccd1 _18534_/Q sky130_fd_sc_hd__dfxtp_1
X_15746_ _13563_/X _19217_/Q _15754_/S vssd1 vssd1 vccd1 vccd1 _15747_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17214__A _17214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12958_ _12958_/A vssd1 vssd1 vccd1 vccd1 _12958_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ _11908_/Y _11904_/A _12179_/B vssd1 vssd1 vccd1 vccd1 _11909_/X sky130_fd_sc_hd__mux2_1
X_15677_ _15677_/A vssd1 vssd1 vccd1 vccd1 _19186_/D sky130_fd_sc_hd__clkbuf_1
X_18465_ _19314_/CLK _18465_/D vssd1 vssd1 vccd1 vccd1 _18465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16945__C1 _16933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12358__A _12358_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ _19744_/Q vssd1 vssd1 vccd1 vccd1 _16021_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__14049__S _14049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14628_ input41/X _18148_/A _14293_/X _14623_/X _09194_/X vssd1 vssd1 vccd1 vccd1
+ _18207_/B sky130_fd_sc_hd__a32o_2
X_17416_ _17603_/A vssd1 vssd1 vccd1 vccd1 _17920_/B sky130_fd_sc_hd__buf_2
XANTENNA__14420__A0 _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13223__A1 _15586_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18396_ _19312_/CLK _18396_/D vssd1 vssd1 vccd1 vccd1 _18396_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16772__B _16778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17347_ _17294_/S _17251_/X _17346_/X vssd1 vssd1 vccd1 vccd1 _17347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12792__S _13143_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ _14559_/A vssd1 vssd1 vccd1 vccd1 _18758_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18162__A1 _09172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17278_ _17512_/S vssd1 vssd1 vccd1 vccd1 _17407_/A sky130_fd_sc_hd__clkbuf_2
X_19017_ _19113_/CLK _19017_/D vssd1 vssd1 vccd1 vccd1 _19017_/Q sky130_fd_sc_hd__dfxtp_1
X_16229_ _13599_/X _19386_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16230_/A sky130_fd_sc_hd__mux2_1
XFILLER_162_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09603_ _09597_/X _09601_/X _09602_/X vssd1 vssd1 vccd1 vccd1 _09603_/X sky130_fd_sc_hd__o21a_1
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09534_ _09632_/A vssd1 vssd1 vccd1 vccd1 _10590_/A sky130_fd_sc_hd__buf_4
XFILLER_83_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15739__A0 _13554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09465_ _09465_/A vssd1 vssd1 vccd1 vccd1 _09614_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16936__C1 _16933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16963__A _16963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10371__S1 _10229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09396_ _09396_/A vssd1 vssd1 vccd1 vccd1 _10824_/S sky130_fd_sc_hd__buf_4
XFILLER_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10028__A1 _09760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13798__S _13798_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16174__S _16180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_164_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12725__A0 _18252_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ _10509_/A vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10171_ _18934_/Q _18700_/Q _19382_/Q _19030_/Q _09782_/A _09956_/A vssd1 vssd1 vccd1
+ vccd1 _10171_/X sky130_fd_sc_hd__mux4_1
XANTENNA__14422__S _14428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14478__A0 _13886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12450__B _12450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13930_ _13930_/A vssd1 vssd1 vccd1 vccd1 _18508_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11347__A _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13861_ _14541_/A vssd1 vssd1 vccd1 vccd1 _13861_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11139__S0 _11173_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15600_ _15565_/X _15598_/X _15599_/Y _12575_/X _18276_/Q vssd1 vssd1 vccd1 vccd1
+ _15600_/X sky130_fd_sc_hd__a32o_2
X_12812_ _13387_/S vssd1 vssd1 vccd1 vccd1 _12887_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_90_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16580_ _19507_/Q _16578_/B _16579_/Y vssd1 vssd1 vccd1 vccd1 _19507_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13792_ _13038_/X _18460_/Q _13798_/S vssd1 vssd1 vccd1 vccd1 _13793_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15531_ _19719_/Q _12669_/X _15543_/S vssd1 vssd1 vccd1 vccd1 _15531_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ _18258_/Q _12739_/X _10895_/X _12740_/X vssd1 vssd1 vccd1 vccd1 _18258_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12661__C1 _12660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12178__A _19412_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10362__S1 _10238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18250_ _19838_/CLK input70/X vssd1 vssd1 vccd1 vccd1 _18250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _13391_/B _11551_/A _13391_/D _11805_/D vssd1 vssd1 vccd1 vccd1 _15463_/B
+ sky130_fd_sc_hd__o31a_1
X_12674_ _12674_/A vssd1 vssd1 vccd1 vccd1 _12674_/X sky130_fd_sc_hd__buf_2
XFILLER_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17201_ _17201_/A vssd1 vssd1 vccd1 vccd1 _17680_/B sky130_fd_sc_hd__clkinv_2
X_14413_ _13896_/X _18695_/Q _14417_/S vssd1 vssd1 vccd1 vccd1 _14414_/A sky130_fd_sc_hd__mux2_1
XFILLER_129_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18181_ _18181_/A vssd1 vssd1 vccd1 vccd1 _19843_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11625_ _12078_/A _11612_/X _11622_/X _11624_/X vssd1 vssd1 vccd1 vccd1 _16243_/B
+ sky130_fd_sc_hd__a31o_1
X_15393_ _15393_/A vssd1 vssd1 vccd1 vccd1 _19104_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_156_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12906__A _15015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17132_ _19697_/Q _17131_/Y _17142_/A vssd1 vssd1 vccd1 vccd1 _19697_/D sky130_fd_sc_hd__o21a_1
XFILLER_11_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13501__S _13503_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ _14344_/A vssd1 vssd1 vccd1 vccd1 _18665_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ _11589_/B _11556_/B vssd1 vssd1 vccd1 vccd1 _11557_/C sky130_fd_sc_hd__nor2_1
XANTENNA__10975__C1 _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17063_ _17085_/A vssd1 vssd1 vccd1 vccd1 _17072_/S sky130_fd_sc_hd__clkbuf_2
X_10507_ _09726_/A _10498_/X _10502_/X _10506_/X _09669_/A vssd1 vssd1 vccd1 vccd1
+ _10507_/X sky130_fd_sc_hd__a311o_4
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14275_ _14275_/A _14275_/B _14275_/C _11649_/B vssd1 vssd1 vccd1 vccd1 _18040_/A
+ sky130_fd_sc_hd__nor4b_2
XFILLER_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11487_ _17117_/A _09142_/A _11487_/S vssd1 vssd1 vccd1 vccd1 _11487_/X sky130_fd_sc_hd__mux2_1
XFILLER_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12716__A0 _12715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16014_ _15481_/X _16013_/Y _16024_/S vssd1 vssd1 vccd1 vccd1 _16014_/X sky130_fd_sc_hd__mux2_1
XFILLER_109_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13226_ _13214_/X _13224_/Y _13225_/Y vssd1 vssd1 vccd1 vccd1 _15070_/A sky130_fd_sc_hd__a21oi_4
X_10438_ _18929_/Q _18695_/Q _19377_/Q _19025_/Q _10341_/S _09886_/A vssd1 vssd1 vccd1
+ vccd1 _10439_/B sky130_fd_sc_hd__mux4_1
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13157_ _19683_/Q _12659_/X _12680_/X _19650_/Q vssd1 vssd1 vccd1 vccd1 _13157_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_124_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10414_/A _10368_/X _10404_/A vssd1 vssd1 vccd1 vccd1 _10369_/X sky130_fd_sc_hd__a21o_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14332__S _14332_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _18114_/A _12021_/X _12022_/X vssd1 vssd1 vccd1 vccd1 _12108_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13088_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__and2_4
X_17965_ _17965_/A vssd1 vssd1 vccd1 vccd1 _19756_/D sky130_fd_sc_hd__clkbuf_1
X_19704_ _19706_/CLK _19704_/D vssd1 vssd1 vccd1 vccd1 _19704_/Q sky130_fd_sc_hd__dfxtp_1
X_16916_ _19618_/Q _16914_/B _16915_/Y vssd1 vssd1 vccd1 vccd1 _19618_/D sky130_fd_sc_hd__o21a_1
X_12039_ _12066_/A _12066_/C vssd1 vssd1 vccd1 vccd1 _12065_/B sky130_fd_sc_hd__and2_1
X_17896_ _17899_/A _17899_/B _17896_/S vssd1 vssd1 vccd1 vccd1 _17896_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16767__B _19562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19635_ _19635_/CLK _19635_/D vssd1 vssd1 vccd1 vccd1 _19635_/Q sky130_fd_sc_hd__dfxtp_1
X_16847_ _16881_/A _16847_/B _16847_/C vssd1 vssd1 vccd1 vccd1 _19593_/D sky130_fd_sc_hd__nor3_1
XFILLER_168_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13472__A _13494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15163__S _15167_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19566_ _19663_/CLK _19566_/D vssd1 vssd1 vccd1 vccd1 _19566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16778_ _16782_/C _19565_/Q _16778_/C _16780_/C vssd1 vssd1 vccd1 vccd1 _16778_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14287__B _18220_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18517_ _19301_/CLK _18517_/D vssd1 vssd1 vccd1 vccd1 _18517_/Q sky130_fd_sc_hd__dfxtp_1
X_15729_ _15729_/A vssd1 vssd1 vccd1 vccd1 _19209_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16783__A _16840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19497_ _19619_/CLK _19497_/D vssd1 vssd1 vccd1 vccd1 _19497_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _16623_/A _16623_/B _16625_/A _09253_/C vssd1 vssd1 vccd1 vccd1 _12605_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_22_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18448_ _19071_/CLK _18448_/D vssd1 vssd1 vccd1 vccd1 _18448_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_167_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ _09207_/A _11526_/A vssd1 vssd1 vccd1 vccd1 _11541_/A sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_146_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18379_ _19386_/CLK _18379_/D vssd1 vssd1 vccd1 vccd1 _18379_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14507__S _14511_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09397__A _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10966__C1 _11160_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18222__B _18222_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12551__A _16245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14242__S _14242_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10071__A _10289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17949__A1 _19781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09860__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10041__S0 _09441_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14197__B _14197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09517_ _10056_/A vssd1 vssd1 vccd1 vccd1 _10347_/A sky130_fd_sc_hd__buf_2
XFILLER_24_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__A1 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ _09448_/A vssd1 vssd1 vccd1 vccd1 _09989_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_158_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14417__S _14417_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09379_ _09442_/A vssd1 vssd1 vccd1 vccd1 _09380_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11410_ _12422_/A _12482_/C vssd1 vssd1 vccd1 vccd1 _11412_/A sky130_fd_sc_hd__or2_1
XFILLER_149_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ _19421_/Q vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__buf_2
XFILLER_149_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_166_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12445__B _12445_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10957__C1 _09448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ _11342_/A _12460_/A vssd1 vssd1 vccd1 vccd1 _11343_/A sky130_fd_sc_hd__nor2_1
XFILLER_125_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14060_ _14060_/A vssd1 vssd1 vccd1 vccd1 _18547_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11272_ _09481_/A _11262_/Y _11267_/X _11271_/Y _09552_/A vssd1 vssd1 vccd1 vccd1
+ _11272_/X sky130_fd_sc_hd__o311a_1
X_13011_ _19148_/Q _13007_/X _12566_/X _19338_/Q _13010_/X vssd1 vssd1 vccd1 vccd1
+ _13011_/X sky130_fd_sc_hd__a221o_2
XANTENNA__15248__S _15256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10223_ _09968_/A _10220_/X _10222_/X vssd1 vssd1 vccd1 vccd1 _10223_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13557__A _15041_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17029__A _17085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14152__S _14158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12461__A _12461_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11382__C1 _09859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input43_A io_ibus_inst[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _10105_/A _10151_/X _10153_/X _09857_/X vssd1 vssd1 vccd1 vccd1 _10154_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16868__A _16868_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11077__A _11232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14962_ _18927_/Q vssd1 vssd1 vccd1 vccd1 _14963_/A sky130_fd_sc_hd__clkbuf_1
X_17750_ _12035_/A _17737_/X _17749_/X _17831_/A vssd1 vssd1 vccd1 vccd1 _17750_/X
+ sky130_fd_sc_hd__o211a_4
XFILLER_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10085_ _11424_/A _11360_/B _10084_/Y _11427_/B vssd1 vssd1 vccd1 vccd1 _11361_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16701_ _16706_/C _16706_/D _16700_/Y vssd1 vssd1 vccd1 vccd1 _19543_/D sky130_fd_sc_hd__o21a_1
XANTENNA__09770__A _10270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10488__A1 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13913_ _13912_/X _18503_/Q _13919_/S vssd1 vssd1 vccd1 vccd1 _13914_/A sky130_fd_sc_hd__mux2_1
X_14893_ _18894_/Q _13994_/X _14893_/S vssd1 vssd1 vccd1 vccd1 _14894_/A sky130_fd_sc_hd__mux2_1
X_17681_ _17910_/A _17676_/Y _17680_/Y _17597_/A vssd1 vssd1 vccd1 vccd1 _17681_/Y
+ sky130_fd_sc_hd__a211oi_1
X_19420_ _19423_/CLK _19420_/D vssd1 vssd1 vccd1 vccd1 _19420_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16632_ _16634_/B _16659_/B vssd1 vssd1 vccd1 vccd1 _16633_/C sky130_fd_sc_hd__and2_1
X_13844_ _13844_/A vssd1 vssd1 vccd1 vccd1 _18481_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19351_ _19357_/CLK _19351_/D vssd1 vssd1 vccd1 vccd1 _19351_/Q sky130_fd_sc_hd__dfxtp_2
X_16563_ _19501_/Q _16561_/B _16562_/Y vssd1 vssd1 vccd1 vccd1 _19501_/D sky130_fd_sc_hd__o21a_1
X_13775_ _13775_/A vssd1 vssd1 vccd1 vccd1 _18452_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10987_ _10895_/X _12450_/B _11288_/A _12449_/B vssd1 vssd1 vccd1 vccd1 _10987_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18302_ _19285_/CLK _18302_/D vssd1 vssd1 vccd1 vccd1 _18302_/Q sky130_fd_sc_hd__dfxtp_1
X_15514_ _15541_/A hold18/A vssd1 vssd1 vccd1 vccd1 _15514_/Y sky130_fd_sc_hd__nand2_1
X_12726_ _12726_/A vssd1 vssd1 vccd1 vccd1 _18252_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_149_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16494_ _16493_/A _16493_/C _19482_/Q vssd1 vssd1 vccd1 vccd1 _16495_/C sky130_fd_sc_hd__a21oi_1
X_19282_ _19282_/CLK _19282_/D vssd1 vssd1 vccd1 vccd1 _19282_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15445_ _15445_/A vssd1 vssd1 vccd1 vccd1 _19128_/D sky130_fd_sc_hd__clkbuf_1
X_18233_ _18233_/A vssd1 vssd1 vccd1 vccd1 _18248_/A sky130_fd_sc_hd__clkbuf_1
X_12657_ _14623_/A vssd1 vssd1 vccd1 vccd1 _12657_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_157_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ _11606_/X _11608_/B vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__and2b_1
X_18164_ _18164_/A vssd1 vssd1 vccd1 vccd1 _19839_/D sky130_fd_sc_hd__clkbuf_1
X_15376_ _15376_/A vssd1 vssd1 vccd1 vccd1 _19097_/D sky130_fd_sc_hd__clkbuf_1
X_12588_ _19606_/Q _12697_/A _12583_/X _19538_/Q _12587_/X vssd1 vssd1 vccd1 vccd1
+ _12589_/B sky130_fd_sc_hd__a221o_1
XFILLER_157_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10948__C1 _10883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14327_ _14327_/A vssd1 vssd1 vccd1 vccd1 _18657_/D sky130_fd_sc_hd__clkbuf_1
X_17115_ _17115_/A vssd1 vssd1 vccd1 vccd1 _17115_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18095_ _14860_/B _18086_/X _18094_/X _18084_/X vssd1 vssd1 vccd1 vccd1 _19813_/D
+ sky130_fd_sc_hd__o211a_1
X_11539_ _11538_/X _17166_/A _11539_/S vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_144_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_116_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17046_ _19671_/Q _16932_/A _17050_/S vssd1 vssd1 vccd1 vccd1 _17047_/A sky130_fd_sc_hd__mux2_1
XFILLER_143_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14258_ _18635_/Q _14033_/X _14264_/S vssd1 vssd1 vccd1 vccd1 _14259_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12165__A1 _10303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13209_ _14589_/A vssd1 vssd1 vccd1 vccd1 _13209_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_174_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12371__A _19420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14189_ _18605_/Q _14039_/X _14191_/S vssd1 vssd1 vccd1 vccd1 _14190_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__A2 _09555_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18997_ _19096_/CLK _18997_/D vssd1 vssd1 vccd1 vccd1 _18997_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17957_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_79_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_173_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19367_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_39_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_72_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__S0 _10022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17879_ _17490_/X _17876_/Y _17878_/Y vssd1 vssd1 vccd1 vccd1 _17879_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_65_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19618_ _19618_/CLK _19618_/D vssd1 vssd1 vccd1 vccd1 _19618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13417__B2 _18253_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19549_ _19549_/CLK _19549_/D vssd1 vssd1 vccd1 vccd1 _19549_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_188_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19308_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09302_ _19703_/Q vssd1 vssd1 vccd1 vccd1 _12975_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ _19700_/Q _19699_/Q vssd1 vssd1 vccd1 vccd1 _09289_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_111_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19845_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09164_ _09325_/A _18100_/A _09176_/A _17114_/C vssd1 vssd1 vccd1 vccd1 _09169_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_159_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12265__B _12289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09095_ _09186_/A _09186_/B _11646_/B _11513_/C vssd1 vssd1 vccd1 vccd1 _09124_/A
+ sky130_fd_sc_hd__or4_4
XANTENNA__14761__A _14772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_126_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19660_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_162_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15068__S _15077_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09997_ _18475_/Q _19066_/Q _19228_/Q _18443_/Q _09850_/A _09977_/X vssd1 vssd1 vccd1
+ vccd1 _09998_/B sky130_fd_sc_hd__mux4_1
XFILLER_131_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09590__A _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10910_ _10910_/A vssd1 vssd1 vccd1 vccd1 _10910_/X sky130_fd_sc_hd__buf_2
XFILLER_56_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11890_ _18144_/A _11890_/B _11890_/C vssd1 vssd1 vccd1 vccd1 _11890_/X sky130_fd_sc_hd__and3_1
XFILLER_151_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10841_ _10848_/A _10840_/X _09482_/A vssd1 vssd1 vccd1 vccd1 _10841_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_71_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13560_ _15044_/A vssd1 vssd1 vccd1 vccd1 _13560_/X sky130_fd_sc_hd__buf_2
X_10772_ _09369_/A _10760_/X _10771_/X _09472_/A _19716_/Q vssd1 vssd1 vccd1 vccd1
+ _10798_/A sky130_fd_sc_hd__a32o_2
XFILLER_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12511_ _12953_/A vssd1 vssd1 vccd1 vccd1 _12511_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10642__A1 _10639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ _13491_/A vssd1 vssd1 vccd1 vccd1 _18344_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15230_ _15230_/A vssd1 vssd1 vccd1 vccd1 _15239_/S sky130_fd_sc_hd__buf_4
XFILLER_139_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ _12447_/A _12442_/B vssd1 vssd1 vccd1 vccd1 _12442_/Y sky130_fd_sc_hd__nor2_1
XFILLER_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12175__B _12175_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13986__S _13995_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ _19002_/Q _15083_/X _15167_/S vssd1 vssd1 vccd1 vccd1 _15162_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15767__A _15767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ _19356_/Q _12274_/B _15632_/S vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14112_ _13925_/X _18571_/Q _14118_/S vssd1 vssd1 vccd1 vccd1 _14113_/A sky130_fd_sc_hd__mux2_1
XFILLER_165_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09765__A _09765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11324_ _10779_/A _11323_/X _09563_/A vssd1 vssd1 vccd1 vccd1 _11324_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_154_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15486__B hold19/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15092_ _15092_/A vssd1 vssd1 vccd1 vccd1 _15092_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_158_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18920_ _19369_/CLK _18920_/D vssd1 vssd1 vccd1 vccd1 _18920_/Q sky130_fd_sc_hd__dfxtp_1
X_14043_ _18542_/Q _14042_/X _14043_/S vssd1 vssd1 vccd1 vccd1 _14044_/A sky130_fd_sc_hd__mux2_1
X_11255_ _19266_/Q _19104_/Q _18513_/Q _18283_/Q _09410_/A _11124_/X vssd1 vssd1 vccd1
+ vccd1 _11255_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17086__A1 _15600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10206_ _19319_/Q _18731_/Q _18768_/Q _18342_/Q _10166_/S _09891_/A vssd1 vssd1 vccd1
+ vccd1 _10206_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_90_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 _19529_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__10253__S0 _10247_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18851_ _19074_/CLK _18851_/D vssd1 vssd1 vccd1 vccd1 _18851_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11519__B _19844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ _11188_/A _11185_/X _11007_/X vssd1 vssd1 vccd1 vccd1 _11186_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16294__C1 _16293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17802_ _17802_/A _17802_/B vssd1 vssd1 vccd1 vccd1 _17802_/X sky130_fd_sc_hd__or2_1
XANTENNA__15706__S _15708_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10137_ _18503_/Q _18998_/Q _10137_/S vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__mux2_1
X_18782_ _19740_/CLK _18782_/D vssd1 vssd1 vccd1 vccd1 _18782_/Q sky130_fd_sc_hd__dfxtp_2
X_15994_ _13611_/X _19328_/Q _15996_/S vssd1 vssd1 vccd1 vccd1 _15995_/A sky130_fd_sc_hd__mux2_1
XFILLER_48_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17733_ _17733_/A _17733_/B vssd1 vssd1 vccd1 vccd1 _17733_/Y sky130_fd_sc_hd__nand2_1
X_14945_ _14945_/A vssd1 vssd1 vccd1 vccd1 _18918_/D sky130_fd_sc_hd__clkbuf_1
X_10068_ _19325_/Q _18737_/Q _18774_/Q _18348_/Q _10017_/S _09507_/A vssd1 vssd1 vccd1
+ vccd1 _10068_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10556__S1 _09443_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17664_ _17812_/A _17664_/B vssd1 vssd1 vccd1 vccd1 _17664_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14876_ _18886_/Q _13969_/X _14882_/S vssd1 vssd1 vccd1 vccd1 _14877_/A sky130_fd_sc_hd__mux2_1
XFILLER_62_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19403_ _19838_/CLK _19403_/D vssd1 vssd1 vccd1 vccd1 _19403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16615_ _19518_/Q _16613_/B _16614_/Y vssd1 vssd1 vccd1 vccd1 _19518_/D sky130_fd_sc_hd__o21a_1
XFILLER_165_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12607__C1 _12584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ _13311_/X _18476_/Q _13831_/S vssd1 vssd1 vccd1 vccd1 _13828_/A sky130_fd_sc_hd__mux2_1
XFILLER_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17595_ _19713_/Q _17570_/X _17594_/X vssd1 vssd1 vccd1 vccd1 _19713_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10308__S1 _09712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19334_ _19796_/CLK _19334_/D vssd1 vssd1 vccd1 vccd1 _19334_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__17222__A _17222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16546_ _16546_/A vssd1 vssd1 vccd1 vccd1 _16546_/X sky130_fd_sc_hd__clkbuf_2
X_13758_ _13349_/X _18446_/Q _13758_/S vssd1 vssd1 vccd1 vccd1 _13759_/A sky130_fd_sc_hd__mux2_1
XFILLER_16_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ _19448_/Q _12700_/X _12708_/X vssd1 vssd1 vccd1 vccd1 _12709_/X sky130_fd_sc_hd__o21a_1
X_19265_ _19329_/CLK _19265_/D vssd1 vssd1 vccd1 vccd1 _19265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16477_ _16868_/A vssd1 vssd1 vccd1 vccd1 _16524_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12366__A _19420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14057__S _14063_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ _13689_/A vssd1 vssd1 vccd1 vccd1 _18415_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18216_ _18224_/A _18216_/B vssd1 vssd1 vccd1 vccd1 _18217_/A sky130_fd_sc_hd__and2_1
XFILLER_129_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15428_ _15428_/A vssd1 vssd1 vccd1 vccd1 _19120_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_19_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19196_ _19386_/CLK _19196_/D vssd1 vssd1 vccd1 vccd1 _19196_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19250_/CLK sky130_fd_sc_hd__clkbuf_16
X_18147_ _16623_/A _18134_/X _18146_/X _16280_/X vssd1 vssd1 vccd1 vccd1 _19834_/D
+ sky130_fd_sc_hd__o211a_1
X_15359_ _19090_/Q _15057_/X _15361_/S vssd1 vssd1 vccd1 vccd1 _15360_/A sky130_fd_sc_hd__mux2_1
XFILLER_117_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_145_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18078_ _19806_/Q _12627_/X _18077_/X _17021_/X vssd1 vssd1 vccd1 vccd1 _19806_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_105_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09920_ _10158_/A _09920_/B vssd1 vssd1 vccd1 vccd1 _09920_/Y sky130_fd_sc_hd__nor2_1
X_17029_ _17085_/A vssd1 vssd1 vccd1 vccd1 _17098_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_116_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10614__A _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19286_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17077__A1 _15582_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ _10500_/S vssd1 vssd1 vccd1 vccd1 _10413_/S sky130_fd_sc_hd__clkbuf_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__A0 _19781_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _09782_/A vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__clkbuf_4
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16301__A _16301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11445__A _11445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11180__A _11195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _09331_/A _13944_/A _19701_/Q vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__o21ai_1
XFILLER_167_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12377__A1 _17125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09147_ _11589_/A _17108_/A _11530_/A vssd1 vssd1 vccd1 vccd1 _17166_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14491__A _14502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__A _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _19838_/Q _19837_/Q _19836_/Q _19835_/Q vssd1 vssd1 vccd1 vccd1 _09166_/B
+ sky130_fd_sc_hd__or4bb_2
XFILLER_107_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12129__A1 _19346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13326__A0 _19735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17068__A1 _12577_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _18390_/Q _18651_/Q _18550_/Q _18885_/Q _11265_/S _11033_/A vssd1 vssd1 vccd1
+ vccd1 _11041_/B sky130_fd_sc_hd__mux4_1
XFILLER_1_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09928__S0 _09840_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _19597_/Q _12697_/X _12503_/A _19465_/Q _12990_/X vssd1 vssd1 vccd1 vccd1
+ _15513_/B sky130_fd_sc_hd__a221o_2
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14730_ _14730_/A vssd1 vssd1 vccd1 vccd1 _18821_/D sky130_fd_sc_hd__clkbuf_1
X_11942_ _11942_/A vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_45_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17240__A1 _12383_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _14544_/X _18791_/Q _14665_/S vssd1 vssd1 vccd1 vccd1 _14662_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _11873_/A _17195_/A vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__or2_1
XFILLER_33_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18138__A _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16400_ _16427_/A _16406_/C vssd1 vssd1 vccd1 vccd1 _16400_/Y sky130_fd_sc_hd__nor2_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13570__A _15054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13612_ _18383_/Q _13611_/X _13615_/S vssd1 vssd1 vccd1 vccd1 _13613_/A sky130_fd_sc_hd__mux2_1
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10824_ _18617_/Q _18952_/Q _10824_/S vssd1 vssd1 vccd1 vccd1 _10824_/X sky130_fd_sc_hd__mux2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14592_/A vssd1 vssd1 vccd1 vccd1 _14592_/X sky130_fd_sc_hd__clkbuf_2
X_17380_ _17550_/S vssd1 vssd1 vccd1 vccd1 _17654_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__12604__A2 _17028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10076__C1 _09829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16331_ _19427_/Q _16331_/B _16331_/C vssd1 vssd1 vccd1 vccd1 _16332_/C sky130_fd_sc_hd__and3_1
X_13543_ _13543_/A vssd1 vssd1 vccd1 vccd1 _18361_/D sky130_fd_sc_hd__clkbuf_1
X_10755_ _11313_/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10755_/X sky130_fd_sc_hd__or2_1
XFILLER_125_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16262_ _16266_/A _16262_/B vssd1 vssd1 vccd1 vccd1 _16263_/A sky130_fd_sc_hd__or2_1
XFILLER_13_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19050_ _19247_/CLK _19050_/D vssd1 vssd1 vccd1 vccd1 _19050_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_20_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13474_ _13474_/A vssd1 vssd1 vccd1 vccd1 _18336_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17696__B _17696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10686_ _10590_/A _10685_/X _09630_/X vssd1 vssd1 vccd1 vccd1 _10686_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_127_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15213_ _19025_/Q _15054_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15214_/A sky130_fd_sc_hd__mux2_1
X_18001_ _19773_/Q _19394_/Q _18005_/S vssd1 vssd1 vccd1 vccd1 _18002_/A sky130_fd_sc_hd__mux2_1
X_12425_ _17917_/B _17232_/A vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__or2_1
XFILLER_173_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16193_ _16239_/S vssd1 vssd1 vccd1 vccd1 _16202_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_154_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15144_ _15144_/A vssd1 vssd1 vccd1 vccd1 _18994_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10474__S0 _10274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12356_ _17886_/B _12356_/B vssd1 vssd1 vccd1 vccd1 _12360_/A sky130_fd_sc_hd__xnor2_1
XFILLER_153_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ _11307_/A _11307_/B _11307_/C vssd1 vssd1 vccd1 vccd1 _11307_/X sky130_fd_sc_hd__or3_4
XFILLER_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15075_ _15075_/A vssd1 vssd1 vccd1 vccd1 _18967_/D sky130_fd_sc_hd__clkbuf_1
X_12287_ _12287_/A _17856_/B vssd1 vssd1 vccd1 vccd1 _12314_/A sky130_fd_sc_hd__nor2_1
XFILLER_141_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17059__A1 _15536_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ _14598_/A vssd1 vssd1 vccd1 vccd1 _14026_/X sky130_fd_sc_hd__clkbuf_2
X_18903_ _19127_/CLK _18903_/D vssd1 vssd1 vccd1 vccd1 _18903_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_output74_A _11968_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ _11238_/A vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__buf_4
XFILLER_171_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15436__S _15444_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18834_ _19378_/CLK _18834_/D vssd1 vssd1 vccd1 vccd1 _18834_/Q sky130_fd_sc_hd__dfxtp_1
X_11169_ _09477_/A _11158_/X _11167_/X _09577_/A _11168_/Y vssd1 vssd1 vccd1 vccd1
+ _12445_/B sky130_fd_sc_hd__o32ai_4
XFILLER_96_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18765_ _19378_/CLK _18765_/D vssd1 vssd1 vccd1 vccd1 _18765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15977_ _13586_/X _19320_/Q _15981_/S vssd1 vssd1 vccd1 vccd1 _15978_/A sky130_fd_sc_hd__mux2_1
XFILLER_82_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17716_ _17551_/X _17549_/Y _17716_/S vssd1 vssd1 vccd1 vccd1 _17716_/X sky130_fd_sc_hd__mux2_1
X_14928_ _18910_/Q _14045_/X _14930_/S vssd1 vssd1 vccd1 vccd1 _14929_/A sky130_fd_sc_hd__mux2_1
X_18696_ _19285_/CLK _18696_/D vssd1 vssd1 vccd1 vccd1 _18696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17231__A1 _12405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _17370_/X _17359_/Y _17716_/S vssd1 vssd1 vccd1 vccd1 _17647_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12795__S _13144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14859_ _14859_/A vssd1 vssd1 vccd1 vccd1 _18879_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15171__S _15171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17578_ _17574_/Y _17577_/X _17625_/S vssd1 vssd1 vccd1 vccd1 _17578_/X sky130_fd_sc_hd__mux2_1
XFILLER_91_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14295__B _18224_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19317_ _19379_/CLK _19317_/D vssd1 vssd1 vccd1 vccd1 _19317_/Q sky130_fd_sc_hd__dfxtp_1
X_16529_ _19491_/Q _16529_/B _16529_/C vssd1 vssd1 vccd1 vccd1 _16530_/C sky130_fd_sc_hd__and3_1
XFILLER_31_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19248_ _19248_/CLK _19248_/D vssd1 vssd1 vccd1 vccd1 _19248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19179_ _19180_/CLK _19179_/D vssd1 vssd1 vccd1 vccd1 _19179_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14515__S _14515_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11031__A1 _18981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12543__B _12543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ _10205_/A vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__buf_2
XFILLER_113_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15346__S _15350_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13655__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10768__S1 _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09834_ _09834_/A vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__clkbuf_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09765_/A vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__buf_2
XFILLER_67_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09696_ _10150_/A vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15081__S _15093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_109_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10058__C1 _10689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ _09761_/A _10529_/X _10538_/X _09834_/A _10539_/Y vssd1 vssd1 vccd1 vccd1
+ _12462_/A sky130_fd_sc_hd__o32a_4
XANTENNA__11270__A1 _11024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16733__B1 _16718_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_194_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10471_ _10471_/A _10471_/B vssd1 vssd1 vccd1 vccd1 _10471_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12210_ _11619_/A _11507_/A _12302_/A vssd1 vssd1 vccd1 vccd1 _12210_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_109_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13190_ _15063_/A vssd1 vssd1 vccd1 vccd1 _14585_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_135_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10376__A3 _10375_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12141_ _12241_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12142_/B sky130_fd_sc_hd__nor2_1
XFILLER_68_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10781__B1 _09484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10208__S0 _09955_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12072_ _19344_/Q _12069_/X _12071_/X vssd1 vssd1 vccd1 vccd1 _12072_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15900_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15909_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__09923__C1 _09831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15256__S _15256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _11116_/A _11021_/X _11022_/X vssd1 vssd1 vccd1 vccd1 _11023_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_150_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16880_ _16879_/B _16879_/C _19605_/Q vssd1 vssd1 vccd1 vccd1 _16881_/C sky130_fd_sc_hd__a21oi_1
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10533__B1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15831_ _13583_/X _19255_/Q _15837_/S vssd1 vssd1 vccd1 vccd1 _15832_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15472__A0 _15471_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11085__A _11085_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18550_ _19076_/CLK _18550_/D vssd1 vssd1 vccd1 vccd1 _18550_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15762_ _15762_/A vssd1 vssd1 vccd1 vccd1 _19224_/D sky130_fd_sc_hd__clkbuf_1
X_12974_ _12974_/A vssd1 vssd1 vccd1 vccd1 _12974_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17213__A1 _12089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17501_ _17340_/A _17345_/Y _17501_/S vssd1 vssd1 vccd1 vccd1 _17609_/B sky130_fd_sc_hd__mux2_1
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _14620_/X _18815_/Q _14713_/S vssd1 vssd1 vccd1 vccd1 _14714_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _19736_/CLK _18481_/D vssd1 vssd1 vccd1 vccd1 _18481_/Q sky130_fd_sc_hd__dfxtp_1
X_11925_ _11924_/Y _11456_/A _11925_/S vssd1 vssd1 vccd1 vccd1 _17201_/A sky130_fd_sc_hd__mux2_2
XFILLER_75_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _14598_/X _19194_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15694_/A sky130_fd_sc_hd__mux2_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17432_/A _17432_/B _17190_/A vssd1 vssd1 vccd1 vccd1 _17871_/A sky130_fd_sc_hd__or3b_1
XANTENNA__11813__A _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11856_ _19400_/Q vssd1 vssd1 vccd1 vccd1 _11879_/A sky130_fd_sc_hd__buf_4
X_14644_ _14700_/A vssd1 vssd1 vccd1 vccd1 _14713_/S sky130_fd_sc_hd__buf_6
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10049__C1 _09752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _10807_/A vssd1 vssd1 vccd1 vccd1 _10953_/A sky130_fd_sc_hd__clkbuf_2
X_14575_ _14575_/A vssd1 vssd1 vccd1 vccd1 _18763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17363_ _17361_/X _17362_/X _17497_/S vssd1 vssd1 vccd1 vccd1 _17364_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11787_ _11822_/A _17247_/A vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__xnor2_4
XFILLER_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19102_ _19296_/CLK _19102_/D vssd1 vssd1 vccd1 vccd1 _19102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16314_ _19473_/Q _19472_/Q _19474_/Q _16461_/A vssd1 vssd1 vccd1 vccd1 _16469_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10738_ _19180_/Q _18794_/Q _19244_/Q _18363_/Q _10654_/A _10655_/A vssd1 vssd1 vccd1
+ vccd1 _10739_/B sky130_fd_sc_hd__mux4_2
XFILLER_13_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13526_ _18356_/Q _13525_/X _13529_/S vssd1 vssd1 vccd1 vccd1 _13527_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10695__S0 _10576_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17294_ _17292_/X _17293_/X _17294_/S vssd1 vssd1 vccd1 vccd1 _17294_/X sky130_fd_sc_hd__mux2_1
XFILLER_158_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_174_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19033_ _19385_/CLK _19033_/D vssd1 vssd1 vccd1 vccd1 _19033_/Q sky130_fd_sc_hd__dfxtp_1
X_16245_ _16245_/A vssd1 vssd1 vccd1 vccd1 _16848_/A sky130_fd_sc_hd__buf_4
X_13457_ _12981_/X _18329_/Q _13459_/S vssd1 vssd1 vccd1 vccd1 _13458_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14335__S _14343_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ _10669_/A _10669_/B vssd1 vssd1 vccd1 vccd1 _10669_/X sky130_fd_sc_hd__and2_1
XFILLER_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11013__A1 _19109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _12408_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12408_/X sky130_fd_sc_hd__xor2_4
XFILLER_115_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16176_ _13522_/X _19362_/Q _16180_/S vssd1 vssd1 vccd1 vccd1 _16177_/A sky130_fd_sc_hd__mux2_1
X_13388_ _13388_/A vssd1 vssd1 vccd1 vccd1 _18314_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput106 _17166_/A vssd1 vssd1 vccd1 vccd1 io_dbus_rd_en sky130_fd_sc_hd__buf_2
XFILLER_115_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput117 _12465_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[17] sky130_fd_sc_hd__buf_2
XFILLER_154_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10998__S1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15127_ _15127_/A vssd1 vssd1 vccd1 vccd1 _18986_/D sky130_fd_sc_hd__clkbuf_1
X_12339_ _19418_/Q _19419_/Q _12339_/C vssd1 vssd1 vccd1 vccd1 _12371_/B sky130_fd_sc_hd__and3_1
Xoutput128 _12477_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[27] sky130_fd_sc_hd__buf_2
XFILLER_114_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput139 _12453_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[8] sky130_fd_sc_hd__buf_2
XFILLER_115_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15058_ _18962_/Q _15057_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15059_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_123_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14009_ _14009_/A vssd1 vssd1 vccd1 vccd1 _18531_/D sky130_fd_sc_hd__clkbuf_1
X_19866_ _19866_/CLK _19866_/D vssd1 vssd1 vccd1 vccd1 _19866_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14070__S _14074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10524__B1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18817_ _19235_/CLK _18817_/D vssd1 vssd1 vccd1 vccd1 _18817_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19797_ _19800_/CLK _19797_/D vssd1 vssd1 vccd1 vccd1 _19797_/Q sky130_fd_sc_hd__dfxtp_1
X_09550_ _09803_/A _09544_/X _09549_/X vssd1 vssd1 vccd1 vccd1 _09550_/Y sky130_fd_sc_hd__o21ai_1
X_18748_ _19235_/CLK _18748_/D vssd1 vssd1 vccd1 vccd1 _18748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17204__A1 _17802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10827__A1 _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09481_ _09481_/A vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18679_ _19724_/CLK _18679_/D vssd1 vssd1 vccd1 vccd1 _18679_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_149_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10438__S0 _10341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10212__C1 _09831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10802__A _11174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09748_ _18477_/Q _19068_/Q _19230_/Q _18445_/Q _11374_/S _09687_/A vssd1 vssd1 vccd1
+ vccd1 _09748_/X sky130_fd_sc_hd__mux4_1
XFILLER_28_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__A1 _19112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ _09980_/S vssd1 vssd1 vccd1 vccd1 _10451_/S sky130_fd_sc_hd__buf_2
XFILLER_28_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12729__A _12769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17746__A2 _17743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ _11810_/S _11706_/X _11707_/Y _11709_/X vssd1 vssd1 vccd1 vccd1 _11710_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ _12689_/X _12675_/X _12716_/S vssd1 vssd1 vccd1 vccd1 _12690_/X sky130_fd_sc_hd__mux2_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12448__B _12448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11738_/A vssd1 vssd1 vccd1 vccd1 _12100_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14360_ _14360_/A vssd1 vssd1 vccd1 vccd1 _18672_/D sky130_fd_sc_hd__clkbuf_1
X_11572_ _11542_/A _11918_/B _11571_/Y _09341_/A vssd1 vssd1 vccd1 vccd1 _11572_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15509__B2 hold12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ _14608_/A vssd1 vssd1 vccd1 vccd1 _13311_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10523_ _18927_/Q _18693_/Q _19375_/Q _19023_/Q _10520_/S _10262_/A vssd1 vssd1 vccd1
+ vccd1 _10523_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput19 io_dbus_rdata[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_2
X_14291_ _14291_/A vssd1 vssd1 vccd1 vccd1 _18644_/D sky130_fd_sc_hd__clkbuf_1
X_13242_ _13242_/A vssd1 vssd1 vccd1 vccd1 _18306_/D sky130_fd_sc_hd__clkbuf_1
X_16030_ _16086_/A vssd1 vssd1 vccd1 vccd1 _16052_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10454_ _10500_/S vssd1 vssd1 vccd1 vccd1 _10499_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__12743__A1 _18258_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _13173_/A vssd1 vssd1 vccd1 vccd1 _18302_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_123_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10385_ _18595_/Q _18866_/Q _19090_/Q _18834_/Q _10339_/S _10482_/A vssd1 vssd1 vccd1
+ vccd1 _10385_/X sky130_fd_sc_hd__mux4_1
XFILLER_163_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _19410_/Q vssd1 vssd1 vccd1 vccd1 _12126_/A sky130_fd_sc_hd__buf_2
XANTENNA__15494__B hold15/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17981_ _17981_/A vssd1 vssd1 vccd1 vccd1 _17990_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_111_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19720_ _19720_/CLK _19720_/D vssd1 vssd1 vccd1 vccd1 _19720_/Q sky130_fd_sc_hd__dfxtp_4
X_16932_ _16932_/A _16931_/X vssd1 vssd1 vccd1 vccd1 _16932_/X sky130_fd_sc_hd__or2b_1
X_12055_ _19787_/Q _10494_/A _12143_/S vssd1 vssd1 vccd1 vccd1 _12089_/A sky130_fd_sc_hd__mux2_4
XFILLER_96_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11006_ _19303_/Q _18715_/Q _18752_/Q _18326_/Q _10940_/S _11005_/X vssd1 vssd1 vccd1
+ vccd1 _11006_/X sky130_fd_sc_hd__mux4_1
X_19651_ _19687_/CLK _19651_/D vssd1 vssd1 vccd1 vccd1 _19651_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16863_ _16862_/B _16862_/C _19599_/Q vssd1 vssd1 vccd1 vccd1 _16864_/C sky130_fd_sc_hd__a21oi_1
XFILLER_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18602_ _19197_/CLK _18602_/D vssd1 vssd1 vccd1 vccd1 _18602_/Q sky130_fd_sc_hd__dfxtp_1
X_15814_ _15814_/A vssd1 vssd1 vccd1 vccd1 _19247_/D sky130_fd_sc_hd__clkbuf_1
X_19582_ _19635_/CLK _19582_/D vssd1 vssd1 vccd1 vccd1 _19582_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16794_ _19572_/Q vssd1 vssd1 vccd1 vccd1 _16800_/B sky130_fd_sc_hd__clkbuf_1
X_18533_ _19027_/CLK _18533_/D vssd1 vssd1 vccd1 vccd1 _18533_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_93_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15745_ _15767_/A vssd1 vssd1 vccd1 vccd1 _15754_/S sky130_fd_sc_hd__clkbuf_8
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _19146_/Q _12956_/B _12956_/Y vssd1 vssd1 vccd1 vccd1 _12957_/X sky130_fd_sc_hd__o21a_1
XFILLER_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15015__A _15015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18464_ _19249_/CLK _18464_/D vssd1 vssd1 vccd1 vccd1 _18464_/Q sky130_fd_sc_hd__dfxtp_1
X_11908_ _11934_/B _11908_/B vssd1 vssd1 vccd1 vccd1 _11908_/Y sky130_fd_sc_hd__nand2_1
X_15676_ _14573_/X _19186_/Q _15682_/S vssd1 vssd1 vccd1 vccd1 _15677_/A sky130_fd_sc_hd__mux2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12888_/A vssd1 vssd1 vccd1 vccd1 _18287_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17415_ _17415_/A _17726_/B vssd1 vssd1 vccd1 vccd1 _17603_/A sky130_fd_sc_hd__nor2_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14627_ _14627_/A vssd1 vssd1 vccd1 vccd1 _18148_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_18395_ _19311_/CLK _18395_/D vssd1 vssd1 vccd1 vccd1 _18395_/Q sky130_fd_sc_hd__dfxtp_1
X_11839_ _11893_/A vssd1 vssd1 vccd1 vccd1 _17630_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18147__C1 _16280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16772__C _16772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17230__A _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11234__A1 _11024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17346_ _17356_/S _17346_/B vssd1 vssd1 vccd1 vccd1 _17346_/X sky130_fd_sc_hd__and2b_1
X_14558_ _14557_/X _18758_/Q _14567_/S vssd1 vssd1 vccd1 vccd1 _14559_/A sky130_fd_sc_hd__mux2_1
XFILLER_174_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _14996_/A vssd1 vssd1 vccd1 vccd1 _13509_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_173_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17277_ _17275_/X _17276_/X _17375_/S vssd1 vssd1 vccd1 vccd1 _17277_/X sky130_fd_sc_hd__mux2_1
XFILLER_174_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14489_ _13902_/X _18729_/Q _14489_/S vssd1 vssd1 vccd1 vccd1 _14490_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19016_ _19113_/CLK _19016_/D vssd1 vssd1 vccd1 vccd1 _19016_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_134_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16228_ _16228_/A vssd1 vssd1 vccd1 vccd1 _19385_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_161_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16159_ _16159_/A _19769_/Q _16159_/C vssd1 vssd1 vccd1 vccd1 _16165_/B sky130_fd_sc_hd__or3_1
XFILLER_138_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10745__B1 _09448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10840__S0 _10854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11718__A _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10622__A _10689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_142_clock_A clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19849_ _19865_/CLK _19849_/D vssd1 vssd1 vccd1 vccd1 _19849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09602_ _09989_/A vssd1 vssd1 vccd1 vccd1 _09602_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09533_ _10839_/A vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__buf_2
XANTENNA__12549__A _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13144__S _13144_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09464_ _09464_/A vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12670__B1 _17102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09395_ _09589_/A vssd1 vssd1 vccd1 vccd1 _09688_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17140__A _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__A2 _10012_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_67_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11084__S0 _10964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14703__S _14709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10170_ _10115_/A _10167_/Y _10169_/Y _09964_/A vssd1 vssd1 vccd1 vccd1 _10170_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_106_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_120_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11347__B _12462_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17315__A _17485_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13860_ _13860_/A vssd1 vssd1 vccd1 vccd1 _18486_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11139__S1 _11124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12811_ _13275_/A vssd1 vssd1 vccd1 vccd1 _13387_/S sky130_fd_sc_hd__buf_6
XFILLER_28_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13791_ _13791_/A vssd1 vssd1 vccd1 vccd1 _18459_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12459__A _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09657__A1 _10680_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15530_ _15530_/A vssd1 vssd1 vccd1 vccd1 _19149_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ hold15/A _12739_/X _11288_/A _12740_/X vssd1 vssd1 vccd1 vccd1 _18257_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13989__S _13995_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15461_ _09309_/X _13404_/X _15482_/S vssd1 vssd1 vccd1 vccd1 _15461_/X sky130_fd_sc_hd__mux2_1
X_12673_ _13392_/A vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18146__A _18146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_169_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17200_ _17197_/X _17199_/X _17336_/A vssd1 vssd1 vccd1 vccd1 _17440_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14412_ _14412_/A vssd1 vssd1 vccd1 vccd1 _18694_/D sky130_fd_sc_hd__clkbuf_1
X_11624_ _11623_/X _11553_/Y _19393_/Q vssd1 vssd1 vccd1 vccd1 _11624_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18180_ _18190_/A _18180_/B vssd1 vssd1 vccd1 vccd1 _18181_/A sky130_fd_sc_hd__and2_1
XANTENNA__09768__A _09768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15392_ _19104_/Q _14996_/X _15400_/S vssd1 vssd1 vccd1 vccd1 _15393_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17131_ _18142_/B _17177_/B _17131_/C _17131_/D vssd1 vssd1 vccd1 vccd1 _17131_/Y
+ sky130_fd_sc_hd__nor4_4
X_14343_ _13902_/X _18665_/Q _14343_/S vssd1 vssd1 vccd1 vccd1 _14344_/A sky130_fd_sc_hd__mux2_1
XFILLER_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11555_ _11565_/A _11513_/A _09327_/A _18104_/A vssd1 vssd1 vccd1 vccd1 _17917_/A
+ sky130_fd_sc_hd__o211a_4
XFILLER_156_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10506_ _10511_/A _10503_/X _10505_/X _09737_/A vssd1 vssd1 vccd1 vccd1 _10506_/X
+ sky130_fd_sc_hd__o211a_1
X_17062_ _17062_/A vssd1 vssd1 vccd1 vccd1 _19678_/D sky130_fd_sc_hd__clkbuf_1
X_14274_ _18197_/A vssd1 vssd1 vccd1 vccd1 _14274_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_171_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11486_ _11412_/A _11492_/D _11485_/X vssd1 vssd1 vccd1 vccd1 _11489_/B sky130_fd_sc_hd__a21oi_1
XFILLER_155_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13913__A0 _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16013_ _16021_/C _16013_/B vssd1 vssd1 vccd1 vccd1 _16013_/Y sky130_fd_sc_hd__nand2_1
X_13225_ input15/X _13166_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _13225_/Y sky130_fd_sc_hd__a21oi_2
X_10437_ _10275_/X _10434_/Y _10436_/Y _10429_/A vssd1 vssd1 vccd1 vccd1 _10437_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17104__B1 _18091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13156_ _19475_/Q vssd1 vssd1 vccd1 vccd1 _16474_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10368_ _18499_/Q _18994_/Q _10368_/S vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__mux2_1
XFILLER_98_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10822__S0 _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _19409_/Q _12093_/X _12103_/X _12106_/Y vssd1 vssd1 vccd1 vccd1 _16282_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__13229__S _13252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13154_/A _13082_/X _13086_/Y _13051_/A vssd1 vssd1 vccd1 vccd1 _13088_/B
+ sky130_fd_sc_hd__a211o_1
X_17964_ _16091_/A _19788_/Q _17968_/S vssd1 vssd1 vccd1 vccd1 _17965_/A sky130_fd_sc_hd__mux2_1
X_10299_ _10288_/Y _10292_/Y _10294_/Y _10298_/Y _09831_/A vssd1 vssd1 vccd1 vccd1
+ _10299_/X sky130_fd_sc_hd__o221a_4
XFILLER_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19703_ _19706_/CLK _19703_/D vssd1 vssd1 vccd1 vccd1 _19703_/Q sky130_fd_sc_hd__dfxtp_1
X_16915_ _16915_/A _16915_/B vssd1 vssd1 vccd1 vccd1 _16915_/Y sky130_fd_sc_hd__nor2_1
X_12038_ _12066_/A _12066_/C vssd1 vssd1 vccd1 vccd1 _12040_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11378__S1 _09715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17895_ _19735_/Q _17831_/X _17894_/X vssd1 vssd1 vccd1 vccd1 _19735_/D sky130_fd_sc_hd__o21a_1
XANTENNA__15444__S _15444_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19634_ _19635_/CLK _19634_/D vssd1 vssd1 vccd1 vccd1 _19634_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18080__A1 _09172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16846_ _16845_/B _16845_/C _19593_/Q vssd1 vssd1 vccd1 vccd1 _16847_/C sky130_fd_sc_hd__a21oi_1
XFILLER_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09360__A3 _17112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19565_ _19667_/CLK _19565_/D vssd1 vssd1 vccd1 vccd1 _19565_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_168_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16777_ _19567_/Q vssd1 vssd1 vccd1 vccd1 _16777_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13989_ _18525_/Q _13988_/X _13995_/S vssd1 vssd1 vccd1 vccd1 _13990_/A sky130_fd_sc_hd__mux2_1
X_18516_ _19108_/CLK _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10258__A2 _10245_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15728_ _13538_/X _19209_/Q _15732_/S vssd1 vssd1 vccd1 vccd1 _15729_/A sky130_fd_sc_hd__mux2_1
X_19496_ _19619_/CLK _19496_/D vssd1 vssd1 vccd1 vccd1 _19496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10663__C1 _09614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18447_ _19390_/CLK _18447_/D vssd1 vssd1 vccd1 vccd1 _18447_/Q sky130_fd_sc_hd__dfxtp_1
X_15659_ _15659_/A vssd1 vssd1 vccd1 vccd1 _19178_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09678__A _09733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ _18102_/A _09186_/B _09180_/C _17124_/B vssd1 vssd1 vccd1 vccd1 _11526_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18378_ _19391_/CLK _18378_/D vssd1 vssd1 vccd1 vccd1 _18378_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17329_ _12488_/Y _17328_/B _09322_/X vssd1 vssd1 vccd1 vccd1 _17329_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17894__A1 _12369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14523__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16304__A _18079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13139__S _13172_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10733__A3 _18826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15409__A0 _19112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_68_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10041__S1 _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16082__A0 _12550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ _09547_/A vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__buf_2
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09447_ _09447_/A vssd1 vssd1 vccd1 vccd1 _09448_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_169_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13199__A1 _19159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13199__B2 _19349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ _09416_/A vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11340_ _09617_/X _11329_/X _11338_/X _09579_/A _11339_/Y vssd1 vssd1 vccd1 vccd1
+ _12460_/A sky130_fd_sc_hd__o32a_4
XFILLER_166_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13838__A _19811_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11271_ _11278_/A _11268_/X _11270_/X vssd1 vssd1 vccd1 vccd1 _11271_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_152_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14433__S _14439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ _19674_/Q _13008_/X _13009_/X _16967_/A vssd1 vssd1 vccd1 vccd1 _13010_/X
+ sky130_fd_sc_hd__a22o_1
X_10222_ _10345_/A _10221_/X _09765_/A vssd1 vssd1 vccd1 vccd1 _10222_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17637__A1 _19715_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13371__A1 _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13049__S _13091_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _10197_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10153_/X sky130_fd_sc_hd__or2_1
XFILLER_0_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input36_A io_ibus_inst[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14961_ _14961_/A vssd1 vssd1 vccd1 vccd1 _18926_/D sky130_fd_sc_hd__clkbuf_1
X_10084_ _11427_/A _11426_/A vssd1 vssd1 vccd1 vccd1 _10084_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16700_ _16706_/C _16706_/D _16675_/X vssd1 vssd1 vccd1 vccd1 _16700_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13573__A _15057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13912_ _14592_/A vssd1 vssd1 vccd1 vccd1 _13912_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__A0 _19711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17680_ _17680_/A _17680_/B vssd1 vssd1 vccd1 vccd1 _17680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14892_ _14892_/A vssd1 vssd1 vccd1 vccd1 _18893_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16631_ _19521_/Q _19520_/Q vssd1 vssd1 vccd1 vccd1 _16659_/B sky130_fd_sc_hd__and2_1
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10893__C1 _10883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13843_ _13837_/X _18481_/Q _13855_/S vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__mux2_1
XFILLER_90_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11093__A _19711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19350_ _19357_/CLK _19350_/D vssd1 vssd1 vccd1 vccd1 _19350_/Q sky130_fd_sc_hd__dfxtp_2
X_16562_ _16570_/A _16567_/C vssd1 vssd1 vccd1 vccd1 _16562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13774_ _12865_/X _18452_/Q _13776_/S vssd1 vssd1 vccd1 vccd1 _13775_/A sky130_fd_sc_hd__mux2_1
X_10986_ _09617_/A _10975_/X _10984_/X _09578_/A _10985_/Y vssd1 vssd1 vccd1 vccd1
+ _12449_/B sky130_fd_sc_hd__o32a_4
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18301_ _19284_/CLK _18301_/D vssd1 vssd1 vccd1 vccd1 _18301_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17022__C1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15513_ hold18/A _15513_/B vssd1 vssd1 vccd1 vccd1 _15513_/X sky130_fd_sc_hd__or2_1
X_19281_ _19282_/CLK _19281_/D vssd1 vssd1 vccd1 vccd1 _19281_/Q sky130_fd_sc_hd__dfxtp_1
X_12725_ _18252_/Q _12724_/X _17520_/S vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__mux2_1
X_16493_ _16493_/A _19482_/Q _16493_/C vssd1 vssd1 vccd1 vccd1 _16495_/B sky130_fd_sc_hd__and3_1
XFILLER_30_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18232_ _18232_/A vssd1 vssd1 vccd1 vccd1 _19861_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09498__A _11318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15444_ _19128_/Q _15076_/X _15444_/S vssd1 vssd1 vccd1 vccd1 _15445_/A sky130_fd_sc_hd__mux2_1
X_12656_ _16341_/A _19586_/Q _16921_/S _12655_/X vssd1 vssd1 vccd1 vccd1 _19586_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_31_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18163_ _18163_/A _18163_/B vssd1 vssd1 vccd1 vccd1 _18164_/A sky130_fd_sc_hd__or2_1
X_11607_ _11607_/A _11607_/B _17230_/A vssd1 vssd1 vccd1 vccd1 _11608_/B sky130_fd_sc_hd__or3_1
XFILLER_90_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12587_ _19442_/Q _12584_/Y _13356_/B _19474_/Q _12586_/X vssd1 vssd1 vccd1 vccd1
+ _12587_/X sky130_fd_sc_hd__a221o_1
XFILLER_129_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15375_ _19097_/Q _15079_/X _15383_/S vssd1 vssd1 vccd1 vccd1 _15376_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17114_ _17114_/A _17120_/B _17114_/C vssd1 vssd1 vccd1 vccd1 _17114_/X sky130_fd_sc_hd__and3_1
XFILLER_117_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14326_ _13877_/X _18657_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14327_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18094_ _19845_/Q _18116_/B vssd1 vssd1 vccd1 vccd1 _18094_/X sky130_fd_sc_hd__or2_1
XFILLER_129_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11538_ _13051_/A vssd1 vssd1 vccd1 vccd1 _11538_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_7_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17045_ _17045_/A vssd1 vssd1 vccd1 vccd1 _19670_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14343__S _14343_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14257_ _14257_/A vssd1 vssd1 vccd1 vccd1 _18634_/D sky130_fd_sc_hd__clkbuf_1
X_11469_ _10082_/X _10083_/B _11468_/X _11418_/Y vssd1 vssd1 vccd1 vccd1 _11469_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12652__A _15632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ _15067_/A vssd1 vssd1 vccd1 vccd1 _14589_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10176__A1 _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14188_ _14188_/A vssd1 vssd1 vccd1 vccd1 _18604_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13139_ _13138_/X _18300_/Q _13172_/S vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__mux2_1
XFILLER_124_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16300__A1 _12321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18996_ _19089_/CLK _18996_/D vssd1 vssd1 vccd1 vccd1 _18996_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09581__A3 _09573_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16778__B _19565_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17947_ _17947_/A vssd1 vssd1 vccd1 vccd1 _19748_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_15_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13483__A _13494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18053__A1 _19417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__S1 _09651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17878_ _17878_/A _17878_/B vssd1 vssd1 vccd1 vccd1 _17878_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10900__A _10965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16829_ _16829_/A vssd1 vssd1 vccd1 vccd1 _19582_/D sky130_fd_sc_hd__clkbuf_1
X_19617_ _19618_/CLK _19617_/D vssd1 vssd1 vccd1 vccd1 _19617_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10884__C1 _10883_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15811__A0 _13554_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19548_ _19549_/CLK _19548_/D vssd1 vssd1 vccd1 vccd1 _19548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09716__S1 _09715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09301_ _09301_/A _09301_/B vssd1 vssd1 vccd1 vccd1 _11551_/A sky130_fd_sc_hd__or2_2
XFILLER_80_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19479_ _19610_/CLK _19479_/D vssd1 vssd1 vccd1 vccd1 _19479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14378__A0 _13845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09232_ _19698_/Q vssd1 vssd1 vccd1 vccd1 _13400_/A sky130_fd_sc_hd__buf_4
XFILLER_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ _11528_/C vssd1 vssd1 vccd1 vccd1 _17114_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__10347__A _10347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17316__B1 _17294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09094_ _09174_/A _09174_/B vssd1 vssd1 vccd1 vccd1 _11513_/C sky130_fd_sc_hd__and2_1
XFILLER_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_135_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10082__A _10082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09996_ _09998_/A _09994_/X _09995_/X vssd1 vssd1 vccd1 vccd1 _09996_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14302__A0 _13837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09871__A _09871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15084__S _15093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18044__A1 _19413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11667__A1 _19394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11906__A _11915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15802__A0 _13541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10840_ _19274_/Q _19112_/Q _18521_/Q _18291_/Q _10854_/S _10837_/X vssd1 vssd1 vccd1
+ vccd1 _10840_/X sky130_fd_sc_hd__mux4_1
XANTENNA__12616__B1 _12714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13840__B _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17312__B _17319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ _09434_/A _10762_/X _10766_/X _10770_/X _09374_/A vssd1 vssd1 vccd1 vccd1
+ _10771_/X sky130_fd_sc_hd__a311o_2
XANTENNA__14428__S _14428_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12510_ _13054_/A vssd1 vssd1 vccd1 vccd1 _12953_/A sky130_fd_sc_hd__clkbuf_2
X_13490_ _13240_/X _18344_/Q _13492_/S vssd1 vssd1 vccd1 vccd1 _13491_/A sky130_fd_sc_hd__mux2_1
XFILLER_139_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _19423_/Q _12319_/X _12437_/X _12440_/Y vssd1 vssd1 vccd1 vccd1 _12441_/X
+ sky130_fd_sc_hd__o22a_4
XANTENNA__13041__A0 _19719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12372_ _12372_/A _12372_/B _12410_/C vssd1 vssd1 vccd1 vccd1 _12372_/X sky130_fd_sc_hd__or3_1
X_15160_ _15160_/A vssd1 vssd1 vccd1 vccd1 _19001_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_166_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11323_ _18925_/Q _18691_/Q _19373_/Q _19021_/Q _09519_/A _09506_/A vssd1 vssd1 vccd1
+ vccd1 _11323_/X sky130_fd_sc_hd__mux4_1
X_14111_ _14111_/A vssd1 vssd1 vccd1 vccd1 _18570_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15091_ _15091_/A vssd1 vssd1 vccd1 vccd1 _18972_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14163__S _14169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11254_ _11254_/A _11254_/B vssd1 vssd1 vccd1 vccd1 _11254_/X sky130_fd_sc_hd__or2_1
X_14042_ _14614_/A vssd1 vssd1 vccd1 vccd1 _14042_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_109_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09643__S0 _10572_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10205_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10205_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18850_ _19074_/CLK _18850_/D vssd1 vssd1 vccd1 vccd1 _18850_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15783__A _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10253__S1 _10238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11185_ _19301_/Q _18713_/Q _18750_/Q _18324_/Q _10873_/S _11177_/X vssd1 vssd1 vccd1
+ vccd1 _11185_/X sky130_fd_sc_hd__mux4_1
XFILLER_79_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11519__C _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17801_ _17724_/A _17798_/X _17800_/Y _17413_/A vssd1 vssd1 vccd1 vccd1 _17801_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_121_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10136_ _18934_/Q _18700_/Q _19382_/Q _19030_/Q _09846_/X _09871_/X vssd1 vssd1 vccd1
+ vccd1 _10136_/X sky130_fd_sc_hd__mux4_1
XFILLER_122_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18781_ _19711_/CLK _18781_/D vssd1 vssd1 vccd1 vccd1 _18781_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15993_ _15993_/A vssd1 vssd1 vccd1 vccd1 _19327_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_95_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13507__S _13507_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ _17400_/X _17731_/X _17732_/S vssd1 vssd1 vccd1 vccd1 _17733_/B sky130_fd_sc_hd__mux2_1
XFILLER_76_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11658__A1 _19627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14944_ _18918_/Q vssd1 vssd1 vccd1 vccd1 _14945_/A sky130_fd_sc_hd__clkbuf_1
X_10067_ _10684_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _10067_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_189_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10866__C1 _09658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17663_ _17661_/X _17664_/B _17744_/S vssd1 vssd1 vccd1 vccd1 _17663_/X sky130_fd_sc_hd__mux2_1
XFILLER_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14875_ _14875_/A vssd1 vssd1 vccd1 vccd1 _18885_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19402_ _19838_/CLK _19402_/D vssd1 vssd1 vccd1 vccd1 _19402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16614_ _16666_/A _16614_/B vssd1 vssd1 vccd1 vccd1 _16614_/Y sky130_fd_sc_hd__nor2_1
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12607__B1 _12606_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13826_ _13826_/A vssd1 vssd1 vccd1 vccd1 _18475_/D sky130_fd_sc_hd__clkbuf_1
X_17594_ _11796_/A _17427_/X _17593_/X _09359_/X vssd1 vssd1 vccd1 vccd1 _17594_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_91_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19333_ _19796_/CLK _19333_/D vssd1 vssd1 vccd1 vccd1 _19333_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__10618__C1 _09450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545_ _19495_/Q _16541_/C _16544_/Y vssd1 vssd1 vccd1 vccd1 _19495_/D sky130_fd_sc_hd__o21a_1
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13757_ _13757_/A vssd1 vssd1 vccd1 vccd1 _18445_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10969_ _10969_/A vssd1 vssd1 vccd1 vccd1 _10969_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ _19576_/Q _12701_/X _12706_/X _12707_/X vssd1 vssd1 vccd1 vccd1 _12708_/X
+ sky130_fd_sc_hd__a211o_1
X_19264_ _19264_/CLK _19264_/D vssd1 vssd1 vccd1 vccd1 _19264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_149_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16476_ _16485_/A _16476_/B _16476_/C vssd1 vssd1 vccd1 vccd1 _19476_/D sky130_fd_sc_hd__nor3_1
X_13688_ _13367_/X _18415_/Q _13690_/S vssd1 vssd1 vccd1 vccd1 _13689_/A sky130_fd_sc_hd__mux2_1
X_18215_ _18233_/A vssd1 vssd1 vccd1 vccd1 _18224_/A sky130_fd_sc_hd__clkbuf_1
X_15427_ _19120_/Q _15051_/X _15433_/S vssd1 vssd1 vccd1 vccd1 _15428_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13032__A0 _19718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12639_ _12639_/A vssd1 vssd1 vccd1 vccd1 _12895_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__11269__S0 _10969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19195_ _19391_/CLK _19195_/D vssd1 vssd1 vccd1 vccd1 _19195_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14862__A _14930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18146_ _18146_/A _18146_/B vssd1 vssd1 vccd1 vccd1 _18146_/X sky130_fd_sc_hd__or2_1
XFILLER_156_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15358_ _15358_/A vssd1 vssd1 vccd1 vccd1 _19089_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15169__S _15171_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14309_ _14309_/A vssd1 vssd1 vccd1 vccd1 _18649_/D sky130_fd_sc_hd__clkbuf_1
X_18077_ _18077_/A _18087_/B vssd1 vssd1 vccd1 vccd1 _18077_/X sky130_fd_sc_hd__or2_1
XFILLER_172_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15289_ _14582_/X _19059_/Q _15289_/S vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__mux2_1
XFILLER_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12138__A2 _12467_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17028_ _17028_/A _17133_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17085_/A sky130_fd_sc_hd__and3_2
XFILLER_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09850_ _09850_/A vssd1 vssd1 vccd1 vccd1 _10500_/S sky130_fd_sc_hd__buf_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11897__A1 _10749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _10217_/S vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__buf_2
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _19012_/CLK _18979_/D vssd1 vssd1 vccd1 vccd1 _18979_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11445__B _12465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17785__B1 _17784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15632__S _15632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10609__C1 _09450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12557__A _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clock clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 _19161_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_167_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09215_ _19856_/Q vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__buf_2
XFILLER_50_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13023__B1 _13022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14772__A _14772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__A _19734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__A _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09146_ _18146_/A _11528_/A _09146_/C _11560_/A vssd1 vssd1 vccd1 vccd1 _11530_/A
+ sky130_fd_sc_hd__or4_2
XANTENNA__10388__A1 _10297_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09873__S0 _09931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12292__A _19417_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13326__A1 _13325_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_163_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11337__B1 _09484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15807__S _15815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17294__S _17294_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14711__S _14713_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09979_ _09993_/A _09979_/B vssd1 vssd1 vccd1 vccd1 _09979_/X sky130_fd_sc_hd__or2_1
XFILLER_130_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12837__B1 _12704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_190_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12990_ _19529_/Q _13004_/A _12953_/A _19497_/Q _12989_/X vssd1 vssd1 vccd1 vccd1
+ _12990_/X sky130_fd_sc_hd__a221o_1
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _11969_/B _11793_/X _11936_/X _11940_/Y vssd1 vssd1 vccd1 vccd1 _16266_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14660_/A vssd1 vssd1 vccd1 vccd1 _18790_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11872_ _11873_/A _17195_/A vssd1 vssd1 vccd1 vccd1 _11872_/X sky130_fd_sc_hd__and2_1
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _15095_/A vssd1 vssd1 vccd1 vccd1 _13611_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10823_ _10823_/A _10823_/B vssd1 vssd1 vccd1 vccd1 _10823_/X sky130_fd_sc_hd__or2_1
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14591_ _14591_/A vssd1 vssd1 vccd1 vccd1 _18768_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14158__S _14158_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16330_ _16331_/B _16331_/C _19427_/Q vssd1 vssd1 vccd1 vccd1 _16332_/B sky130_fd_sc_hd__a21oi_1
XFILLER_125_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11812__A1 _11826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13542_ _18361_/Q _13541_/X _13545_/S vssd1 vssd1 vccd1 vccd1 _13543_/A sky130_fd_sc_hd__mux2_1
X_10754_ _19307_/Q _18719_/Q _18756_/Q _18330_/Q _10650_/X _11298_/A vssd1 vssd1 vccd1
+ vccd1 _10755_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16261_ _16261_/A vssd1 vssd1 vccd1 vccd1 _19400_/D sky130_fd_sc_hd__clkbuf_1
X_13473_ _13107_/X _18336_/Q _13481_/S vssd1 vssd1 vccd1 vccd1 _13474_/A sky130_fd_sc_hd__mux2_1
X_10685_ _19309_/Q _18721_/Q _18758_/Q _18332_/Q _10022_/X _10567_/X vssd1 vssd1 vccd1
+ vccd1 _10685_/X sky130_fd_sc_hd__mux4_1
XFILLER_9_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18000_ _18000_/A vssd1 vssd1 vccd1 vccd1 _19772_/D sky130_fd_sc_hd__clkbuf_1
X_15212_ _15212_/A vssd1 vssd1 vccd1 vccd1 _19024_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_172_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19365_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_138_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09776__A _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ _17917_/B _17232_/A vssd1 vssd1 vccd1 vccd1 _17920_/A sky130_fd_sc_hd__nand2_1
X_16192_ _16192_/A vssd1 vssd1 vccd1 vccd1 _19369_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09864__S0 _09846_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15143_ _18994_/Q _15057_/X _15145_/S vssd1 vssd1 vccd1 vccd1 _15144_/A sky130_fd_sc_hd__mux2_1
X_12355_ _17312_/A _17878_/A _12332_/B vssd1 vssd1 vccd1 vccd1 _12356_/B sky130_fd_sc_hd__a21boi_1
XFILLER_154_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10474__S1 _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11306_ _09982_/A _11303_/X _11305_/X _09989_/A vssd1 vssd1 vccd1 vccd1 _11307_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_153_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15074_ _18967_/Q _15073_/X _15077_/S vssd1 vssd1 vccd1 vccd1 _15075_/A sky130_fd_sc_hd__mux2_1
XFILLER_99_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12286_ _12286_/A vssd1 vssd1 vccd1 vccd1 _17856_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_142_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11328__B1 _09484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_187_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19307_/CLK sky130_fd_sc_hd__clkbuf_16
X_18902_ _18902_/CLK _18902_/D vssd1 vssd1 vccd1 vccd1 _18902_/Q sky130_fd_sc_hd__dfxtp_1
X_14025_ _14025_/A vssd1 vssd1 vccd1 vccd1 _18536_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15717__S _15721_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11237_ _09476_/A _11226_/X _11235_/X _09576_/A _11236_/Y vssd1 vssd1 vccd1 vccd1
+ _11238_/A sky130_fd_sc_hd__o32a_1
XANTENNA__14621__S _14621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16402__A _16546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10000__B1 _09737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18833_ _19315_/CLK _18833_/D vssd1 vssd1 vccd1 vccd1 _18833_/Q sky130_fd_sc_hd__dfxtp_1
X_11168_ _19710_/Q vssd1 vssd1 vccd1 vccd1 _11168_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_110_clock _19586_/CLK vssd1 vssd1 vccd1 vccd1 _19834_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__11546__A _14272_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10119_ _18408_/Q _18669_/Q _18568_/Q _18903_/Q _09786_/A _10169_/A vssd1 vssd1 vccd1
+ vccd1 _10120_/B sky130_fd_sc_hd__mux4_1
XANTENNA__18008__A1 _19397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18764_ _19315_/CLK _18764_/D vssd1 vssd1 vccd1 vccd1 _18764_/Q sky130_fd_sc_hd__dfxtp_1
X_15976_ _15976_/A vssd1 vssd1 vccd1 vccd1 _19319_/D sky130_fd_sc_hd__clkbuf_1
X_11099_ _18611_/Q _18946_/Q _11265_/S vssd1 vssd1 vccd1 vccd1 _11100_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09919__S1 _09905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17715_ _17715_/A vssd1 vssd1 vccd1 vccd1 _17715_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_36_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14927_ _14927_/A vssd1 vssd1 vccd1 vccd1 _18909_/D sky130_fd_sc_hd__clkbuf_1
X_18695_ _19377_/CLK _18695_/D vssd1 vssd1 vccd1 vccd1 _18695_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17646_ _17646_/A vssd1 vssd1 vccd1 vccd1 _17646_/X sky130_fd_sc_hd__clkbuf_2
X_14858_ _18879_/Q _14048_/X _14858_/S vssd1 vssd1 vccd1 vccd1 _14859_/A sky130_fd_sc_hd__mux2_1
XFILLER_51_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_125_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19423_/CLK sky130_fd_sc_hd__clkbuf_16
X_13809_ _13171_/X _18468_/Q _13809_/S vssd1 vssd1 vccd1 vccd1 _13810_/A sky130_fd_sc_hd__mux2_1
XFILLER_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14068__S _14074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17577_ _17730_/A _17576_/X _17577_/S vssd1 vssd1 vccd1 vccd1 _17577_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16990__A1 _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14789_ _14845_/A vssd1 vssd1 vccd1 vccd1 _14858_/S sky130_fd_sc_hd__buf_6
XFILLER_44_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19316_ _19378_/CLK _19316_/D vssd1 vssd1 vccd1 vccd1 _19316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16528_ _16529_/B _16529_/C _19491_/Q vssd1 vssd1 vccd1 vccd1 _16530_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12096__B _19399_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19247_ _19247_/CLK _19247_/D vssd1 vssd1 vccd1 vccd1 _19247_/Q sky130_fd_sc_hd__dfxtp_1
X_16459_ _16458_/A _16458_/C _19470_/Q vssd1 vssd1 vccd1 vccd1 _16460_/C sky130_fd_sc_hd__a21oi_1
XFILLER_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19178_ _19306_/CLK _19178_/D vssd1 vssd1 vccd1 vccd1 _19178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_145_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09855__S0 _09854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18129_ _12494_/A _18120_/X _18128_/Y _18123_/X vssd1 vssd1 vccd1 vccd1 _19826_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10465__S1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13308__A1 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09607__S0 _09599_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _10345_/A vssd1 vssd1 vccd1 vccd1 _10205_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__18247__A1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18247__B2 _18146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09932__B1 _10195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09833_ _09833_/A vssd1 vssd1 vccd1 vccd1 _09834_/A sky130_fd_sc_hd__clkbuf_2
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12819__B1 _12784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _09764_/A vssd1 vssd1 vccd1 vccd1 _09765_/A sky130_fd_sc_hd__buf_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15481__B2 _18255_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12295__A1 _12291_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ _09866_/A vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__A1 _09194_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16733__A1 _16736_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_137_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09596__A _09596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10470_ _18465_/Q _19056_/Q _19218_/Q _18433_/Q _10260_/A _10521_/A vssd1 vssd1 vccd1
+ vccd1 _10471_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ _19702_/Q _09305_/B vssd1 vssd1 vccd1 vccd1 _09235_/B sky130_fd_sc_hd__or2_1
XANTENNA__10456__S1 _09672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10535__A _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12140_ _12140_/A _12140_/B _17779_/A _12140_/D vssd1 vssd1 vccd1 vccd1 _12141_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_135_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10781__A1 _10639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__18238__A1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ _15632_/S vssd1 vssd1 vccd1 vccd1 _12071_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__10208__S1 _09905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18238__B2 _18140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14441__S _14443_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_132_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11022_ _11022_/A vssd1 vssd1 vccd1 vccd1 _11022_/X sky130_fd_sc_hd__buf_2
XFILLER_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10533__A1 _10535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15830_ _15830_/A vssd1 vssd1 vccd1 vccd1 _19254_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10270__A _10270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ _13586_/X _19224_/Q _15765_/S vssd1 vssd1 vccd1 vccd1 _15762_/A sky130_fd_sc_hd__mux2_1
XFILLER_66_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12973_ _13153_/A _12968_/X _12972_/X vssd1 vssd1 vccd1 vccd1 _12973_/X sky130_fd_sc_hd__a21bo_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_42_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19314_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_100_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15272__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17500_ _17613_/B _17499_/Y _17500_/S vssd1 vssd1 vccd1 vccd1 _17500_/X sky130_fd_sc_hd__mux2_1
XFILLER_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14712_/A vssd1 vssd1 vccd1 vccd1 _18814_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11924_ _19782_/Q vssd1 vssd1 vccd1 vccd1 _11924_/Y sky130_fd_sc_hd__inv_2
X_18480_ _19297_/CLK _18480_/D vssd1 vssd1 vccd1 vccd1 _18480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15692_ _15692_/A vssd1 vssd1 vccd1 vccd1 _19193_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16421__B1 _16402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _17425_/X _17428_/Y _09315_/B _17430_/X vssd1 vssd1 vccd1 vccd1 _19708_/D
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14643_ _15245_/B _15782_/B vssd1 vssd1 vccd1 vccd1 _14700_/A sky130_fd_sc_hd__nand2_4
XANTENNA__13235__A0 _19730_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11855_ _11855_/A vssd1 vssd1 vccd1 vccd1 _11855_/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__16892__A _16915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16972__A1 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output105_A _17174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17362_ _17265_/X _17260_/X _17372_/S vssd1 vssd1 vccd1 vccd1 _17362_/X sky130_fd_sc_hd__mux2_1
X_10806_ _11257_/A vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__buf_2
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19027_/CLK sky130_fd_sc_hd__clkbuf_16
X_14574_ _14573_/X _18763_/Q _14583_/S vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10144__S0 _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11786_ _19777_/Q _11288_/A _11925_/S vssd1 vssd1 vccd1 vccd1 _17247_/A sky130_fd_sc_hd__mux2_8
X_19101_ _19292_/CLK _19101_/D vssd1 vssd1 vccd1 vccd1 _19101_/Q sky130_fd_sc_hd__dfxtp_1
X_16313_ _19469_/Q _19471_/Q _19470_/Q _16453_/A vssd1 vssd1 vccd1 vccd1 _16461_/A
+ sky130_fd_sc_hd__and4_1
X_13525_ _15009_/A vssd1 vssd1 vccd1 vccd1 _13525_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_158_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17293_ _12405_/A _17410_/B _17293_/S vssd1 vssd1 vccd1 vccd1 _17293_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10737_ _09995_/A _10728_/X _10732_/X _10736_/X _11307_/A vssd1 vssd1 vccd1 vccd1
+ _10737_/X sky130_fd_sc_hd__a311o_2
XFILLER_13_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10695__S1 _10577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13520__S _13529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19032_ _19384_/CLK _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/Q sky130_fd_sc_hd__dfxtp_1
X_16244_ _16244_/A vssd1 vssd1 vccd1 vccd1 _19393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13456_ _13456_/A vssd1 vssd1 vccd1 vccd1 _18328_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_51_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10668_ _18620_/Q _18955_/Q _11299_/S vssd1 vssd1 vccd1 vccd1 _10669_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09206__A2 _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12407_ _12388_/A _12388_/B _12387_/A _12386_/A vssd1 vssd1 vccd1 vccd1 _12408_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_12_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16175_ _16175_/A vssd1 vssd1 vccd1 vccd1 _19361_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12210__A1 _11619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10445__A _19724_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _11452_/A vssd1 vssd1 vccd1 vccd1 _10599_/Y sky130_fd_sc_hd__inv_2
X_13387_ _13386_/X _18314_/Q _13387_/S vssd1 vssd1 vccd1 vccd1 _13388_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput107 _12482_/B vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[0] sky130_fd_sc_hd__buf_2
XFILLER_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15126_ _18986_/Q _15031_/X _15134_/S vssd1 vssd1 vccd1 vccd1 _15127_/A sky130_fd_sc_hd__mux2_1
Xoutput118 _12466_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[18] sky130_fd_sc_hd__buf_2
Xoutput129 _12478_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[28] sky130_fd_sc_hd__buf_2
X_12338_ _19418_/Q _12339_/C _19419_/Q vssd1 vssd1 vccd1 vccd1 _12340_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10772__B2 _19716_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15447__S _15455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15057_ _15057_/A vssd1 vssd1 vccd1 vccd1 _15057_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12269_ _12269_/A vssd1 vssd1 vccd1 vccd1 _12269_/Y sky130_fd_sc_hd__inv_2
X_14008_ _18531_/Q _14007_/X _14011_/S vssd1 vssd1 vccd1 vccd1 _14009_/A sky130_fd_sc_hd__mux2_1
XFILLER_141_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19865_ _19865_/CLK _19865_/D vssd1 vssd1 vccd1 vccd1 _19865_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11721__A0 _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18816_ _19235_/CLK _18816_/D vssd1 vssd1 vccd1 vccd1 _18816_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10180__A _10181_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19796_ _19796_/CLK _19796_/D vssd1 vssd1 vccd1 vccd1 _19796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15959_ _13560_/X _19312_/Q _15959_/S vssd1 vssd1 vccd1 vccd1 _15960_/A sky130_fd_sc_hd__mux2_1
X_18747_ _19202_/CLK _18747_/D vssd1 vssd1 vccd1 vccd1 _18747_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15182__S _15184_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09480_ _10914_/A vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__clkbuf_4
X_18678_ _19361_/CLK _18678_/D vssd1 vssd1 vccd1 vccd1 _18678_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15215__A1 _15057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17629_ _17627_/X _17628_/Y _17855_/S vssd1 vssd1 vccd1 vccd1 _17629_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_149_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14526__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13529__A1 _13528_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_117_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10355__A _11351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15357__S _15361_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13666__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13162__C1 _13161_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09816_ _19198_/Q _18812_/Q _19262_/Q _18381_/Q _09815_/X _09799_/X vssd1 vssd1 vccd1
+ vccd1 _09817_/B sky130_fd_sc_hd__mux4_1
XFILLER_74_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09747_ _11368_/A _09747_/B vssd1 vssd1 vccd1 vccd1 _09747_/X sky130_fd_sc_hd__or2_1
XFILLER_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09678_ _09733_/A vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16403__B1 _16402_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15820__S _15826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _12093_/A vssd1 vssd1 vccd1 vccd1 _11640_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__17601__A _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10964__S _10964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ _11672_/S _17168_/B vssd1 vssd1 vccd1 vccd1 _11571_/Y sky130_fd_sc_hd__nor2_1
XFILLER_22_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13310_ _15086_/A vssd1 vssd1 vccd1 vccd1 _14608_/A sky130_fd_sc_hd__clkbuf_1
X_10522_ _10348_/A _10519_/Y _10521_/Y _10277_/A vssd1 vssd1 vccd1 vccd1 _10522_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_168_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14290_ _14290_/A _18222_/B vssd1 vssd1 vccd1 vccd1 _14291_/A sky130_fd_sc_hd__and2_2
XFILLER_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12464__B _12464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10453_ _09674_/A _10450_/X _10452_/X vssd1 vssd1 vccd1 vccd1 _10453_/X sky130_fd_sc_hd__a21o_1
X_13241_ _13240_/X _18306_/Q _13252_/S vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__mux2_1
XFILLER_171_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10265__A _10378_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12743__A2 _12739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ _13171_/X _18302_/Q _13172_/S vssd1 vssd1 vccd1 vccd1 _13173_/A sky130_fd_sc_hd__mux2_1
X_10384_ _18403_/Q _18664_/Q _18563_/Q _18898_/Q _10274_/X _10263_/X vssd1 vssd1 vccd1
+ vccd1 _10384_/X sky130_fd_sc_hd__mux4_1
XANTENNA_input66_A io_ibus_valid vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13576__A _15060_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ _12123_/A vssd1 vssd1 vccd1 vccd1 _12123_/Y sky130_fd_sc_hd__clkinv_2
X_17980_ _17980_/A vssd1 vssd1 vccd1 vccd1 _19763_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16931_ _16931_/A _16937_/C _17149_/A vssd1 vssd1 vccd1 vccd1 _16931_/X sky130_fd_sc_hd__and3_1
X_12054_ _17756_/B _12054_/B vssd1 vssd1 vccd1 vccd1 _12056_/A sky130_fd_sc_hd__xnor2_2
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11005_ _11012_/A vssd1 vssd1 vccd1 vccd1 _11005_/X sky130_fd_sc_hd__clkbuf_4
X_19650_ _19687_/CLK _19650_/D vssd1 vssd1 vccd1 vccd1 _19650_/Q sky130_fd_sc_hd__dfxtp_1
X_16862_ _19599_/Q _16862_/B _16862_/C vssd1 vssd1 vccd1 vccd1 _16864_/B sky130_fd_sc_hd__and3_1
XFILLER_120_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18601_ _19096_/CLK _18601_/D vssd1 vssd1 vccd1 vccd1 _18601_/Q sky130_fd_sc_hd__dfxtp_1
X_15813_ _13557_/X _19247_/Q _15815_/S vssd1 vssd1 vccd1 vccd1 _15814_/A sky130_fd_sc_hd__mux2_1
X_19581_ _19581_/CLK _19581_/D vssd1 vssd1 vccd1 vccd1 _19581_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12259__A1 _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16793_ _19571_/Q _16791_/B _16792_/Y vssd1 vssd1 vccd1 vccd1 _19571_/D sky130_fd_sc_hd__o21a_1
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18532_ _19285_/CLK _18532_/D vssd1 vssd1 vccd1 vccd1 _18532_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15744_ _15744_/A vssd1 vssd1 vccd1 vccd1 _19216_/D sky130_fd_sc_hd__clkbuf_1
X_12956_ _12956_/A _12956_/B vssd1 vssd1 vccd1 vccd1 _12956_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14200__A _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10365__S0 _10315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18463_ _19248_/CLK _18463_/D vssd1 vssd1 vccd1 vccd1 _18463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_73_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11907_ _11915_/A _11969_/D vssd1 vssd1 vccd1 vccd1 _11908_/B sky130_fd_sc_hd__or2_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15675_ _15675_/A vssd1 vssd1 vccd1 vccd1 _19185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16945__A1 _13410_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _12886_/X _18287_/Q _12887_/S vssd1 vssd1 vccd1 vccd1 _12888_/A sky130_fd_sc_hd__mux2_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17406_/X _17418_/B _17411_/X _17413_/X vssd1 vssd1 vccd1 vccd1 _17414_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14626_ _14626_/A vssd1 vssd1 vccd1 vccd1 _18779_/D sky130_fd_sc_hd__clkbuf_1
X_18394_ _19308_/CLK _18394_/D vssd1 vssd1 vccd1 vccd1 _18394_/Q sky130_fd_sc_hd__dfxtp_1
X_11838_ _11890_/B _12453_/A _11890_/C _19863_/Q vssd1 vssd1 vccd1 vccd1 _11893_/A
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17291_/S _17238_/X _17344_/X vssd1 vssd1 vccd1 vccd1 _17345_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14557_ _14557_/A vssd1 vssd1 vccd1 vccd1 _14557_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14346__S _14354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09832__C1 _09831_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _11769_/A vssd1 vssd1 vccd1 vccd1 _12098_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_147_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15031__A _15031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13508_ _13508_/A vssd1 vssd1 vccd1 vccd1 _18352_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_147_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17276_ _17802_/B _17680_/B _17283_/S vssd1 vssd1 vccd1 vccd1 _17276_/X sky130_fd_sc_hd__mux2_1
X_14488_ _14488_/A vssd1 vssd1 vccd1 vccd1 _18728_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_146_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19015_ _19329_/CLK _19015_/D vssd1 vssd1 vccd1 vccd1 _19015_/Q sky130_fd_sc_hd__dfxtp_1
X_16227_ _13595_/X _19385_/Q _16235_/S vssd1 vssd1 vccd1 vccd1 _16228_/A sky130_fd_sc_hd__mux2_1
X_13439_ _13507_/S vssd1 vssd1 vccd1 vccd1 _13448_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09964__A _09964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16158_ _16158_/A vssd1 vssd1 vccd1 vccd1 _19357_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_138_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _15109_/A vssd1 vssd1 vccd1 vccd1 _18978_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14081__S _14085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16089_ _16087_/X _19345_/Q _16112_/S vssd1 vssd1 vccd1 vccd1 _16090_/A sky130_fd_sc_hd__mux2_1
XFILLER_130_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15905__S _15909_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10114__S _10114_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19848_ _19865_/CLK _19848_/D vssd1 vssd1 vccd1 vccd1 _19848_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09601_ _18607_/Q _18878_/Q _19102_/Q _18846_/Q _09599_/X _09977_/A vssd1 vssd1 vccd1
+ vccd1 _09601_/X sky130_fd_sc_hd__mux4_1
XFILLER_95_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19779_ _19779_/CLK _19779_/D vssd1 vssd1 vccd1 vccd1 _19779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ _11164_/A vssd1 vssd1 vccd1 vccd1 _10839_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10356__S0 _10315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09463_ _18783_/Q vssd1 vssd1 vccd1 vccd1 _09464_/A sky130_fd_sc_hd__inv_2
XFILLER_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12670__B2 _12696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09394_ _09394_/A vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__buf_2
XFILLER_52_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10028__A3 _10026_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14256__S _14264_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09874__A _10197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15087__S _15093_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_105_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15815__S _15815_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12810_ _14715_/C _15173_/A _13947_/B vssd1 vssd1 vccd1 vccd1 _13275_/A sky130_fd_sc_hd__or3_4
X_13790_ _13025_/X _18459_/Q _13798_/S vssd1 vssd1 vccd1 vccd1 _13791_/A sky130_fd_sc_hd__mux2_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09114__A _18083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ hold19/A _12739_/X _11016_/X _12740_/X vssd1 vssd1 vccd1 vccd1 _18256_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12661__B2 _19340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15460_ _15460_/A vssd1 vssd1 vccd1 vccd1 _19135_/D sky130_fd_sc_hd__clkbuf_1
X_12672_ _12672_/A vssd1 vssd1 vccd1 vccd1 _13392_/A sky130_fd_sc_hd__inv_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411_ _13893_/X _18694_/Q _14417_/S vssd1 vssd1 vccd1 vccd1 _14412_/A sky130_fd_sc_hd__mux2_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__clkbuf_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12413__A1 _19358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15391_ _15459_/S vssd1 vssd1 vccd1 vccd1 _15400_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__C1 _09813_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17130_ _17130_/A _17130_/B _17130_/C _17130_/D vssd1 vssd1 vccd1 vccd1 _17131_/D
+ sky130_fd_sc_hd__or4_1
X_14342_ _14342_/A vssd1 vssd1 vccd1 vccd1 _18664_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_129_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11554_ _12134_/A _11553_/Y _19392_/Q vssd1 vssd1 vccd1 vccd1 _16241_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09290__B1 _12548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12194__B _12195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17061_ _19678_/Q _15542_/X _17061_/S vssd1 vssd1 vccd1 vccd1 _17062_/A sky130_fd_sc_hd__mux2_1
X_10505_ _10514_/A _10505_/B vssd1 vssd1 vccd1 vccd1 _10505_/X sky130_fd_sc_hd__or2_1
XFILLER_10_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14273_ _14627_/A vssd1 vssd1 vccd1 vccd1 _18197_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_156_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11485_ _17120_/A _17183_/A vssd1 vssd1 vccd1 vccd1 _11485_/X sky130_fd_sc_hd__and2_1
XFILLER_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16012_ _16011_/A _16011_/C _16011_/B vssd1 vssd1 vccd1 vccd1 _16013_/B sky130_fd_sc_hd__o21ai_1
XFILLER_171_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13224_ _13154_/X _13223_/X _13164_/X vssd1 vssd1 vccd1 vccd1 _13224_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_137_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10436_ _10436_/A _10436_/B vssd1 vssd1 vccd1 vccd1 _10436_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17104__B2 _11557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15115__A0 _18981_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_128_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13155_ _19607_/Q vssd1 vssd1 vccd1 vccd1 _16887_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10367_ _18627_/Q _18962_/Q _10367_/S vssd1 vssd1 vccd1 vccd1 _10367_/X sky130_fd_sc_hd__mux2_1
XFILLER_124_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10822__S1 _10802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _11884_/X _12104_/Y _12156_/C _11835_/X vssd1 vssd1 vccd1 vccd1 _12106_/Y
+ sky130_fd_sc_hd__o31ai_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10378_/A _10295_/X _10297_/X vssd1 vssd1 vccd1 vccd1 _10298_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _13111_/C _13086_/B vssd1 vssd1 vccd1 vccd1 _13086_/Y sky130_fd_sc_hd__nor2_1
X_17963_ _17963_/A vssd1 vssd1 vccd1 vccd1 _19755_/D sky130_fd_sc_hd__clkbuf_1
X_19702_ _19706_/CLK _19702_/D vssd1 vssd1 vccd1 vccd1 _19702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16914_ _16914_/A _16914_/B _16914_/C vssd1 vssd1 vccd1 vccd1 _19617_/D sky130_fd_sc_hd__nor3_1
X_12037_ _12037_/A vssd1 vssd1 vccd1 vccd1 _12037_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11152__A1 _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17894_ _12369_/B _17786_/X _17893_/X _17795_/X vssd1 vssd1 vccd1 vccd1 _17894_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19633_ _19669_/CLK _19633_/D vssd1 vssd1 vccd1 vccd1 _19633_/Q sky130_fd_sc_hd__dfxtp_2
X_16845_ _19593_/Q _16845_/B _16845_/C vssd1 vssd1 vccd1 vccd1 _16847_/B sky130_fd_sc_hd__and3_1
XANTENNA__18080__A2 _12739_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19564_ _19564_/CLK _19564_/D vssd1 vssd1 vccd1 vccd1 _19564_/Q sky130_fd_sc_hd__dfxtp_1
X_16776_ _16782_/C _16782_/D _16775_/Y vssd1 vssd1 vccd1 vccd1 _19566_/D sky130_fd_sc_hd__o21a_1
X_13988_ _14560_/A vssd1 vssd1 vccd1 vccd1 _13988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_92_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12369__B _12369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18515_ _19074_/CLK _18515_/D vssd1 vssd1 vccd1 vccd1 _18515_/Q sky130_fd_sc_hd__dfxtp_1
X_15727_ _15727_/A vssd1 vssd1 vccd1 vccd1 _19208_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_46_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12939_ _12938_/X _19527_/Q _12939_/S vssd1 vssd1 vccd1 vccd1 _12939_/X sky130_fd_sc_hd__mux2_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10258__A3 _10257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19495_ _19619_/CLK _19495_/D vssd1 vssd1 vccd1 vccd1 _19495_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15658_ _14547_/X _19178_/Q _15660_/S vssd1 vssd1 vccd1 vccd1 _15659_/A sky130_fd_sc_hd__mux2_1
X_18446_ _19261_/CLK _18446_/D vssd1 vssd1 vccd1 vccd1 _18446_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17125__C_N _18125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14609_ _14608_/X _18774_/Q _14615_/S vssd1 vssd1 vccd1 vccd1 _14610_/A sky130_fd_sc_hd__mux2_1
X_18377_ _19610_/CLK _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12404__A1 _11413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15589_ _19729_/Q _15588_/X _15595_/S vssd1 vssd1 vccd1 vccd1 _15589_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_147_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17328_ _17328_/A _17328_/B _17328_/C vssd1 vssd1 vccd1 vccd1 _17328_/X sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_11_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10966__A1 _10965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17259_ _17229_/X _17257_/X _17504_/S vssd1 vssd1 vccd1 vccd1 _17740_/A sky130_fd_sc_hd__mux2_1
XFILLER_128_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_162_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09515_ _10623_/A vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__buf_2
XFILLER_25_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15370__S _15372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09869__A _09931_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ _18782_/Q vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__buf_2
XFILLER_80_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ _10990_/A vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__buf_4
XFILLER_40_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_153_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13838__B _14297_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ _11024_/A _11269_/X _10914_/A vssd1 vssd1 vccd1 vccd1 _11270_/X sky130_fd_sc_hd__o21a_1
XFILLER_134_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10221_ _18406_/Q _18667_/Q _18566_/Q _18901_/Q _09952_/S _09891_/A vssd1 vssd1 vccd1
+ vccd1 _10221_/X sky130_fd_sc_hd__mux4_1
XANTENNA__11639__A _11639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10152_ _19288_/Q _19126_/Q _18535_/Q _18305_/Q _09931_/S _09871_/A vssd1 vssd1 vccd1
+ vccd1 _10153_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14960_ _18926_/Q vssd1 vssd1 vccd1 vccd1 _14961_/A sky130_fd_sc_hd__clkbuf_1
X_10083_ _11426_/A _10083_/B _10082_/X vssd1 vssd1 vccd1 vccd1 _11360_/B sky130_fd_sc_hd__or3b_1
XFILLER_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA__10568__S0 _10566_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13911_ _13911_/A vssd1 vssd1 vccd1 vccd1 _18502_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_102_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12882__A1 _15479_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input29_A io_dbus_rdata[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _18893_/Q _13991_/X _14893_/S vssd1 vssd1 vccd1 vccd1 _14892_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17270__A0 _12245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16630_ _19520_/Q _16634_/B _19521_/Q vssd1 vssd1 vccd1 vccd1 _16633_/B sky130_fd_sc_hd__a21oi_1
XFILLER_114_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13842_ _13941_/S vssd1 vssd1 vccd1 vccd1 _13855_/S sky130_fd_sc_hd__buf_2
XFILLER_75_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16561_ _19501_/Q _16561_/B vssd1 vssd1 vccd1 vccd1 _16567_/C sky130_fd_sc_hd__and2_1
XFILLER_90_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13773_ _13773_/A vssd1 vssd1 vccd1 vccd1 _18451_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_128_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ _19713_/Q vssd1 vssd1 vccd1 vccd1 _10985_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18300_ _19377_/CLK _18300_/D vssd1 vssd1 vccd1 vccd1 _18300_/Q sky130_fd_sc_hd__dfxtp_1
X_15512_ _15512_/A vssd1 vssd1 vccd1 vccd1 _19146_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09779__A _10381_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19280_ _19280_/CLK _19280_/D vssd1 vssd1 vccd1 vccd1 _19280_/Q sky130_fd_sc_hd__dfxtp_1
X_12724_ _09194_/X _11239_/A _12735_/S vssd1 vssd1 vccd1 vccd1 _12724_/X sky130_fd_sc_hd__mux2_1
X_16492_ _16549_/A vssd1 vssd1 vccd1 vccd1 _16541_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10740__S0 _10660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18231_ _18231_/A _18231_/B vssd1 vssd1 vccd1 vccd1 _18232_/A sky130_fd_sc_hd__and2_1
X_15443_ _15443_/A vssd1 vssd1 vccd1 vccd1 _19127_/D sky130_fd_sc_hd__clkbuf_1
X_12655_ _16929_/B _12651_/X _12653_/X _17102_/B _19584_/Q vssd1 vssd1 vccd1 vccd1
+ _12655_/X sky130_fd_sc_hd__o32a_1
XANTENNA__17996__A _18029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16781__C1 _16293_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_169_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18162_ _09172_/C _12674_/A _18148_/Y input60/X vssd1 vssd1 vccd1 vccd1 _18163_/B
+ sky130_fd_sc_hd__o22a_1
X_11606_ _11607_/A _11607_/B _17230_/A vssd1 vssd1 vccd1 vccd1 _11606_/X sky130_fd_sc_hd__o21a_1
X_15374_ _15374_/A vssd1 vssd1 vccd1 vccd1 _15383_/S sky130_fd_sc_hd__buf_4
X_12586_ _19506_/Q _12586_/B vssd1 vssd1 vccd1 vccd1 _12586_/X sky130_fd_sc_hd__and2_1
XFILLER_129_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_185_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ _17120_/A vssd1 vssd1 vccd1 vccd1 _17114_/A sky130_fd_sc_hd__buf_2
X_14325_ _14325_/A vssd1 vssd1 vccd1 vccd1 _18656_/D sky130_fd_sc_hd__clkbuf_1
X_18093_ _18121_/A vssd1 vssd1 vccd1 vccd1 _18116_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ _18744_/Q vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_172_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15887__A1 _14566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17044_ _19670_/Q _15495_/X _17050_/S vssd1 vssd1 vccd1 vccd1 _17045_/A sky130_fd_sc_hd__mux2_1
X_14256_ _18634_/Q _14029_/X _14264_/S vssd1 vssd1 vccd1 vccd1 _14257_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output97_A _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _11468_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11468_/X sky130_fd_sc_hd__and2_1
XFILLER_48_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ _13197_/X _13205_/Y _13206_/Y vssd1 vssd1 vccd1 vccd1 _15067_/A sky130_fd_sc_hd__a21oi_4
X_10419_ _10419_/A _10419_/B vssd1 vssd1 vccd1 vccd1 _10419_/X sky130_fd_sc_hd__or2_1
XFILLER_48_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14187_ _18604_/Q _14036_/X _14191_/S vssd1 vssd1 vccd1 vccd1 _14188_/A sky130_fd_sc_hd__mux2_1
X_11399_ _19297_/Q _19135_/Q _18544_/Q _18314_/Q _09815_/X _09799_/X vssd1 vssd1 vccd1
+ vccd1 _11400_/B sky130_fd_sc_hd__mux4_1
XFILLER_152_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _14576_/A vssd1 vssd1 vccd1 vccd1 _13138_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _19089_/CLK _18995_/D vssd1 vssd1 vccd1 vccd1 _18995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15455__S _15455_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16778__C _16778_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _15041_/A vssd1 vssd1 vccd1 vccd1 _14563_/A sky130_fd_sc_hd__clkbuf_2
X_17946_ _12994_/A _19780_/Q _17946_/S vssd1 vssd1 vccd1 vccd1 _17947_/A sky130_fd_sc_hd__mux2_1
XFILLER_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_94_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17877_ _17875_/X _17876_/Y _17898_/S vssd1 vssd1 vccd1 vccd1 _17877_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17261__A0 _12089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09238__C_N _09172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__A _11284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19616_ _19618_/CLK _19616_/D vssd1 vssd1 vccd1 vccd1 _19616_/Q sky130_fd_sc_hd__dfxtp_1
X_16828_ _18136_/A _16828_/B _16830_/B vssd1 vssd1 vccd1 vccd1 _16829_/A sky130_fd_sc_hd__and3_1
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19547_ _19549_/CLK _19547_/D vssd1 vssd1 vccd1 vccd1 _19547_/Q sky130_fd_sc_hd__dfxtp_1
X_16759_ _16799_/A _16759_/B _16767_/C vssd1 vssd1 vccd1 vccd1 _19561_/D sky130_fd_sc_hd__nor3_1
XFILLER_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09300_ _16623_/A _16623_/B _16937_/C _09299_/X vssd1 vssd1 vccd1 vccd1 _09301_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13703__S _13703_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19478_ _19610_/CLK _19478_/D vssd1 vssd1 vccd1 vccd1 _19478_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09231_ _09207_/X _11942_/A _09230_/X vssd1 vssd1 vccd1 vccd1 _09231_/X sky130_fd_sc_hd__o21a_1
XFILLER_22_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18429_ _19248_/CLK _18429_/D vssd1 vssd1 vccd1 vccd1 _18429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09201__B _19814_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09162_ _09182_/C _09182_/B _09113_/A vssd1 vssd1 vccd1 vccd1 _11528_/C sky130_fd_sc_hd__nor3b_1
XFILLER_148_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ _19848_/Q vssd1 vssd1 vccd1 vccd1 _09174_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_119_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_163_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_131_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09995_ _09995_/A vssd1 vssd1 vccd1 vccd1 _09995_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__10082__B _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_131_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12616__A1 _13397_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16196__S _16202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14709__S _14709_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09599__A _10654_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _09597_/X _10767_/X _10769_/X _09602_/X vssd1 vssd1 vccd1 vccd1 _10770_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09429_ _18782_/Q vssd1 vssd1 vccd1 vccd1 _11007_/A sky130_fd_sc_hd__inv_2
XFILLER_158_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _12440_/A _12440_/B vssd1 vssd1 vccd1 vccd1 _12440_/Y sky130_fd_sc_hd__nand2_1
XFILLER_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12371_ _19420_/Q _12371_/B vssd1 vssd1 vccd1 vccd1 _12410_/C sky130_fd_sc_hd__and2_1
XANTENNA__11572__A1_N _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14110_ _13921_/X _18570_/Q _14118_/S vssd1 vssd1 vccd1 vccd1 _14111_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11322_ _09651_/A _11319_/Y _11321_/Y _10575_/A vssd1 vssd1 vccd1 vccd1 _11322_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_4_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15090_ _18972_/Q _15089_/X _15093_/S vssd1 vssd1 vccd1 vccd1 _15091_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12472__B _12472_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14041_ _14041_/A vssd1 vssd1 vccd1 vccd1 _18541_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_106_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ _19298_/Q _18710_/Q _18747_/Q _18321_/Q _09410_/A _10801_/A vssd1 vssd1 vccd1
+ vccd1 _11254_/B sky130_fd_sc_hd__mux4_1
XFILLER_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09643__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16818__B1 _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _19191_/Q _18805_/Q _19255_/Q _18374_/Q _09955_/S _09954_/A vssd1 vssd1 vccd1
+ vccd1 _10205_/B sky130_fd_sc_hd__mux4_1
XFILLER_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11184_ _11184_/A _11184_/B vssd1 vssd1 vccd1 vccd1 _11184_/X sky130_fd_sc_hd__or2_1
XANTENNA__10563__C1 _09989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11519__D _18087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17800_ _17800_/A _17800_/B vssd1 vssd1 vccd1 vccd1 _17800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10135_ _11357_/A _12472_/B vssd1 vssd1 vccd1 vccd1 _11422_/A sky130_fd_sc_hd__or2_1
XFILLER_95_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18780_ _19711_/CLK _18780_/D vssd1 vssd1 vccd1 vccd1 _18780_/Q sky130_fd_sc_hd__dfxtp_4
X_15992_ _13608_/X _19327_/Q _15992_/S vssd1 vssd1 vccd1 vccd1 _15993_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17731_ _17730_/Y _17572_/X _17731_/S vssd1 vssd1 vccd1 vccd1 _17731_/X sky130_fd_sc_hd__mux2_1
X_14943_ _14943_/A vssd1 vssd1 vccd1 vccd1 _18917_/D sky130_fd_sc_hd__clkbuf_1
X_10066_ _19197_/Q _18811_/Q _19261_/Q _18380_/Q _09500_/A _10693_/A vssd1 vssd1 vccd1
+ vccd1 _10067_/B sky130_fd_sc_hd__mux4_1
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14057__A0 _13845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14874_ _18885_/Q _13965_/X _14882_/S vssd1 vssd1 vccd1 vccd1 _14875_/A sky130_fd_sc_hd__mux2_1
X_17662_ _17662_/A _17662_/B vssd1 vssd1 vccd1 vccd1 _17664_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19401_ _19838_/CLK _19401_/D vssd1 vssd1 vccd1 vccd1 _19401_/Q sky130_fd_sc_hd__dfxtp_4
X_16613_ _19518_/Q _16613_/B vssd1 vssd1 vccd1 vccd1 _16614_/B sky130_fd_sc_hd__and2_1
X_13825_ _13294_/X _18475_/Q _13831_/S vssd1 vssd1 vccd1 vccd1 _13826_/A sky130_fd_sc_hd__mux2_1
X_17593_ _17571_/X _17578_/X _17591_/X _17592_/X vssd1 vssd1 vccd1 vccd1 _17593_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_63_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13523__S _13529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16544_ _16570_/A _16551_/C vssd1 vssd1 vccd1 vccd1 _16544_/Y sky130_fd_sc_hd__nor2_1
X_19332_ _19802_/CLK _19332_/D vssd1 vssd1 vccd1 vccd1 _19332_/Q sky130_fd_sc_hd__dfxtp_2
X_13756_ _13330_/X _18445_/Q _13758_/S vssd1 vssd1 vccd1 vccd1 _13757_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10968_ _10968_/A vssd1 vssd1 vccd1 vccd1 _11085_/A sky130_fd_sc_hd__buf_2
XFILLER_44_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17546__A1 _11732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10713__S0 _09645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ _13265_/A vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_16475_ _16474_/A _16474_/C _19476_/Q vssd1 vssd1 vccd1 vccd1 _16476_/C sky130_fd_sc_hd__a21oi_1
X_19263_ _19389_/CLK _19263_/D vssd1 vssd1 vccd1 vccd1 _19263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ _13687_/A vssd1 vssd1 vccd1 vccd1 _18414_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_148_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ _18616_/Q _18951_/Q _10964_/S vssd1 vssd1 vccd1 vccd1 _10900_/B sky130_fd_sc_hd__mux2_1
X_15426_ _15426_/A vssd1 vssd1 vccd1 vccd1 _19119_/D sky130_fd_sc_hd__clkbuf_1
X_18214_ _18214_/A vssd1 vssd1 vccd1 vccd1 _19854_/D sky130_fd_sc_hd__clkbuf_1
X_12638_ _13055_/A vssd1 vssd1 vccd1 vccd1 _12638_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_19194_ _19610_/CLK _19194_/D vssd1 vssd1 vccd1 vccd1 _19194_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13032__A1 _12649_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11269__S1 _09511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18145_ _16623_/B _18134_/X _18144_/X _18136_/X vssd1 vssd1 vccd1 vccd1 _19833_/D
+ sky130_fd_sc_hd__o211a_1
X_15357_ _19089_/Q _15054_/X _15361_/S vssd1 vssd1 vccd1 vccd1 _15358_/A sky130_fd_sc_hd__mux2_1
X_12569_ _19622_/Q _12496_/C _12565_/X _19648_/Q _12568_/X vssd1 vssd1 vccd1 vccd1
+ _12569_/X sky130_fd_sc_hd__a221o_1
XANTENNA__14354__S _14354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14308_ _13851_/X _18649_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _14309_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18076_ _19805_/Q _12627_/X _18075_/X _17021_/X vssd1 vssd1 vccd1 vccd1 _19805_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_116_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15288_ _15288_/A vssd1 vssd1 vccd1 vccd1 _19058_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17027_ _17027_/A vssd1 vssd1 vccd1 vccd1 _19663_/D sky130_fd_sc_hd__clkbuf_1
X_14239_ _14239_/A vssd1 vssd1 vccd1 vccd1 _18626_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09972__A _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10554__C1 _09450_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13494__A _13494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ _10215_/S vssd1 vssd1 vccd1 vccd1 _10217_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _19012_/CLK _18978_/D vssd1 vssd1 vccd1 vccd1 _18978_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17929_ _19740_/Q _19772_/Q _17935_/S vssd1 vssd1 vccd1 vccd1 _17930_/A sky130_fd_sc_hd__mux2_1
XFILLER_67_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16037__A1 _19336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15796__A0 _13531_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14529__S _14535_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13271__A1 _12848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11282__B1 _09576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _17184_/C _17176_/A _17145_/A vssd1 vssd1 vccd1 vccd1 _11942_/A sky130_fd_sc_hd__or3b_4
XANTENNA__13023__A1 _11538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ _09182_/C _09182_/B _09113_/A vssd1 vssd1 vccd1 vccd1 _11560_/A sky130_fd_sc_hd__or3b_1
XANTENNA__14264__S _14264_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09873__S1 _09871_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_107_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_opt_1_0_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09978_ _18938_/Q _18704_/Q _19386_/Q _19034_/Q _10602_/S _09977_/X vssd1 vssd1 vccd1
+ vccd1 _09979_/B sky130_fd_sc_hd__mux4_1
XFILLER_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_133_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11636__B _17239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11128__S _11128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11940_ _12230_/A _11938_/Y _11994_/C _11962_/A vssd1 vssd1 vccd1 vccd1 _11940_/Y
+ sky130_fd_sc_hd__o31ai_1
XANTENNA__10032__S _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_73_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15787__A0 _13519_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _19780_/Q _10798_/A _11925_/S vssd1 vssd1 vccd1 vccd1 _17195_/A sky130_fd_sc_hd__mux2_4
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14439__S _14439_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _13610_/A vssd1 vssd1 vccd1 vccd1 _18382_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ _18920_/Q _18686_/Q _19368_/Q _19016_/Q _09598_/A _10802_/X vssd1 vssd1 vccd1
+ vccd1 _10823_/B sky130_fd_sc_hd__mux4_1
XFILLER_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14590_ _14589_/X _18768_/Q _14599_/S vssd1 vssd1 vccd1 vccd1 _14591_/A sky130_fd_sc_hd__mux2_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17528__A1 _17731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12467__B _12467_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13541_ _15025_/A vssd1 vssd1 vccd1 vccd1 _13541_/X sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_1_clock clkbuf_1_1_1_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_111_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10753_ _11309_/A _10753_/B vssd1 vssd1 vccd1 vccd1 _10753_/X sky130_fd_sc_hd__or2_1
XFILLER_13_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16260_ _16266_/A _16260_/B vssd1 vssd1 vccd1 vccd1 _16261_/A sky130_fd_sc_hd__or2_1
X_13472_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13481_/S sky130_fd_sc_hd__buf_4
X_10684_ _10684_/A _10684_/B vssd1 vssd1 vccd1 vccd1 _10684_/Y sky130_fd_sc_hd__nor2_1
X_15211_ _19024_/Q _15051_/X _15217_/S vssd1 vssd1 vccd1 vccd1 _15212_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13579__A _15063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _19802_/Q _12422_/Y _12423_/S vssd1 vssd1 vccd1 vccd1 _17232_/A sky130_fd_sc_hd__mux2_8
XANTENNA__14174__S _14180_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16191_ _13544_/X _19369_/Q _16191_/S vssd1 vssd1 vccd1 vccd1 _16192_/A sky130_fd_sc_hd__mux2_1
XFILLER_127_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_58_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15142_ _15142_/A vssd1 vssd1 vccd1 vccd1 _18993_/D sky130_fd_sc_hd__clkbuf_1
X_12354_ _12301_/X _12478_/B _12353_/Y vssd1 vssd1 vccd1 vccd1 _17886_/B sky130_fd_sc_hd__o21ai_4
XFILLER_127_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11305_ _11305_/A _11305_/B vssd1 vssd1 vccd1 vccd1 _11305_/X sky130_fd_sc_hd__or2_1
XFILLER_154_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15073_ _15073_/A vssd1 vssd1 vccd1 vccd1 _15073_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__14902__S _14904_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12285_ _12287_/A _12286_/A vssd1 vssd1 vccd1 vccd1 _12288_/A sky130_fd_sc_hd__and2_1
XFILLER_141_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11328__A1 _10639_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18901_ _19286_/CLK _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_113_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14024_ _18536_/Q _14023_/X _14027_/S vssd1 vssd1 vccd1 vccd1 _14025_/A sky130_fd_sc_hd__mux2_1
X_11236_ _19708_/Q vssd1 vssd1 vccd1 vccd1 _11236_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold7_A hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18832_ _19314_/CLK _18832_/D vssd1 vssd1 vccd1 vccd1 _18832_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_121_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11167_ _11160_/Y _11162_/Y _11164_/Y _11166_/Y _11044_/A vssd1 vssd1 vccd1 vccd1
+ _11167_/X sky130_fd_sc_hd__o221a_1
XFILLER_110_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10118_ _10174_/A _10117_/X _09823_/X vssd1 vssd1 vccd1 vccd1 _10118_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_49_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18763_ _19314_/CLK _18763_/D vssd1 vssd1 vccd1 vccd1 _18763_/Q sky130_fd_sc_hd__dfxtp_1
X_15975_ _13583_/X _19319_/Q _15981_/S vssd1 vssd1 vccd1 vccd1 _15976_/A sky130_fd_sc_hd__mux2_1
X_11098_ _11098_/A vssd1 vssd1 vccd1 vccd1 _11098_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16019__A1 _19333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17216__A0 _17722_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11187__S0 _11127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17714_ _17673_/X _17707_/X _17713_/Y _17571_/A vssd1 vssd1 vccd1 vccd1 _17714_/X
+ sky130_fd_sc_hd__o211a_1
X_14926_ _18909_/Q _14042_/X _14926_/S vssd1 vssd1 vccd1 vccd1 _14927_/A sky130_fd_sc_hd__mux2_1
X_10049_ _10042_/X _10044_/X _10046_/X _10048_/X _09752_/A vssd1 vssd1 vccd1 vccd1
+ _10049_/X sky130_fd_sc_hd__a221o_2
X_18694_ _19250_/CLK _18694_/D vssd1 vssd1 vccd1 vccd1 _18694_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17645_ _17390_/X _17827_/B _17644_/X _17333_/X vssd1 vssd1 vccd1 vccd1 _17645_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14857_ _14857_/A vssd1 vssd1 vccd1 vccd1 _18878_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13808_ _13808_/A vssd1 vssd1 vccd1 vccd1 _18467_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14788_ _15317_/B _15389_/B vssd1 vssd1 vccd1 vccd1 _14845_/A sky130_fd_sc_hd__nor2_2
XANTENNA__14450__A0 _13845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17576_ _17445_/X _17448_/X _17576_/S vssd1 vssd1 vccd1 vccd1 _17576_/X sky130_fd_sc_hd__mux2_1
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17519__B2 _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19315_ _19315_/CLK _19315_/D vssd1 vssd1 vccd1 vccd1 _19315_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16527_ _16529_/B _16529_/C _16526_/Y vssd1 vssd1 vccd1 vccd1 _19490_/D sky130_fd_sc_hd__o21a_1
XFILLER_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13739_ _13191_/X _18437_/Q _13747_/S vssd1 vssd1 vccd1 vccd1 _13740_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10178__A _19729_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10606__A3 _18828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14873__A _14930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12096__C _19402_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19246_ _19248_/CLK _19246_/D vssd1 vssd1 vccd1 vccd1 _19246_/Q sky130_fd_sc_hd__dfxtp_1
X_16458_ _16458_/A _19470_/Q _16458_/C vssd1 vssd1 vccd1 vccd1 _16460_/B sky130_fd_sc_hd__and3_1
XANTENNA__11016__B1 _09469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15409_ _19112_/Q _15025_/X _15411_/S vssd1 vssd1 vccd1 vccd1 _15410_/A sky130_fd_sc_hd__mux2_1
X_16389_ _19446_/Q _16389_/B vssd1 vssd1 vccd1 vccd1 _16396_/C sky130_fd_sc_hd__and2_1
X_19177_ _19239_/CLK _19177_/D vssd1 vssd1 vccd1 vccd1 _19177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_118_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10906__A _11220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12764__B1 _11354_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__S1 _09676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18128_ _18128_/A _18128_/B vssd1 vssd1 vccd1 vccd1 _18128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_129_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18059_ _19799_/Q _19420_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18060_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09607__S1 _09977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09901_ _10169_/A _09895_/Y _09900_/Y _09964_/A vssd1 vssd1 vccd1 vccd1 _09901_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_132_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09932__A1 _09690_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ _09817_/Y _09824_/Y _09826_/Y _09828_/Y _09831_/X vssd1 vssd1 vccd1 vccd1
+ _09832_/X sky130_fd_sc_hd__o221a_1
XFILLER_141_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _10296_/A vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__clkbuf_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11456__B _12457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11178__S0 _11127_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15643__S _15649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09694_ _10404_/A vssd1 vssd1 vccd1 vccd1 _09866_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10925__S0 _10862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12287__B _17856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10058__A1 _10056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15598__B _15598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13399__A hold21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14744__A1 _18828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ _19704_/Q _19703_/Q vssd1 vssd1 vccd1 vccd1 _09305_/B sky130_fd_sc_hd__or2_1
XFILLER_136_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_108_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15818__S _15826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14722__S _14726_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12070_ _12074_/A vssd1 vssd1 vccd1 vccd1 _15632_/S sky130_fd_sc_hd__buf_4
XFILLER_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11021_ _19303_/Q _18715_/Q _18752_/Q _18326_/Q _09624_/A _11020_/X vssd1 vssd1 vccd1
+ vccd1 _11021_/X sky130_fd_sc_hd__mux4_1
XFILLER_89_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10551__A _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__C1 _09465_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17997__A1 _19392_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15760_ _15760_/A vssd1 vssd1 vccd1 vccd1 _19223_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_131_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12972_ _13033_/A _12972_/B _13019_/C vssd1 vssd1 vccd1 vccd1 _12972_/X sky130_fd_sc_hd__or3_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input11_A io_dbus_rdata[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _11923_/A _17680_/A vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__xnor2_1
X_14711_ _14617_/X _18814_/Q _14713_/S vssd1 vssd1 vccd1 vccd1 _14712_/A sky130_fd_sc_hd__mux2_1
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15691_ _14595_/X _19193_/Q _15693_/S vssd1 vssd1 vccd1 vccd1 _15692_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14169__S _14169_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14371_/B _18091_/A _14642_/C _14642_/D vssd1 vssd1 vccd1 vccd1 _15782_/B
+ sky130_fd_sc_hd__and4b_2
X_17430_ _17831_/A vssd1 vssd1 vccd1 vccd1 _17430_/X sky130_fd_sc_hd__buf_2
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13235__A1 _12687_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11854_ _11854_/A _11854_/B vssd1 vssd1 vccd1 vccd1 _11855_/A sky130_fd_sc_hd__xnor2_4
XFILLER_73_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _11211_/A vssd1 vssd1 vccd1 vccd1 _11257_/A sky130_fd_sc_hd__clkbuf_2
X_14573_ _14573_/A vssd1 vssd1 vccd1 vccd1 _14573_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_17361_ _17261_/X _17213_/X _17372_/S vssd1 vssd1 vccd1 vccd1 _17361_/X sky130_fd_sc_hd__mux2_1
X_11785_ _11818_/S vssd1 vssd1 vccd1 vccd1 _11925_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_159_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10144__S1 _10090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13801__S _13809_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19100_ _19388_/CLK _19100_/D vssd1 vssd1 vccd1 vccd1 _19100_/Q sky130_fd_sc_hd__dfxtp_1
X_16312_ _19467_/Q _19466_/Q _19468_/Q _16443_/A vssd1 vssd1 vccd1 vccd1 _16453_/A
+ sky130_fd_sc_hd__and4_1
X_13524_ _13524_/A vssd1 vssd1 vccd1 vccd1 _18355_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16185__A0 _13535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17292_ _17232_/A _12487_/B _17293_/S vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__mux2_1
X_10736_ _10743_/A _10733_/X _10735_/X _09989_/A vssd1 vssd1 vccd1 vccd1 _10736_/X
+ sky130_fd_sc_hd__o211a_1
X_16243_ _16282_/A _16243_/B vssd1 vssd1 vccd1 vccd1 _16244_/A sky130_fd_sc_hd__and2_1
X_19031_ _19391_/CLK _19031_/D vssd1 vssd1 vccd1 vccd1 _19031_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13455_ _12945_/X _18328_/Q _13459_/S vssd1 vssd1 vccd1 vccd1 _13456_/A sky130_fd_sc_hd__mux2_1
XFILLER_12_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ _10667_/A _10667_/B vssd1 vssd1 vccd1 vccd1 _10667_/X sky130_fd_sc_hd__or2_1
XFILLER_127_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ _12419_/A _17906_/B vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__xnor2_4
XFILLER_173_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16174_ _13519_/X _19361_/Q _16180_/S vssd1 vssd1 vccd1 vccd1 _16175_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13386_ _14620_/A vssd1 vssd1 vccd1 vccd1 _13386_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10598_ _10598_/A _10598_/B vssd1 vssd1 vccd1 vccd1 _11452_/A sky130_fd_sc_hd__or2_1
XFILLER_154_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15125_ _15171_/S vssd1 vssd1 vccd1 vccd1 _15134_/S sky130_fd_sc_hd__buf_2
Xoutput108 _17175_/A vssd1 vssd1 vccd1 vccd1 io_dbus_st_type[1] sky130_fd_sc_hd__buf_2
X_12337_ _12347_/B _12337_/B vssd1 vssd1 vccd1 vccd1 _12337_/Y sky130_fd_sc_hd__xnor2_4
Xoutput119 _12467_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[19] sky130_fd_sc_hd__buf_2
XFILLER_141_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10772__A2 _10760_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15056_ _15056_/A vssd1 vssd1 vccd1 vccd1 _18961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12268_ _12312_/A _12268_/B vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__xnor2_4
X_14007_ _14579_/A vssd1 vssd1 vccd1 vccd1 _14007_/X sky130_fd_sc_hd__clkbuf_2
X_11219_ _18610_/Q _18945_/Q _11219_/S vssd1 vssd1 vccd1 vccd1 _11220_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11557__A _17175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19864_ _19865_/CLK _19864_/D vssd1 vssd1 vccd1 vccd1 _19864_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_122_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_96_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12199_ _12199_/A _12199_/B vssd1 vssd1 vccd1 vccd1 _12200_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11182__C1 _10949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 _12337_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[27] sky130_fd_sc_hd__buf_2
XFILLER_150_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18815_ _19297_/CLK _18815_/D vssd1 vssd1 vccd1 vccd1 _18815_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15999__B1 _13419_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10180__B _12471_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19795_ _19796_/CLK _19795_/D vssd1 vssd1 vccd1 vccd1 _19795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18746_ _19807_/CLK _18746_/D vssd1 vssd1 vccd1 vccd1 _18746_/Q sky130_fd_sc_hd__dfxtp_1
X_15958_ _15958_/A vssd1 vssd1 vccd1 vccd1 _19311_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10907__S0 _10904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ _18901_/Q _14017_/X _14915_/S vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16948__C1 _16933_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14079__S _14085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18677_ _18975_/CLK _18677_/D vssd1 vssd1 vccd1 vccd1 _18677_/Q sky130_fd_sc_hd__dfxtp_1
X_15889_ _15911_/A vssd1 vssd1 vccd1 vccd1 _15898_/S sky130_fd_sc_hd__buf_4
XFILLER_64_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17628_ _17630_/A _17630_/B vssd1 vssd1 vccd1 vccd1 _17628_/Y sky130_fd_sc_hd__nand2_1
XFILLER_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11237__B1 _09576_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17559_ _17563_/A _17563_/B _17775_/S vssd1 vssd1 vccd1 vccd1 _17559_/X sky130_fd_sc_hd__mux2_1
XANTENNA__18165__B2 _18081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__S0 _10579_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16176__A0 _13522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19229_ _19325_/CLK _19229_/D vssd1 vssd1 vccd1 vccd1 _19229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_164_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10355__B _12467_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16323__A _16848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17428__B1 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_141_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11712__A1 _19395_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input3_A io_dbus_rdata[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _11387_/A vssd1 vssd1 vccd1 vccd1 _09815_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09746_ _19326_/Q _18738_/Q _18775_/Q _18349_/Q _11374_/S _09687_/A vssd1 vssd1 vccd1
+ vccd1 _09747_/B sky130_fd_sc_hd__mux4_1
XFILLER_101_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_171_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ _09839_/A vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17600__A0 _17605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_186_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19180_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11323__S0 _09519_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15402__A _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11570_ _11575_/A _17175_/C vssd1 vssd1 vccd1 vccd1 _17168_/B sky130_fd_sc_hd__or2_1
XFILLER_23_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _10521_/A _10521_/B vssd1 vssd1 vccd1 vccd1 _10521_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13240_ _14595_/A vssd1 vssd1 vccd1 vccd1 _13240_/X sky130_fd_sc_hd__clkbuf_2
X_10452_ _10414_/A _10451_/X _10236_/A vssd1 vssd1 vccd1 vccd1 _10452_/X sky130_fd_sc_hd__a21o_1
XFILLER_108_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ _14582_/A vssd1 vssd1 vccd1 vccd1 _13171_/X sky130_fd_sc_hd__clkbuf_2
X_10383_ _10272_/A _10380_/Y _10382_/Y _10439_/A vssd1 vssd1 vccd1 vccd1 _10383_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14452__S _14456_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12122_ _12122_/A _12122_/B vssd1 vssd1 vccd1 vccd1 _12123_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_input59_A io_ibus_inst[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_124_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19416_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_123_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12480__B _12480_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16930_ _19628_/Q _12674_/X _16929_/X _16269_/X vssd1 vssd1 vccd1 vccd1 _19628_/D
+ sky130_fd_sc_hd__o211a_1
X_12053_ _12241_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _12054_/B sky130_fd_sc_hd__nor2_1
XFILLER_105_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11004_ _11171_/A _11004_/B vssd1 vssd1 vccd1 vccd1 _11004_/X sky130_fd_sc_hd__or2_1
XANTENNA__10062__S0 _09538_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16861_ _16862_/B _16862_/C _16860_/Y vssd1 vssd1 vccd1 vccd1 _19598_/D sky130_fd_sc_hd__o21a_1
XFILLER_78_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13592__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15283__S _15289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18600_ _19291_/CLK _18600_/D vssd1 vssd1 vccd1 vccd1 _18600_/Q sky130_fd_sc_hd__dfxtp_1
X_15812_ _15812_/A vssd1 vssd1 vccd1 vccd1 _19246_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_139_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19775_/CLK sky130_fd_sc_hd__clkbuf_16
X_19580_ _19583_/CLK _19580_/D vssd1 vssd1 vccd1 vccd1 _19580_/Q sky130_fd_sc_hd__dfxtp_1
X_16792_ _16840_/A _16800_/C vssd1 vssd1 vccd1 vccd1 _16792_/Y sky130_fd_sc_hd__nor2_1
XFILLER_92_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18531_ _19284_/CLK _18531_/D vssd1 vssd1 vccd1 vccd1 _18531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17186__B_N _17432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12955_ _13391_/A _12955_/B vssd1 vssd1 vccd1 vccd1 _12956_/B sky130_fd_sc_hd__nand2_1
X_15743_ _13560_/X _19216_/Q _15743_/S vssd1 vssd1 vccd1 vccd1 _15744_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10365__S1 _10229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _11915_/A _11969_/D vssd1 vssd1 vccd1 vccd1 _11934_/B sky130_fd_sc_hd__nand2_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _19309_/CLK _18462_/D vssd1 vssd1 vccd1 vccd1 _18462_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ _14569_/X _19185_/Q _15682_/S vssd1 vssd1 vccd1 vccd1 _15675_/A sky130_fd_sc_hd__mux2_1
X_12886_ _14534_/A vssd1 vssd1 vccd1 vccd1 _12886_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_34_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17413_/A vssd1 vssd1 vccd1 vccd1 _17413_/X sky130_fd_sc_hd__clkbuf_2
X_11837_ _19399_/Q _11793_/X _11829_/X _11836_/Y vssd1 vssd1 vccd1 vccd1 _16258_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14625_ _14635_/A _18205_/B vssd1 vssd1 vccd1 vccd1 _14626_/A sky130_fd_sc_hd__and2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18393_ _19308_/CLK _18393_/D vssd1 vssd1 vccd1 vccd1 _18393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11314__S0 _10030_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11840__A _11840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14556_ _14556_/A vssd1 vssd1 vccd1 vccd1 _18757_/D sky130_fd_sc_hd__clkbuf_1
X_17344_ _17367_/S _17344_/B vssd1 vssd1 vccd1 vccd1 _17344_/X sky130_fd_sc_hd__and2b_1
XFILLER_60_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11768_ _19397_/Q _11768_/B vssd1 vssd1 vccd1 vccd1 _11769_/A sky130_fd_sc_hd__and2_1
XFILLER_146_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10719_ _10719_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10719_/Y sky130_fd_sc_hd__nor2_1
X_13507_ _13386_/X _18352_/Q _13507_/S vssd1 vssd1 vccd1 vccd1 _13508_/A sky130_fd_sc_hd__mux2_1
X_14487_ _13899_/X _18728_/Q _14489_/S vssd1 vssd1 vccd1 vccd1 _14488_/A sky130_fd_sc_hd__mux2_1
X_17275_ _17810_/B _17662_/B _17293_/S vssd1 vssd1 vccd1 vccd1 _17275_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12719__A0 _18107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11699_ _11699_/A vssd1 vssd1 vccd1 vccd1 _12974_/A sky130_fd_sc_hd__buf_2
XFILLER_173_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19014_ _19329_/CLK _19014_/D vssd1 vssd1 vccd1 vccd1 _19014_/Q sky130_fd_sc_hd__dfxtp_1
X_13438_ _13494_/A vssd1 vssd1 vccd1 vccd1 _13507_/S sky130_fd_sc_hd__buf_6
X_16226_ _16226_/A vssd1 vssd1 vccd1 vccd1 _16235_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_174_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16157_ _16156_/X _19357_/Q _16167_/S vssd1 vssd1 vccd1 vccd1 _16158_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13767__A _13835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17239__A _17239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ _13369_/A vssd1 vssd1 vccd1 vccd1 _18313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19161__CLK _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15108_ _18978_/Q _15006_/X _15112_/S vssd1 vssd1 vccd1 vccd1 _15109_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16088_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16112_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_88_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_142_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15039_ _18956_/Q _15038_/X _15045_/S vssd1 vssd1 vccd1 vccd1 _15040_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10191__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19847_ _19865_/CLK _19847_/D vssd1 vssd1 vccd1 vccd1 _19847_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09994__S0 _09850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09600_ _09600_/A vssd1 vssd1 vccd1 vccd1 _09977_/A sky130_fd_sc_hd__buf_2
XFILLER_84_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19778_ _19780_/CLK _19778_/D vssd1 vssd1 vccd1 vccd1 _19778_/Q sky130_fd_sc_hd__dfxtp_1
X_09531_ _09531_/A vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__buf_2
X_18729_ _19124_/CLK _18729_/D vssd1 vssd1 vccd1 vccd1 _18729_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17189__A2 _12432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10356__S1 _10229_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _10236_/A _09459_/X _09461_/X _09737_/A vssd1 vssd1 vccd1 vccd1 _09462_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _09393_/A vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_52_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11630__A0 _11619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15368__S _15372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19282_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__13677__A _13677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17149__A _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19285_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_86_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14301__A _14369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09729_ _09844_/A vssd1 vssd1 vccd1 vccd1 _09730_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__11644__B _11644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15831__S _15837_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12740_ _12747_/A vssd1 vssd1 vccd1 vccd1 _12740_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_83_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09114__B _18081_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12671_ _16341_/A _19587_/Q _16921_/S _12670_/X vssd1 vssd1 vccd1 vccd1 _19587_/D
+ sky130_fd_sc_hd__o31a_1
XFILLER_15_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17331__B _17432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14410_/A vssd1 vssd1 vccd1 vccd1 _18693_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ _13411_/A _11794_/A _12175_/A vssd1 vssd1 vccd1 vccd1 _11622_/X sky130_fd_sc_hd__and3_1
XFILLER_169_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15390_ _15446_/A vssd1 vssd1 vccd1 vccd1 _15459_/S sky130_fd_sc_hd__buf_6
XFILLER_23_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14341_ _13899_/X _18664_/Q _14343_/S vssd1 vssd1 vccd1 vccd1 _14342_/A sky130_fd_sc_hd__mux2_1
X_11553_ _12175_/A _14275_/C vssd1 vssd1 vccd1 vccd1 _11553_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09290__A1 _12543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17060_ _17060_/A vssd1 vssd1 vccd1 vccd1 _19677_/D sky130_fd_sc_hd__clkbuf_1
X_10504_ _18400_/Q _18661_/Q _18560_/Q _18895_/Q _09980_/S _10310_/A vssd1 vssd1 vccd1
+ vccd1 _10505_/B sky130_fd_sc_hd__mux4_1
X_14272_ _14272_/A _18250_/Q vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__nor2_1
XFILLER_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11484_ _11567_/A vssd1 vssd1 vccd1 vccd1 _17183_/A sky130_fd_sc_hd__clkbuf_2
X_16011_ _16011_/A _16011_/B _16011_/C vssd1 vssd1 vccd1 vccd1 _16021_/C sky130_fd_sc_hd__or3_2
XFILLER_171_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13223_ _19729_/Q _15586_/B _13306_/A vssd1 vssd1 vccd1 vccd1 _13223_/X sky130_fd_sc_hd__mux2_1
XANTENNA__15278__S _15278_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10435_ _18626_/Q _18961_/Q _10435_/S vssd1 vssd1 vccd1 vccd1 _10436_/B sky130_fd_sc_hd__mux2_1
XFILLER_109_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12491__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_3_7_0_clock clkbuf_3_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_7_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_128_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13154_ _13154_/A vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10366_ _10419_/A _10366_/B vssd1 vssd1 vccd1 vccd1 _10366_/X sky130_fd_sc_hd__or2_1
XANTENNA__11819__B _17245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output165_A _12418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16898__A _16914_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12105_ _19648_/Q _19647_/Q _12105_/C vssd1 vssd1 vccd1 vccd1 _12156_/C sky130_fd_sc_hd__and3_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10215__S _10215_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _16069_/A _13083_/B _12861_/A vssd1 vssd1 vccd1 vccd1 _13086_/B sky130_fd_sc_hd__o21ai_1
X_17962_ _19755_/Q _19787_/Q _17968_/S vssd1 vssd1 vccd1 vccd1 _17963_/A sky130_fd_sc_hd__mux2_1
X_10297_ _10297_/A vssd1 vssd1 vccd1 vccd1 _10297_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_105_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19701_ _19706_/CLK _19701_/D vssd1 vssd1 vccd1 vccd1 _19701_/Q sky130_fd_sc_hd__dfxtp_4
X_16913_ _16912_/B _16912_/C _19617_/Q vssd1 vssd1 vccd1 vccd1 _16914_/C sky130_fd_sc_hd__a21oi_1
X_12036_ _19407_/Q vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__buf_2
XFILLER_78_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17893_ _17852_/X _17484_/Y _17892_/Y _17860_/X vssd1 vssd1 vccd1 vccd1 _17893_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13526__S _13529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19632_ _19635_/CLK _19632_/D vssd1 vssd1 vccd1 vccd1 _19632_/Q sky130_fd_sc_hd__dfxtp_1
X_16844_ _18079_/B vssd1 vssd1 vccd1 vccd1 _16881_/A sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_181_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14211__A _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19563_ _19564_/CLK _19563_/D vssd1 vssd1 vccd1 vccd1 _19563_/Q sky130_fd_sc_hd__dfxtp_1
X_16775_ _16782_/C _16782_/D _16764_/X vssd1 vssd1 vccd1 vccd1 _16775_/Y sky130_fd_sc_hd__a21oi_1
X_13987_ _13987_/A vssd1 vssd1 vccd1 vccd1 _18524_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_81_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12101__A1 _12092_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15741__S _15743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18514_ _19267_/CLK _18514_/D vssd1 vssd1 vccd1 vccd1 _18514_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15726_ _13535_/X _19208_/Q _15732_/S vssd1 vssd1 vccd1 vccd1 _15727_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12938_ _19495_/Q _13054_/A _12936_/X _12937_/X vssd1 vssd1 vccd1 vccd1 _12938_/X
+ sky130_fd_sc_hd__a22o_1
X_19494_ _19619_/CLK _19494_/D vssd1 vssd1 vccd1 vccd1 _19494_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18445_ _19264_/CLK _18445_/D vssd1 vssd1 vccd1 vccd1 _18445_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15657_ _15657_/A vssd1 vssd1 vccd1 vccd1 _19177_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14357__S _14365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12869_ _16011_/B _12891_/C vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__xor2_1
XFILLER_61_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14608_ _14608_/A vssd1 vssd1 vccd1 vccd1 _14608_/X sky130_fd_sc_hd__clkbuf_2
X_18376_ _19383_/CLK _18376_/D vssd1 vssd1 vccd1 vccd1 _18376_/Q sky130_fd_sc_hd__dfxtp_1
X_15588_ _15565_/X _15586_/X _15587_/Y _12575_/X _18273_/Q vssd1 vssd1 vccd1 vccd1
+ _15588_/X sky130_fd_sc_hd__a32o_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17327_ _17471_/A _17327_/B vssd1 vssd1 vccd1 vccd1 _17328_/C sky130_fd_sc_hd__nand2_1
XFILLER_105_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ _14537_/X _18752_/Q _14551_/S vssd1 vssd1 vccd1 vccd1 _14540_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10510__S1 _09710_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09975__A _09975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17258_ _17480_/A vssd1 vssd1 vccd1 vccd1 _17504_/S sky130_fd_sc_hd__buf_2
XFILLER_146_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16209_ _13570_/X _19377_/Q _16213_/S vssd1 vssd1 vccd1 vccd1 _16210_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14092__S _14096_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17189_ _12429_/A _12432_/A _12432_/B _17188_/X vssd1 vssd1 vccd1 vccd1 _17328_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15106__A1 _15003_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_103_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15916__S _15920_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09741__C1 _09740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _10855_/A vssd1 vssd1 vccd1 vccd1 _10623_/A sky130_fd_sc_hd__buf_2
XFILLER_65_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17031__A1 _13404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09445_ _10042_/A _09445_/B vssd1 vssd1 vccd1 vccd1 _09445_/X sky130_fd_sc_hd__or2_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15593__A1 _19161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09376_ _11012_/A vssd1 vssd1 vccd1 vccd1 _10990_/A sky130_fd_sc_hd__buf_2
XFILLER_21_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09885__A _10521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_166_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_153_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10220_ _18598_/Q _18869_/Q _19093_/Q _18837_/Q _10112_/S _09905_/A vssd1 vssd1 vccd1
+ vccd1 _10220_/X sky130_fd_sc_hd__mux4_1
XFILLER_165_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15826__S _15826_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10151_ _18471_/Q _19062_/Q _19224_/Q _18439_/Q _09930_/S _10090_/X vssd1 vssd1 vccd1
+ vccd1 _10151_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11119__C1 _10929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09958__S0 _10168_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ _10082_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _10082_/X sky130_fd_sc_hd__or2_1
XFILLER_102_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10568__S1 _10567_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ _13909_/X _18502_/Q _13919_/S vssd1 vssd1 vccd1 vccd1 _13911_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14890_ _14890_/A vssd1 vssd1 vccd1 vccd1 _18892_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_87_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17270__A1 _17630_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _13922_/A vssd1 vssd1 vccd1 vccd1 _13941_/S sky130_fd_sc_hd__buf_6
XFILLER_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16560_ _16585_/A _16560_/B _16561_/B vssd1 vssd1 vccd1 vccd1 _19500_/D sky130_fd_sc_hd__nor3_1
X_13772_ _12851_/X _18451_/Q _13776_/S vssd1 vssd1 vccd1 vccd1 _13773_/A sky130_fd_sc_hd__mux2_1
X_10984_ _10977_/Y _10979_/Y _10981_/Y _10983_/Y _09571_/A vssd1 vssd1 vccd1 vccd1
+ _10984_/X sky130_fd_sc_hd__o221a_2
XFILLER_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17022__A1 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15511_ _15510_/X _19146_/Q _15517_/S vssd1 vssd1 vccd1 vccd1 _15512_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12723_ _12723_/A vssd1 vssd1 vccd1 vccd1 _18251_/D sky130_fd_sc_hd__clkbuf_1
X_16491_ _16493_/A _16493_/C _16490_/Y vssd1 vssd1 vccd1 vccd1 _19481_/D sky130_fd_sc_hd__o21a_1
XFILLER_128_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18230_ input52/X _18197_/X _18229_/X _18193_/X _18135_/A vssd1 vssd1 vccd1 vccd1
+ _18231_/B sky130_fd_sc_hd__a32o_1
XANTENNA__15584__A1 _19159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12654_ _14275_/A _12654_/B vssd1 vssd1 vccd1 vccd1 _17102_/B sky130_fd_sc_hd__or2_2
X_15442_ _19127_/Q _15073_/X _15444_/S vssd1 vssd1 vccd1 vccd1 _15443_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12398__A1 _18144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11605_ _19772_/Q _11239_/A _11678_/A vssd1 vssd1 vccd1 vccd1 _17230_/A sky130_fd_sc_hd__mux2_4
XFILLER_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18161_ _18161_/A vssd1 vssd1 vccd1 vccd1 _19838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_169_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12585_ _16622_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _12586_/B sky130_fd_sc_hd__nor2_2
X_15373_ _15373_/A vssd1 vssd1 vccd1 vccd1 _19096_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_128_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17112_ _17112_/A vssd1 vssd1 vccd1 vccd1 _17130_/B sky130_fd_sc_hd__inv_2
XANTENNA__09795__A _09964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14324_ _13873_/X _18656_/Q _14332_/S vssd1 vssd1 vccd1 vccd1 _14325_/A sky130_fd_sc_hd__mux2_1
X_11536_ _11536_/A vssd1 vssd1 vccd1 vccd1 _18742_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18092_ _19844_/Q _12694_/X _18091_/Y _18084_/X vssd1 vssd1 vccd1 vccd1 _19812_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11070__B2 _19711_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17043_ _17043_/A vssd1 vssd1 vccd1 vccd1 _19669_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14255_ _14255_/A vssd1 vssd1 vccd1 vccd1 _14264_/S sky130_fd_sc_hd__buf_4
XFILLER_144_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11467_ _11467_/A _11467_/B _11467_/C vssd1 vssd1 vccd1 vccd1 _11470_/B sky130_fd_sc_hd__or3_1
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13206_ input14/X _13166_/X _13167_/X vssd1 vssd1 vccd1 vccd1 _13206_/Y sky130_fd_sc_hd__a21oi_2
X_10418_ _18402_/Q _18663_/Q _18562_/Q _18897_/Q _10368_/S _09674_/A vssd1 vssd1 vccd1
+ vccd1 _10419_/B sky130_fd_sc_hd__mux4_1
XFILLER_136_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_125_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14186_ _14186_/A vssd1 vssd1 vccd1 vccd1 _18603_/D sky130_fd_sc_hd__clkbuf_1
X_11398_ _09767_/X _11391_/X _11393_/Y _11397_/Y _09813_/X vssd1 vssd1 vccd1 vccd1
+ _11398_/X sky130_fd_sc_hd__o311a_1
XFILLER_152_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16297__C1 _16269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13137_ _15054_/A vssd1 vssd1 vccd1 vccd1 _14576_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__09971__C1 _09831_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _18596_/Q _18867_/Q _19091_/Q _18835_/Q _10341_/S _10436_/A vssd1 vssd1 vccd1
+ vccd1 _10349_/X sky130_fd_sc_hd__mux4_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17517__A _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18994_ _19089_/CLK _18994_/D vssd1 vssd1 vccd1 vccd1 _18994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_98_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18038__A0 _19790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10008__S0 _09776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17945_/A vssd1 vssd1 vccd1 vccd1 _19747_/D sky130_fd_sc_hd__clkbuf_1
X_13068_ _13051_/X _13066_/X _13067_/X vssd1 vssd1 vccd1 vccd1 _15041_/A sky130_fd_sc_hd__o21a_4
XFILLER_39_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12019_ _19406_/Q _11665_/X _12014_/Y _12018_/X vssd1 vssd1 vccd1 vccd1 _16274_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_39_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10333__B1 _09822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17876_ _17878_/A _17878_/B vssd1 vssd1 vccd1 vccd1 _17876_/Y sky130_fd_sc_hd__nand2_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19615_ _19618_/CLK _19615_/D vssd1 vssd1 vccd1 vccd1 _19615_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17261__A1 _17743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16827_ _19582_/Q _16827_/B vssd1 vssd1 vccd1 vccd1 _16830_/B sky130_fd_sc_hd__nand2_1
XFILLER_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11284__B _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_94_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17252__A _17252_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19546_ _19549_/CLK _19546_/D vssd1 vssd1 vccd1 vccd1 _19546_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16758_ _19561_/Q _19560_/Q _16758_/C vssd1 vssd1 vccd1 vccd1 _16767_/C sky130_fd_sc_hd__and3_1
XFILLER_0_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15709_ _15709_/A vssd1 vssd1 vccd1 vccd1 _19201_/D sky130_fd_sc_hd__clkbuf_1
X_19477_ _19610_/CLK _19477_/D vssd1 vssd1 vccd1 vccd1 _19477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16689_ _19539_/Q _19538_/Q _16689_/C _16689_/D vssd1 vssd1 vccd1 vccd1 _16697_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_22_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09230_ _09575_/B _09230_/B _11508_/A vssd1 vssd1 vccd1 vccd1 _09230_/X sky130_fd_sc_hd__and3b_1
X_18428_ _19309_/CLK _18428_/D vssd1 vssd1 vccd1 vccd1 _18428_/Q sky130_fd_sc_hd__dfxtp_1
X_09161_ _11528_/A vssd1 vssd1 vccd1 vccd1 _18100_/A sky130_fd_sc_hd__buf_4
X_18359_ _19241_/CLK _18359_/D vssd1 vssd1 vccd1 vccd1 _18359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18083__A _18083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14815__S _14821_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17316__A2 _12487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09092_ _19841_/Q _09182_/B _19839_/Q vssd1 vssd1 vccd1 vccd1 _11646_/B sky130_fd_sc_hd__or3_2
XFILLER_148_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12010__B1 _19406_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09962__C1 _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09994_ _19324_/Q _18736_/Q _18773_/Q _18347_/Q _09850_/A _09977_/X vssd1 vssd1 vccd1
+ vccd1 _09994_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15381__S _15383_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17004__A1 _12689_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10819__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10722__S1 _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09428_ _10042_/A vssd1 vssd1 vccd1 vccd1 _10514_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_40_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09359_ _17795_/A vssd1 vssd1 vccd1 vccd1 _09359_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_138_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11052__A1 _09416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10486__S0 _10274_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ _19420_/Q _12371_/B vssd1 vssd1 vccd1 vccd1 _12372_/B sky130_fd_sc_hd__nor2_1
XFILLER_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_138_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11321_ _11321_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11321_/Y sky130_fd_sc_hd__nand2_1
XFILLER_60_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14040_ _18541_/Q _14039_/X _14043_/S vssd1 vssd1 vccd1 vccd1 _14041_/A sky130_fd_sc_hd__mux2_1
XFILLER_153_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11252_ _11252_/A _11252_/B vssd1 vssd1 vccd1 vccd1 _11252_/X sky130_fd_sc_hd__or2_1
XFILLER_107_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _09667_/A _10193_/X _10202_/X _09758_/A _19728_/Q vssd1 vssd1 vccd1 vccd1
+ _11354_/A sky130_fd_sc_hd__a32o_4
XANTENNA__10012__C1 _09829_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ _19173_/Q _18787_/Q _19237_/Q _18356_/Q _11127_/S _11177_/X vssd1 vssd1 vccd1
+ vccd1 _11184_/B sky130_fd_sc_hd__mux4_1
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input41_A io_ibus_inst[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10134_ _09762_/X _10123_/X _10132_/X _09835_/X _10133_/Y vssd1 vssd1 vccd1 vccd1
+ _12472_/B sky130_fd_sc_hd__o32a_4
XFILLER_122_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15991_ _15991_/A vssd1 vssd1 vccd1 vccd1 _19326_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17730_ _17730_/A vssd1 vssd1 vccd1 vccd1 _17730_/Y sky130_fd_sc_hd__clkinv_2
X_14942_ _18917_/Q vssd1 vssd1 vccd1 vccd1 _14943_/A sky130_fd_sc_hd__clkbuf_1
X_10065_ _09485_/A _10052_/Y _10058_/X _10064_/Y _09811_/A vssd1 vssd1 vccd1 vccd1
+ _10065_/X sky130_fd_sc_hd__o311a_4
XFILLER_102_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10866__A1 _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17661_ _17662_/A _17662_/B _17842_/S vssd1 vssd1 vccd1 vccd1 _17661_/X sky130_fd_sc_hd__mux2_1
X_14873_ _14930_/S vssd1 vssd1 vccd1 vccd1 _14882_/S sky130_fd_sc_hd__buf_2
XFILLER_75_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18168__A _18188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19400_ _19838_/CLK _19400_/D vssd1 vssd1 vccd1 vccd1 _19400_/Q sky130_fd_sc_hd__dfxtp_1
X_16612_ _16714_/A vssd1 vssd1 vccd1 vccd1 _16666_/A sky130_fd_sc_hd__buf_2
XFILLER_29_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13824_ _13824_/A vssd1 vssd1 vccd1 vccd1 _18474_/D sky130_fd_sc_hd__clkbuf_1
X_17592_ _17592_/A vssd1 vssd1 vccd1 vccd1 _17592_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_91_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19331_ _19423_/CLK _19331_/D vssd1 vssd1 vccd1 vccd1 _19331_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_90_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16543_ _16553_/D vssd1 vssd1 vccd1 vccd1 _16551_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10967_ _18583_/Q _18854_/Q _19078_/Q _18822_/Q _10862_/X _09513_/A vssd1 vssd1 vccd1
+ vccd1 _10967_/X sky130_fd_sc_hd__mux4_1
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13755_ _13755_/A vssd1 vssd1 vccd1 vccd1 _18444_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12706_ _12696_/A _12619_/A _12702_/X _12705_/X vssd1 vssd1 vccd1 vccd1 _12706_/X
+ sky130_fd_sc_hd__a211o_1
X_19262_ _19388_/CLK _19262_/D vssd1 vssd1 vccd1 vccd1 _19262_/Q sky130_fd_sc_hd__dfxtp_1
X_16474_ _16474_/A _19476_/Q _16474_/C vssd1 vssd1 vccd1 vccd1 _16476_/B sky130_fd_sc_hd__and3_1
X_10898_ _11151_/S vssd1 vssd1 vccd1 vccd1 _10964_/S sky130_fd_sc_hd__clkbuf_4
X_13686_ _13349_/X _18414_/Q _13686_/S vssd1 vssd1 vccd1 vccd1 _13687_/A sky130_fd_sc_hd__mux2_1
XFILLER_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18213_ _18213_/A _18213_/B vssd1 vssd1 vccd1 vccd1 _18214_/A sky130_fd_sc_hd__and2_1
XFILLER_31_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15425_ _19119_/Q _15047_/X _15433_/S vssd1 vssd1 vccd1 vccd1 _15426_/A sky130_fd_sc_hd__mux2_1
X_12637_ _19563_/Q vssd1 vssd1 vccd1 vccd1 _16772_/C sky130_fd_sc_hd__clkbuf_2
X_19193_ _19383_/CLK _19193_/D vssd1 vssd1 vccd1 vccd1 _19193_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12944__A _15022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18144_ _18144_/A _18146_/B vssd1 vssd1 vccd1 vccd1 _18144_/X sky130_fd_sc_hd__or2_1
X_12568_ _19627_/Q _16931_/A _12526_/X _19155_/Q _12567_/X vssd1 vssd1 vccd1 vccd1
+ _12568_/X sky130_fd_sc_hd__a221o_1
X_15356_ _15356_/A vssd1 vssd1 vccd1 vccd1 _19088_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_172_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14307_ _14307_/A vssd1 vssd1 vccd1 vccd1 _18648_/D sky130_fd_sc_hd__clkbuf_1
X_11519_ _19845_/Q _19844_/Q _19843_/Q _18087_/A vssd1 vssd1 vccd1 vccd1 _11521_/C
+ sky130_fd_sc_hd__or4_1
X_18075_ _18075_/A _18087_/B vssd1 vssd1 vccd1 vccd1 _18075_/X sky130_fd_sc_hd__or2_1
XFILLER_129_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15287_ _14579_/X _19058_/Q _15289_/S vssd1 vssd1 vccd1 vccd1 _15288_/A sky130_fd_sc_hd__mux2_1
XFILLER_145_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12499_ _19604_/Q vssd1 vssd1 vccd1 vccd1 _16879_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17026_ _19663_/Q _16935_/A _17026_/S vssd1 vssd1 vccd1 vccd1 _17027_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14238_ _18626_/Q _14004_/X _14242_/S vssd1 vssd1 vccd1 vccd1 _14239_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14169_ _18596_/Q _14010_/X _14169_/S vssd1 vssd1 vccd1 vccd1 _14170_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17247__A _17247_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17482__A1 _17731_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _19724_/CLK _18977_/D vssd1 vssd1 vccd1 vccd1 _18977_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17928_ _17928_/A vssd1 vssd1 vccd1 vccd1 _19739_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17859_ _17478_/X _17578_/X _17858_/X _17633_/X vssd1 vssd1 vccd1 vccd1 _17859_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_27_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17785__A2 _17652_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10952__S1 _10937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10609__A1 _10614_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19529_ _19529_/CLK _19529_/D vssd1 vssd1 vccd1 vccd1 _19529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11282__A1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__B2 _09311_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09213_ _09213_/A vssd1 vssd1 vccd1 vccd1 _17145_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_139_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10490__C1 _09812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12854__A _18744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16326__A _16344_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09144_ _19866_/Q vssd1 vssd1 vccd1 vccd1 _18146_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12231__B1 _12230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_162_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10793__B1 _09484_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_146_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12534__A1 _19628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09977_ _09977_/A vssd1 vssd1 vccd1 vccd1 _09977_/X sky130_fd_sc_hd__buf_2
XFILLER_77_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10313__S _10315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12837__A2 _12703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_opt_5_0_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_6_0_clock clkbuf_4_7_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_73_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11870_ _17642_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _11873_/A sky130_fd_sc_hd__xor2_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _09432_/A _10804_/X _10809_/X _10820_/X _09614_/A vssd1 vssd1 vccd1 vccd1
+ _10821_/X sky130_fd_sc_hd__a311o_2
XANTENNA__09403__A _11254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ _19179_/Q _18793_/Q _19243_/Q _18362_/Q _10729_/S _11298_/A vssd1 vssd1 vccd1
+ vccd1 _10753_/B sky130_fd_sc_hd__mux4_1
X_13540_ _13540_/A vssd1 vssd1 vccd1 vccd1 _18360_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13471_ _13471_/A vssd1 vssd1 vccd1 vccd1 _18335_/D sky130_fd_sc_hd__clkbuf_1
X_10683_ _19181_/Q _18795_/Q _19245_/Q _18364_/Q _10576_/X _10577_/X vssd1 vssd1 vccd1
+ vccd1 _10684_/B sky130_fd_sc_hd__mux4_1
X_15210_ _15210_/A vssd1 vssd1 vccd1 vccd1 _19023_/D sky130_fd_sc_hd__clkbuf_1
X_12422_ _12422_/A vssd1 vssd1 vccd1 vccd1 _12422_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16190_ _16190_/A vssd1 vssd1 vccd1 vccd1 _19368_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15141_ _18993_/Q _15054_/X _15145_/S vssd1 vssd1 vccd1 vccd1 _15142_/A sky130_fd_sc_hd__mux2_1
X_12353_ _18140_/A _11516_/X _12302_/X vssd1 vssd1 vccd1 vccd1 _12353_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_153_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11304_ _18398_/Q _18659_/Q _18558_/Q _18893_/Q _10660_/A _09442_/A vssd1 vssd1 vccd1
+ vccd1 _11305_/B sky130_fd_sc_hd__mux4_1
X_15072_ _15072_/A vssd1 vssd1 vccd1 vccd1 _18966_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_142_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12284_ _19796_/Q _09975_/A _12357_/S vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__mux2_8
X_18900_ _18902_/CLK _18900_/D vssd1 vssd1 vccd1 vccd1 _18900_/Q sky130_fd_sc_hd__dfxtp_1
X_14023_ _14595_/A vssd1 vssd1 vccd1 vccd1 _14023_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11235_ _11228_/Y _11230_/Y _11232_/Y _11234_/Y _10929_/A vssd1 vssd1 vccd1 vccd1
+ _11235_/X sky130_fd_sc_hd__o221a_1
XANTENNA__13595__A _15079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18831_ _19249_/CLK _18831_/D vssd1 vssd1 vccd1 vccd1 _18831_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17464__A1 _17907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ _11085_/A _11165_/X _10915_/X vssd1 vssd1 vccd1 vccd1 _11166_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15475__B1 _13423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10117_ _18935_/Q _18701_/Q _19383_/Q _19031_/Q _09918_/X _09900_/A vssd1 vssd1 vccd1
+ vccd1 _10117_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18762_ _19249_/CLK _18762_/D vssd1 vssd1 vccd1 vccd1 _18762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15974_ _15974_/A vssd1 vssd1 vccd1 vccd1 _19318_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11097_ _18483_/Q _18978_/Q _11263_/S vssd1 vssd1 vccd1 vccd1 _11098_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17216__A1 _17215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17713_ _17413_/X _17710_/X _17712_/X vssd1 vssd1 vccd1 vccd1 _17713_/Y sky130_fd_sc_hd__o21ai_1
X_10048_ _09993_/A _10047_/X _09989_/X vssd1 vssd1 vccd1 vccd1 _10048_/X sky130_fd_sc_hd__o21a_1
X_14925_ _14925_/A vssd1 vssd1 vccd1 vccd1 _18908_/D sky130_fd_sc_hd__clkbuf_1
X_18693_ _19119_/CLK _18693_/D vssd1 vssd1 vccd1 vccd1 _18693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17644_ _17413_/X _17641_/X _17643_/Y _17532_/X vssd1 vssd1 vccd1 vccd1 _17644_/X
+ sky130_fd_sc_hd__o211a_1
X_14856_ _18878_/Q _14045_/X _14858_/S vssd1 vssd1 vccd1 vccd1 _14857_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13807_ _13148_/X _18467_/Q _13809_/S vssd1 vssd1 vccd1 vccd1 _13808_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17575_ _17446_/X _17439_/A _17575_/S vssd1 vssd1 vccd1 vccd1 _17730_/A sky130_fd_sc_hd__mux2_1
XFILLER_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14787_ _18089_/A _14787_/B vssd1 vssd1 vccd1 vccd1 _15389_/B sky130_fd_sc_hd__nand2_2
XFILLER_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11999_ _17696_/A _12025_/B _17709_/A _12111_/A vssd1 vssd1 vccd1 vccd1 _12000_/B
+ sky130_fd_sc_hd__o31a_1
X_19314_ _19314_/CLK _19314_/D vssd1 vssd1 vccd1 vccd1 _19314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16526_ _16529_/B _16529_/C _16489_/X vssd1 vssd1 vccd1 vccd1 _16526_/Y sky130_fd_sc_hd__a21oi_1
X_13738_ _13749_/A vssd1 vssd1 vccd1 vccd1 _13747_/S sky130_fd_sc_hd__buf_6
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17924__C1 _12744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19245_ _19245_/CLK _19245_/D vssd1 vssd1 vccd1 vccd1 _19245_/Q sky130_fd_sc_hd__dfxtp_1
X_16457_ _16458_/A _16458_/C _16456_/Y vssd1 vssd1 vccd1 vccd1 _19469_/D sky130_fd_sc_hd__o21a_1
X_13669_ _13209_/X _18406_/Q _13675_/S vssd1 vssd1 vccd1 vccd1 _13670_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14365__S _14365_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16146__A _16146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11016__A1 _09366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15408_ _15408_/A vssd1 vssd1 vccd1 vccd1 _19111_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_118_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19176_ _19241_/CLK _19176_/D vssd1 vssd1 vccd1 vccd1 _19176_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11016__B2 _19712_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16388_ _16388_/A _16388_/B _16389_/B vssd1 vssd1 vccd1 vccd1 _19445_/D sky130_fd_sc_hd__nor3_1
XFILLER_157_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18127_ _18127_/A vssd1 vssd1 vccd1 vccd1 _18128_/A sky130_fd_sc_hd__inv_2
XANTENNA__10224__C1 _09813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15339_ _19081_/Q _15028_/X _15339_/S vssd1 vssd1 vccd1 vccd1 _15340_/A sky130_fd_sc_hd__mux2_1
XFILLER_144_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18058_ _18058_/A vssd1 vssd1 vccd1 vccd1 _19798_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10870__S0 _10873_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17009_ _15600_/X _16997_/X _17007_/X _17008_/X vssd1 vssd1 vccd1 vccd1 _19656_/D
+ sky130_fd_sc_hd__o211a_1
X_09900_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_125_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10922__A _11116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18101__C1 _18097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09831_ _09831_/A vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_140_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_141_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15924__S _15924_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09762_/A vssd1 vssd1 vccd1 vccd1 _09762_/X sky130_fd_sc_hd__buf_2
XANTENNA__12819__A2 _12603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _10511_/A vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13444__S _13448_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10925__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17915__C1 _12744_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13399__B _13399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ input70/X vssd1 vssd1 vccd1 vccd1 _16245_/A sky130_fd_sc_hd__buf_4
XFILLER_109_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11020_ _11020_/A vssd1 vssd1 vccd1 vccd1 _11020_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_173_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10613__S0 _10546_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _19747_/Q _12971_/B vssd1 vssd1 vccd1 vccd1 _13019_/C sky130_fd_sc_hd__and2_1
XANTENNA__12759__A _12773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14710_ _14710_/A vssd1 vssd1 vccd1 vccd1 _18813_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11922_ _11942_/A _12457_/B _11890_/C _11921_/X vssd1 vssd1 vccd1 vccd1 _17680_/A
+ sky130_fd_sc_hd__a22o_2
XFILLER_57_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15690_ _15690_/A vssd1 vssd1 vccd1 vccd1 _19192_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12478__B _12478_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14641_ _14641_/A vssd1 vssd1 vccd1 vccd1 _18783_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _11791_/A _11790_/A _11824_/A _11852_/X vssd1 vssd1 vccd1 vccd1 _11854_/B
+ sky130_fd_sc_hd__a31o_4
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10279__A _10479_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17360_ _17351_/Y _17359_/Y _17653_/A vssd1 vssd1 vccd1 vccd1 _17360_/X sky130_fd_sc_hd__mux2_1
X_10804_ _10951_/A _10804_/B vssd1 vssd1 vccd1 vccd1 _10804_/X sky130_fd_sc_hd__or2_1
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14572_ _14572_/A vssd1 vssd1 vccd1 vccd1 _18762_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_14_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11784_ _17587_/A _11784_/B vssd1 vssd1 vccd1 vccd1 _11822_/A sky130_fd_sc_hd__xnor2_2
XFILLER_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16311_ _19463_/Q _19465_/Q _19464_/Q _16435_/A vssd1 vssd1 vccd1 vccd1 _16443_/A
+ sky130_fd_sc_hd__and4_1
X_13523_ _18355_/Q _13522_/X _13529_/S vssd1 vssd1 vccd1 vccd1 _13524_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17291_ _17289_/X _17290_/X _17291_/S vssd1 vssd1 vccd1 vccd1 _17291_/X sky130_fd_sc_hd__mux2_1
X_10735_ _10823_/A _10735_/B vssd1 vssd1 vccd1 vccd1 _10735_/X sky130_fd_sc_hd__or2_1
XFILLER_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14185__S _14191_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19030_ _19320_/CLK _19030_/D vssd1 vssd1 vccd1 vccd1 _19030_/Q sky130_fd_sc_hd__dfxtp_1
X_16242_ _16242_/A vssd1 vssd1 vccd1 vccd1 _19392_/D sky130_fd_sc_hd__clkbuf_1
X_13454_ _13454_/A vssd1 vssd1 vccd1 vccd1 _18327_/D sky130_fd_sc_hd__clkbuf_1
X_10666_ _18396_/Q _18657_/Q _18556_/Q _18891_/Q _10650_/X _09380_/A vssd1 vssd1 vccd1
+ vccd1 _10667_/B sky130_fd_sc_hd__mux4_1
XFILLER_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12746__A1 hold18/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12405_ _12405_/A vssd1 vssd1 vccd1 vccd1 _17906_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_126_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16173_ _16173_/A vssd1 vssd1 vccd1 vccd1 _19360_/D sky130_fd_sc_hd__clkbuf_1
X_13385_ _15098_/A vssd1 vssd1 vccd1 vccd1 _14620_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__17134__B1 _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ _10597_/A _12461_/A vssd1 vssd1 vccd1 vccd1 _10598_/B sky130_fd_sc_hd__nor2_1
XFILLER_126_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15124_ _15124_/A vssd1 vssd1 vccd1 vccd1 _18985_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput109 _12442_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_wdata[0] sky130_fd_sc_hd__buf_2
X_12336_ _12347_/A _12316_/B _12335_/X vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__a21oi_2
XFILLER_126_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_99_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13529__S _13529_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__A3 _10771_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15055_ _18961_/Q _15054_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__mux2_1
X_12267_ _12267_/A _12267_/B vssd1 vssd1 vccd1 vccd1 _12268_/B sky130_fd_sc_hd__nand2_2
XFILLER_123_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14006_ _14006_/A vssd1 vssd1 vccd1 vccd1 _18530_/D sky130_fd_sc_hd__clkbuf_1
X_11218_ _11218_/A vssd1 vssd1 vccd1 vccd1 _11218_/Y sky130_fd_sc_hd__inv_2
X_19863_ _19865_/CLK _19863_/D vssd1 vssd1 vccd1 vccd1 _19863_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__09308__A _19708_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11557__B _17917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12198_ _12173_/A _12173_/B _12168_/A vssd1 vssd1 vccd1 vccd1 _12199_/B sky130_fd_sc_hd__a21oi_2
Xoutput80 _12123_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[18] sky130_fd_sc_hd__buf_2
XFILLER_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11049__S _11049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 _12369_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[28] sky130_fd_sc_hd__buf_2
X_11149_ _11149_/A _18484_/Q vssd1 vssd1 vccd1 vccd1 _11149_/Y sky130_fd_sc_hd__nor2_1
X_18814_ _19264_/CLK _18814_/D vssd1 vssd1 vccd1 vccd1 _18814_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19794_ _19796_/CLK _19794_/D vssd1 vssd1 vccd1 vccd1 _19794_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18745_ _19201_/CLK _18745_/D vssd1 vssd1 vccd1 vccd1 _18745_/Q sky130_fd_sc_hd__dfxtp_1
X_15957_ _13557_/X _19311_/Q _15959_/S vssd1 vssd1 vccd1 vccd1 _15958_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10907__S1 _11072_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ _14908_/A vssd1 vssd1 vccd1 vccd1 _18900_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18676_ _19296_/CLK _18676_/D vssd1 vssd1 vccd1 vccd1 _18676_/Q sky130_fd_sc_hd__dfxtp_1
X_15888_ _15888_/A vssd1 vssd1 vccd1 vccd1 _19280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_64_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17627_ _17630_/A _17630_/B _17832_/S vssd1 vssd1 vccd1 vccd1 _17627_/X sky130_fd_sc_hd__mux2_1
X_14839_ _18870_/Q _14020_/X _14843_/S vssd1 vssd1 vccd1 vccd1 _14840_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14884__A _14930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__A1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17558_ _17864_/S vssd1 vssd1 vccd1 vccd1 _17775_/S sky130_fd_sc_hd__buf_2
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16509_ _19593_/Q _19592_/Q _19594_/Q _16839_/A vssd1 vssd1 vccd1 vccd1 _16849_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__11332__S1 _10705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17489_ _17486_/X _17487_/Y _17898_/S vssd1 vssd1 vccd1 vccd1 _17489_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19228_ _19324_/CLK _19228_/D vssd1 vssd1 vccd1 vccd1 _19228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_165_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_176_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19159_ _19603_/CLK _19159_/D vssd1 vssd1 vccd1 vccd1 _19159_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18091__A _18091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14124__A _18096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_99_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17428__A1 _11612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_1_0_clock clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1_1_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_98_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15654__S _15660_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09814_ _09767_/X _09797_/X _09801_/Y _09810_/Y _09813_/X vssd1 vssd1 vccd1 vccd1
+ _09814_/X sky130_fd_sc_hd__o311a_1
XANTENNA__16100__A1 _12233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09745_ _11373_/A _09745_/B vssd1 vssd1 vccd1 vccd1 _09745_/X sky130_fd_sc_hd__or2_1
XFILLER_100_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ _09676_/A vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17170__A _17319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09888__A _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11323__S1 _09506_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16167__A1 _19359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__B1 _11288_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ _18624_/Q _18959_/Q _10520_/S vssd1 vssd1 vccd1 vccd1 _10521_/B sky130_fd_sc_hd__mux2_1
XFILLER_168_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15829__S _15837_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10451_ _18497_/Q _18992_/Q _10451_/S vssd1 vssd1 vccd1 vccd1 _10451_/X sky130_fd_sc_hd__mux2_1
XFILLER_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14733__S _14737_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11936__C1 _16109_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13170_ _15060_/A vssd1 vssd1 vccd1 vccd1 _14582_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10203__A2 _10193_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10382_ _10382_/A _10382_/B vssd1 vssd1 vccd1 vccd1 _10382_/Y sky130_fd_sc_hd__nand2_1
XFILLER_163_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _12059_/A _12059_/B _12091_/A _12120_/Y vssd1 vssd1 vccd1 vccd1 _12122_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14350__A0 _13912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _17743_/A _12140_/B vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11003_ _19175_/Q _18789_/Q _19239_/Q _18358_/Q _10940_/S _10990_/A vssd1 vssd1 vccd1
+ vccd1 _11004_/B sky130_fd_sc_hd__mux4_1
XANTENNA__18092__A1 _19844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12900__B2 _16540_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16860_ _16862_/B _16862_/C _16812_/X vssd1 vssd1 vccd1 vccd1 _16860_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10062__S1 _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15811_ _13554_/X _19246_/Q _15815_/S vssd1 vssd1 vccd1 vccd1 _15812_/A sky130_fd_sc_hd__mux2_1
XFILLER_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16791_ _19571_/Q _16791_/B vssd1 vssd1 vccd1 vccd1 _16800_/C sky130_fd_sc_hd__and2_1
XFILLER_19_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18530_ _19377_/CLK _18530_/D vssd1 vssd1 vccd1 vccd1 _18530_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15742_ _15742_/A vssd1 vssd1 vccd1 vccd1 _19215_/D sky130_fd_sc_hd__clkbuf_1
X_12954_ _19496_/Q vssd1 vssd1 vccd1 vccd1 _16551_/B sky130_fd_sc_hd__clkbuf_2
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11905_ _19402_/Q vssd1 vssd1 vccd1 vccd1 _11915_/A sky130_fd_sc_hd__buf_2
X_18461_ _19248_/CLK _18461_/D vssd1 vssd1 vccd1 vccd1 _18461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_clock clkbuf_3_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
X_15673_ _15695_/A vssd1 vssd1 vccd1 vccd1 _15682_/S sky130_fd_sc_hd__buf_6
XFILLER_34_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15602__A0 _19732_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ _15012_/A vssd1 vssd1 vccd1 vccd1 _14534_/A sky130_fd_sc_hd__clkbuf_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13812__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17659_/A vssd1 vssd1 vccd1 vccd1 _17413_/A sky130_fd_sc_hd__clkbuf_2
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14624_ input40/X _14282_/X _14293_/X _14623_/X _18107_/A vssd1 vssd1 vccd1 vccd1
+ _18205_/B sky130_fd_sc_hd__a32o_2
X_11836_ _11886_/C _11834_/Y _11835_/X vssd1 vssd1 vccd1 vccd1 _11836_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ _19305_/CLK _18392_/D vssd1 vssd1 vccd1 vccd1 _18392_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_159_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11314__S1 _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17343_ _17500_/S vssd1 vssd1 vccd1 vccd1 _17609_/A sky130_fd_sc_hd__clkbuf_2
X_14555_ _14553_/X _18757_/Q _14567_/S vssd1 vssd1 vccd1 vccd1 _14556_/A sky130_fd_sc_hd__mux2_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _19397_/Q _11768_/B vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13506_ _13506_/A vssd1 vssd1 vccd1 vccd1 _18351_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_159_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17274_ _17274_/A vssd1 vssd1 vccd1 vccd1 _17293_/S sky130_fd_sc_hd__clkbuf_2
X_10718_ _18459_/Q _19050_/Q _19212_/Q _18427_/Q _09645_/S _09541_/A vssd1 vssd1 vccd1
+ vccd1 _10719_/B sky130_fd_sc_hd__mux4_1
X_14486_ _14486_/A vssd1 vssd1 vccd1 vccd1 _18727_/D sky130_fd_sc_hd__clkbuf_1
X_11698_ _09295_/X _11698_/B vssd1 vssd1 vccd1 vccd1 _11801_/B sky130_fd_sc_hd__and2b_1
XFILLER_174_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13916__A0 _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19013_ _19109_/CLK _19013_/D vssd1 vssd1 vccd1 vccd1 _19013_/Q sky130_fd_sc_hd__dfxtp_1
X_16225_ _16225_/A vssd1 vssd1 vccd1 vccd1 _19384_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15739__S _15743_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13437_ _14998_/A _15926_/B vssd1 vssd1 vccd1 vccd1 _13494_/A sky130_fd_sc_hd__nand2_4
XFILLER_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10649_ _10649_/A _10649_/B vssd1 vssd1 vccd1 vccd1 _11453_/A sky130_fd_sc_hd__and2_1
XFILLER_10_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_127_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16156_ _15625_/X _16155_/Y _16156_/S vssd1 vssd1 vccd1 vccd1 _16156_/X sky130_fd_sc_hd__mux2_1
XFILLER_142_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13368_ _13367_/X _18313_/Q _13387_/S vssd1 vssd1 vccd1 vccd1 _13369_/A sky130_fd_sc_hd__mux2_1
XFILLER_115_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15107_ _15107_/A vssd1 vssd1 vccd1 vccd1 _18977_/D sky130_fd_sc_hd__clkbuf_1
X_12319_ _16278_/A vssd1 vssd1 vccd1 vccd1 _12319_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16087_ _12577_/B _16085_/Y _16156_/S vssd1 vssd1 vccd1 vccd1 _16087_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13299_ _16142_/B _13315_/C vssd1 vssd1 vccd1 vccd1 _13299_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_170_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15038_ _15038_/A vssd1 vssd1 vccd1 vccd1 _15038_/X sky130_fd_sc_hd__buf_2
XFILLER_130_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19846_ _19846_/CLK _19846_/D vssd1 vssd1 vccd1 vccd1 _19846_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold12_A hold12/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16989_ _16989_/A _16998_/B vssd1 vssd1 vccd1 vccd1 _16989_/X sky130_fd_sc_hd__or2_1
XFILLER_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19777_ _19780_/CLK _19777_/D vssd1 vssd1 vccd1 vccd1 _19777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_95_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _10920_/A vssd1 vssd1 vccd1 vccd1 _09531_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18728_ _19284_/CLK _18728_/D vssd1 vssd1 vccd1 vccd1 _18728_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12655__B1 _17102_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17189__A3 _12432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09461_ _10042_/A _09461_/B vssd1 vssd1 vccd1 vccd1 _09461_/X sky130_fd_sc_hd__or2_1
X_18659_ _19311_/CLK _18659_/D vssd1 vssd1 vccd1 vccd1 _18659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_92_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12670__A3 _12669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09392_ _11242_/A vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__buf_2
XFILLER_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09501__A _18642_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10647__A _10648_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__A1 _18112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13907__A0 _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15649__S _15649_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13383__A1 input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10382__A _10382_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_154_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14332__A0 _13886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13135__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11146__B1 _09469_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13693__A _13749_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_101_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09728_ _09728_/A vssd1 vssd1 vccd1 vccd1 _09844_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09659_ _09640_/X _09644_/Y _09653_/X _09657_/Y _09658_/X vssd1 vssd1 vccd1 vccd1
+ _09659_/X sky130_fd_sc_hd__o311a_2
XANTENNA__09114__C _09172_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15413__A _15459_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12657_/X _12653_/X _12669_/X _17102_/B _12696_/A vssd1 vssd1 vccd1 vccd1
+ _12670_/X sky130_fd_sc_hd__o32a_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09411__A _10873_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _18127_/A _18125_/A _11684_/C _11684_/D vssd1 vssd1 vccd1 vccd1 _11794_/A
+ sky130_fd_sc_hd__or4_4
XFILLER_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14340_ _14340_/A vssd1 vssd1 vccd1 vccd1 _18663_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ _16000_/B _11652_/A vssd1 vssd1 vccd1 vccd1 _14275_/C sky130_fd_sc_hd__nand2_1
XFILLER_168_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ _18592_/Q _18863_/Q _19087_/Q _18831_/Q _10496_/X _09710_/A vssd1 vssd1 vccd1
+ vccd1 _10503_/X sky130_fd_sc_hd__mux4_1
XFILLER_11_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14271_ _18172_/A vssd1 vssd1 vccd1 vccd1 _14290_/A sky130_fd_sc_hd__clkbuf_4
X_11483_ _11487_/S vssd1 vssd1 vccd1 vccd1 _17120_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_16010_ _16010_/A vssd1 vssd1 vccd1 vccd1 _19331_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_143_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13222_ _16896_/B _12950_/X _12951_/X _16483_/B _13221_/X vssd1 vssd1 vccd1 vccd1
+ _15586_/B sky130_fd_sc_hd__a221o_2
X_10434_ _10434_/A vssd1 vssd1 vccd1 vccd1 _10434_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13374__B2 _19359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10188__A1 _10090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10365_ _18930_/Q _18696_/Q _19378_/Q _19026_/Q _10315_/S _10229_/X vssd1 vssd1 vccd1
+ vccd1 _10366_/B sky130_fd_sc_hd__mux4_2
X_13153_ _13153_/A _13153_/B _13176_/B vssd1 vssd1 vccd1 vccd1 _13153_/X sky130_fd_sc_hd__or3_1
XFILLER_151_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12104_ _19648_/Q _12104_/B vssd1 vssd1 vccd1 vccd1 _12104_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13084_ _19753_/Q vssd1 vssd1 vccd1 vccd1 _16069_/A sky130_fd_sc_hd__clkbuf_2
X_17961_ _17961_/A vssd1 vssd1 vccd1 vccd1 _19754_/D sky130_fd_sc_hd__clkbuf_1
X_10296_ _10296_/A vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__clkbuf_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output158_A _12279_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15294__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13807__S _13809_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16912_ _19617_/Q _16912_/B _16912_/C vssd1 vssd1 vccd1 vccd1 _16914_/B sky130_fd_sc_hd__and3_1
X_19700_ _19866_/CLK _19700_/D vssd1 vssd1 vccd1 vccd1 _19700_/Q sky130_fd_sc_hd__dfxtp_1
X_12035_ _12035_/A vssd1 vssd1 vccd1 vccd1 _12035_/Y sky130_fd_sc_hd__inv_2
XFILLER_78_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11688__A1 _11683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17892_ _17673_/X _17517_/B _17891_/Y vssd1 vssd1 vccd1 vccd1 _17892_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16076__A0 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19631_ _19669_/CLK _19631_/D vssd1 vssd1 vccd1 vccd1 _19631_/Q sky130_fd_sc_hd__dfxtp_1
X_16843_ _16845_/B _16845_/C _16842_/Y vssd1 vssd1 vccd1 vccd1 _19592_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_124_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19562_ _19564_/CLK _19562_/D vssd1 vssd1 vccd1 vccd1 _19562_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13108__A _13275_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16774_ _19565_/Q _16770_/C _16773_/Y vssd1 vssd1 vccd1 vccd1 _19565_/D sky130_fd_sc_hd__o21a_1
XFILLER_168_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_92_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13986_ _18524_/Q _13985_/X _13995_/S vssd1 vssd1 vccd1 vccd1 _13987_/A sky130_fd_sc_hd__mux2_1
XFILLER_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17025__C1 _17021_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18513_ _19268_/CLK _18513_/D vssd1 vssd1 vccd1 vccd1 _18513_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15725_ _15725_/A vssd1 vssd1 vccd1 vccd1 _19207_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ _19431_/Q _12962_/A vssd1 vssd1 vccd1 vccd1 _12937_/X sky130_fd_sc_hd__or2_1
X_19493_ _19619_/CLK _19493_/D vssd1 vssd1 vccd1 vccd1 _19493_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13542__S _13545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18444_ _19197_/CLK _18444_/D vssd1 vssd1 vccd1 vccd1 _18444_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11860__A1 _19336_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15656_ _14544_/X _19177_/Q _15660_/S vssd1 vssd1 vccd1 vccd1 _15657_/A sky130_fd_sc_hd__mux2_1
X_12868_ _19743_/Q vssd1 vssd1 vccd1 vccd1 _16011_/B sky130_fd_sc_hd__clkbuf_2
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09321__A _12720_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14607_ _14607_/A vssd1 vssd1 vccd1 vccd1 _18773_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13062__A0 _19720_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18375_ _19382_/CLK _18375_/D vssd1 vssd1 vccd1 vccd1 _18375_/Q sky130_fd_sc_hd__dfxtp_1
X_11819_ _11850_/A _17245_/A vssd1 vssd1 vccd1 vccd1 _11821_/A sky130_fd_sc_hd__and2_1
XFILLER_33_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15587_ _15599_/A _18273_/Q vssd1 vssd1 vccd1 vccd1 _15587_/Y sky130_fd_sc_hd__nand2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ input1/X _12781_/X _12795_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _14996_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17326_ _17304_/X _17324_/X _17771_/A vssd1 vssd1 vccd1 vccd1 _17327_/B sky130_fd_sc_hd__mux2_1
X_14538_ _14621_/S vssd1 vssd1 vccd1 vccd1 _14551_/S sky130_fd_sc_hd__buf_2
XFILLER_119_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_105_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17257_ _17244_/X _17255_/X _17572_/S vssd1 vssd1 vccd1 vccd1 _17257_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13778__A _13835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__C1 _09448_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14469_ _14515_/S vssd1 vssd1 vccd1 vccd1 _14478_/S sky130_fd_sc_hd__buf_2
XANTENNA__09975__B _12474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_49_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16208_ _16208_/A vssd1 vssd1 vccd1 vccd1 _19376_/D sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_170_clock clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 _19329_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17188_ _17920_/A _12426_/B _17172_/Y _17173_/X _17471_/A vssd1 vssd1 vccd1 vccd1
+ _17188_/X sky130_fd_sc_hd__a41o_1
XFILLER_155_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11298__A _11298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16139_ _15608_/X _16138_/Y _16156_/S vssd1 vssd1 vccd1 vccd1 _16139_/X sky130_fd_sc_hd__mux2_1
XFILLER_170_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_102_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14865__A1 _13953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_185_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19243_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_142_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13717__S _13725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11679__A1 _11677_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11223__S0 _11219_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_97_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_97_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19829_ _19830_/CLK _19829_/D vssd1 vssd1 vccd1 vccd1 _19829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_110_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09930__S _09930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ _09513_/A vssd1 vssd1 vccd1 vccd1 _10855_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__17432__B _17432_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_92_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09444_ _18414_/Q _18675_/Q _18574_/Q _18909_/Q _09441_/X _09443_/X vssd1 vssd1 vccd1
+ vccd1 _09445_/B sky130_fd_sc_hd__mux4_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_123_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19421_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _18780_/Q vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__buf_2
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11603__A1 _11840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15379__S _15383_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_138_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19740_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09655__S0 _10785_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10150_ _10150_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _10150_/X sky130_fd_sc_hd__or2_1
XFILLER_161_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_160_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13627__S _13631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _11427_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _10083_/B sky130_fd_sc_hd__nand2_1
XFILLER_102_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14312__A _14369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09406__A _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15842__S _15848_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ _14197_/C _16622_/B vssd1 vssd1 vccd1 vccd1 _13922_/A sky130_fd_sc_hd__or2_2
XFILLER_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09840__S _09840_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13771_ _13771_/A vssd1 vssd1 vccd1 vccd1 _18450_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10983_ _10977_/A _10982_/X _09482_/A vssd1 vssd1 vccd1 vccd1 _10983_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15510_ _19715_/Q _15509_/X _15516_/S vssd1 vssd1 vccd1 vccd1 _15510_/X sky130_fd_sc_hd__mux2_1
X_12722_ hold21/A _12719_/X _17520_/S vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__mux2_1
X_16490_ _16493_/A _16493_/C _16489_/X vssd1 vssd1 vccd1 vccd1 _16490_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15441_ _15441_/A vssd1 vssd1 vccd1 vccd1 _19126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13044__A0 _13041_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ _12716_/S _12653_/B vssd1 vssd1 vccd1 vccd1 _12653_/X sky130_fd_sc_hd__or2_1
XFILLER_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18160_ _18170_/A _18160_/B vssd1 vssd1 vccd1 vccd1 _18161_/A sky130_fd_sc_hd__and2_1
X_11604_ _17438_/S _11840_/A _11668_/B vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__and3_1
X_15372_ _19096_/Q _15076_/X _15372_/S vssd1 vssd1 vccd1 vccd1 _15373_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12584_ _12584_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _12584_/Y sky130_fd_sc_hd__nor2_4
XFILLER_11_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17111_ _17168_/A _09168_/X vssd1 vssd1 vccd1 vccd1 _17130_/A sky130_fd_sc_hd__or2b_1
XANTENNA__15289__S _15289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14323_ _14369_/S vssd1 vssd1 vccd1 vccd1 _14332_/S sky130_fd_sc_hd__buf_2
XFILLER_12_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_157_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18091_ _18091_/A _18091_/B vssd1 vssd1 vccd1 vccd1 _18091_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14193__S _14195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11535_ _18742_/Q _11534_/X _11539_/S vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_50_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17042_ _19669_/Q _15487_/X _17050_/S vssd1 vssd1 vccd1 vccd1 _17043_/A sky130_fd_sc_hd__mux2_1
X_14254_ _14254_/A vssd1 vssd1 vccd1 vccd1 _18633_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11466_ _11239_/A _12443_/B _11260_/X _12442_/B _11284_/Y vssd1 vssd1 vccd1 vccd1
+ _11467_/C sky130_fd_sc_hd__a221o_1
XFILLER_165_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13205_ _13154_/X _13204_/X _13164_/X vssd1 vssd1 vccd1 vccd1 _13205_/Y sky130_fd_sc_hd__a21oi_1
X_10417_ _10406_/A _10412_/X _10414_/X _10416_/X vssd1 vssd1 vccd1 vccd1 _10417_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_152_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14185_ _18603_/Q _14033_/X _14191_/S vssd1 vssd1 vccd1 vccd1 _14186_/A sky130_fd_sc_hd__mux2_1
X_11397_ _11404_/A _11394_/X _11396_/X vssd1 vssd1 vccd1 vccd1 _11397_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_174_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16702__A _16806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13136_ _12855_/X _13130_/Y _13133_/X _13135_/X vssd1 vssd1 vccd1 vccd1 _15054_/A
+ sky130_fd_sc_hd__o31a_4
X_10348_ _10348_/A vssd1 vssd1 vccd1 vccd1 _10436_/A sky130_fd_sc_hd__clkbuf_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18993_ _19376_/CLK _18993_/D vssd1 vssd1 vccd1 vccd1 _18993_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10581__A1 _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_135_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18038__A1 _19411_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11205__S0 _11128_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10008__S1 _10056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10279_ _10479_/S vssd1 vssd1 vccd1 vccd1 _10433_/S sky130_fd_sc_hd__clkbuf_4
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ input5/X _12974_/X _12977_/X vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__a21o_2
X_17944_ _16039_/A _19779_/Q _17946_/S vssd1 vssd1 vccd1 vccd1 _17945_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14222__A _14268_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09316__A _11743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12018_ _11773_/X _12016_/X _12017_/Y _11623_/A vssd1 vssd1 vccd1 vccd1 _12018_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_94_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17875_ _17878_/A _17878_/B _17896_/S vssd1 vssd1 vccd1 vccd1 _17875_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10333__A1 _10335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15752__S _15754_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19614_ _19618_/CLK _19614_/D vssd1 vssd1 vccd1 vccd1 _19614_/Q sky130_fd_sc_hd__dfxtp_1
X_16826_ _19582_/Q _16827_/B vssd1 vssd1 vccd1 vccd1 _16828_/B sky130_fd_sc_hd__or2_1
XFILLER_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16757_ _16760_/B _16758_/C _19561_/Q vssd1 vssd1 vccd1 vccd1 _16759_/B sky130_fd_sc_hd__a21oi_1
X_19545_ _19549_/CLK _19545_/D vssd1 vssd1 vccd1 vccd1 _19545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10896__S _11071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_clock clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 _19249_/CLK sky130_fd_sc_hd__clkbuf_16
X_13969_ _14541_/A vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15708_ _14620_/X _19201_/Q _15708_/S vssd1 vssd1 vccd1 vccd1 _15709_/A sky130_fd_sc_hd__mux2_1
XFILLER_94_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16688_ _16696_/A _16688_/B _16695_/D vssd1 vssd1 vccd1 vccd1 _19538_/D sky130_fd_sc_hd__nor3_1
X_19476_ _19610_/CLK _19476_/D vssd1 vssd1 vccd1 vccd1 _19476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_clock clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_3_1_0_clock/A
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_61_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18427_ _19309_/CLK _18427_/D vssd1 vssd1 vccd1 vccd1 _18427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15639_ _15695_/A vssd1 vssd1 vccd1 vccd1 _15708_/S sky130_fd_sc_hd__buf_6
XANTENNA__10197__A _10197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09160_ _17108_/A _17165_/A vssd1 vssd1 vccd1 vccd1 _09169_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_55_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19124_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18358_ _19239_/CLK _18358_/D vssd1 vssd1 vccd1 vccd1 _18358_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09986__A _10769_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17309_ _17483_/A _17309_/B vssd1 vssd1 vccd1 vccd1 _17309_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__15500__B _18258_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09091_ _19840_/Q vssd1 vssd1 vccd1 vccd1 _09182_/B sky130_fd_sc_hd__clkbuf_1
X_18289_ _19272_/CLK _18289_/D vssd1 vssd1 vccd1 vccd1 _18289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_174_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12010__A1 _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_127_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16612__A _16714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_116_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09993_ _09993_/A _09993_/B vssd1 vssd1 vccd1 vccd1 _09993_/X sky130_fd_sc_hd__or2_1
XFILLER_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10660__A _10660_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__B1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18201__B2 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10183__S0 _09854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09427_ _10667_/A vssd1 vssd1 vccd1 vccd1 _10042_/A sky130_fd_sc_hd__buf_2
XFILLER_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16763__A1 _19562_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09896__A _10342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__C1 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09358_ _12751_/A vssd1 vssd1 vccd1 vccd1 _17795_/A sky130_fd_sc_hd__buf_2
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_138_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ _19698_/Q _09289_/B vssd1 vssd1 vccd1 vccd1 _12548_/A sky130_fd_sc_hd__and2_2
XFILLER_165_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _18622_/Q _18957_/Q _11320_/S vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__mux2_1
XFILLER_154_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_clock clkbuf_4_3_0_clock/A vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_clock/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15837__S _15837_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11251_ _19170_/Q _18784_/Q _19234_/Q _18353_/Q _09410_/A _10801_/A vssd1 vssd1 vccd1
+ vccd1 _11252_/B sky130_fd_sc_hd__mux4_1
XFILLER_162_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10202_ _09844_/X _10195_/X _10197_/X _10201_/X _09754_/A vssd1 vssd1 vccd1 vccd1
+ _10202_/X sky130_fd_sc_hd__a311o_2
X_11182_ _09431_/A _11171_/X _11175_/X _11181_/X _10949_/A vssd1 vssd1 vccd1 vccd1
+ _11182_/X sky130_fd_sc_hd__a311o_2
XFILLER_162_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10133_ _19730_/Q vssd1 vssd1 vccd1 vccd1 _10133_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15990_ _13605_/X _19326_/Q _15992_/S vssd1 vssd1 vccd1 vccd1 _15991_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12304__A2 _12476_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A io_ibus_inst[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14941_ _14941_/A vssd1 vssd1 vccd1 vccd1 _18916_/D sky130_fd_sc_hd__clkbuf_1
X_10064_ _10289_/A _10061_/X _10063_/X vssd1 vssd1 vccd1 vccd1 _10064_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17660_ _17864_/S vssd1 vssd1 vccd1 vccd1 _17842_/S sky130_fd_sc_hd__buf_2
X_14872_ _14872_/A vssd1 vssd1 vccd1 vccd1 _18884_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16611_ _19517_/Q _16607_/B _16610_/Y vssd1 vssd1 vccd1 vccd1 _19517_/D sky130_fd_sc_hd__o21a_1
X_13823_ _13274_/X _18474_/Q _13831_/S vssd1 vssd1 vccd1 vccd1 _13824_/A sky130_fd_sc_hd__mux2_1
XFILLER_78_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17591_ _17390_/A _17580_/Y _17590_/X _17542_/X vssd1 vssd1 vccd1 vccd1 _17591_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11605__S _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ _19495_/Q _19494_/Q _19493_/Q _16542_/D vssd1 vssd1 vccd1 vccd1 _16553_/D
+ sky130_fd_sc_hd__and4_1
X_19330_ _19421_/CLK _19330_/D vssd1 vssd1 vccd1 vccd1 _19330_/Q sky130_fd_sc_hd__dfxtp_2
X_13754_ _13311_/X _18444_/Q _13758_/S vssd1 vssd1 vccd1 vccd1 _13755_/A sky130_fd_sc_hd__mux2_1
X_10966_ _10965_/A _10963_/Y _10965_/Y _11160_/A vssd1 vssd1 vccd1 vccd1 _10966_/X
+ sky130_fd_sc_hd__o211a_1
X_12705_ _19688_/Q _12703_/X _12704_/X _19655_/Q vssd1 vssd1 vccd1 vccd1 _12705_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13017__A0 _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19261_ _19261_/CLK _19261_/D vssd1 vssd1 vccd1 vccd1 _19261_/Q sky130_fd_sc_hd__dfxtp_1
X_16473_ _16474_/A _16474_/C _16472_/Y vssd1 vssd1 vccd1 vccd1 _19475_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13685_ _13685_/A vssd1 vssd1 vccd1 vccd1 _18413_/D sky130_fd_sc_hd__clkbuf_1
X_10897_ _10897_/A vssd1 vssd1 vccd1 vccd1 _10897_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13820__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18212_ _18212_/A vssd1 vssd1 vccd1 vccd1 _19853_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__15601__A _15601_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15424_ _15446_/A vssd1 vssd1 vccd1 vccd1 _15433_/S sky130_fd_sc_hd__clkbuf_4
X_12636_ _12962_/A vssd1 vssd1 vccd1 vccd1 _12636_/X sky130_fd_sc_hd__clkbuf_2
X_19192_ _19382_/CLK _19192_/D vssd1 vssd1 vccd1 vccd1 _19192_/Q sky130_fd_sc_hd__dfxtp_1
X_18143_ _17125_/A _18091_/B _18142_/Y _18136_/X vssd1 vssd1 vccd1 vccd1 _19832_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15355_ _19088_/Q _15051_/X _15361_/S vssd1 vssd1 vccd1 vccd1 _15356_/A sky130_fd_sc_hd__mux2_1
XFILLER_15_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ _19681_/Q _12601_/A _12566_/X _19345_/Q vssd1 vssd1 vccd1 vccd1 _12567_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14306_ _13848_/X _18648_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _14307_/A sky130_fd_sc_hd__mux2_1
XFILLER_172_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18074_ _18121_/A vssd1 vssd1 vccd1 vccd1 _18087_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_11518_ _19842_/Q vssd1 vssd1 vccd1 vccd1 _18087_/A sky130_fd_sc_hd__buf_2
X_15286_ _15286_/A vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_144_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12498_ _17026_/S vssd1 vssd1 vccd1 vccd1 _12498_/Y sky130_fd_sc_hd__inv_2
XFILLER_172_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_171_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17025_ hold5/X _16970_/A _17024_/X _17021_/X vssd1 vssd1 vccd1 vccd1 _19662_/D sky130_fd_sc_hd__o211a_1
X_14237_ _14237_/A vssd1 vssd1 vccd1 vccd1 _18625_/D sky130_fd_sc_hd__clkbuf_1
X_11449_ _10599_/Y _11452_/B _10598_/A vssd1 vssd1 vccd1 vccd1 _11449_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_113_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17467__C1 _17466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ _14168_/A vssd1 vssd1 vccd1 vccd1 _18595_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15048__A _15080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _13119_/A _13254_/A vssd1 vssd1 vccd1 vccd1 _13167_/A sky130_fd_sc_hd__or2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14099_ _13905_/X _18565_/Q _14107_/S vssd1 vssd1 vccd1 vccd1 _14100_/A sky130_fd_sc_hd__mux2_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _19736_/CLK _18976_/D vssd1 vssd1 vccd1 vccd1 _18976_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11295__B _12457_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _19739_/Q _19771_/Q _17935_/S vssd1 vssd1 vccd1 vccd1 _17928_/A sky130_fd_sc_hd__mux2_1
XFILLER_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15482__S _15482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17858_ _17626_/X _17855_/X _17857_/Y _17532_/A vssd1 vssd1 vccd1 vccd1 _17858_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16809_ _19576_/Q _19575_/Q _19574_/Q _16809_/D vssd1 vssd1 vccd1 vccd1 _16810_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17789_ _17787_/X _17788_/Y _17855_/S vssd1 vssd1 vccd1 vccd1 _17789_/X sky130_fd_sc_hd__mux2_1
XFILLER_82_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19528_ _19543_/CLK _19528_/D vssd1 vssd1 vccd1 vccd1 _19528_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11267__C1 _11232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16745__A1 _16752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19459_ _19529_/CLK _19459_/D vssd1 vssd1 vccd1 vccd1 _19459_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18094__A _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14826__S _14832_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13730__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09212_ _09210_/X _09211_/Y _09168_/X vssd1 vssd1 vccd1 vccd1 _17176_/A sky130_fd_sc_hd__o21ai_1
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09143_ _09179_/A vssd1 vssd1 vccd1 vccd1 _17108_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__12231__A1 _19350_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14127__A _14195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_108_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_129_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10793__A1 _11335_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13966__A _14049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14561__S _14567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10390__A _10390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ _09926_/Y _10088_/A _10086_/A vssd1 vssd1 vccd1 vccd1 _11424_/A sky130_fd_sc_hd__a21o_1
XFILLER_89_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15392__S _15400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13247__A0 _19731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ _10953_/A _10810_/X _10819_/X _09448_/A vssd1 vssd1 vccd1 vccd1 _10820_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _10751_/A _10751_/B vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13470_ _13090_/X _18335_/Q _13470_/S vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__mux2_1
X_10682_ _10682_/A _10682_/B vssd1 vssd1 vccd1 vccd1 _10682_/Y sky130_fd_sc_hd__nor2_1
XFILLER_71_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_139_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _12020_/X _12482_/C _11919_/Y vssd1 vssd1 vccd1 vccd1 _17917_/B sky130_fd_sc_hd__a21o_1
XFILLER_139_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12222__B2 _12195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_166_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15140_ _15140_/A vssd1 vssd1 vccd1 vccd1 _18992_/D sky130_fd_sc_hd__clkbuf_1
X_12352_ _12314_/A _12314_/B _12348_/B _12350_/Y _12351_/Y vssd1 vssd1 vccd1 vccd1
+ _12363_/B sky130_fd_sc_hd__o311a_1
XANTENNA__11981__A0 _19784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11303_ _18590_/Q _18861_/Q _19085_/Q _18829_/Q _10764_/S _09380_/A vssd1 vssd1 vccd1
+ vccd1 _11303_/X sky130_fd_sc_hd__mux4_1
X_15071_ _18966_/Q _15070_/X _15077_/S vssd1 vssd1 vccd1 vccd1 _15072_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12283_ _17856_/A _12283_/B vssd1 vssd1 vccd1 vccd1 _12287_/A sky130_fd_sc_hd__xnor2_1
XFILLER_153_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_153_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14022_ _14022_/A vssd1 vssd1 vccd1 vccd1 _18535_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11234_ _11024_/A _11233_/X _10914_/A vssd1 vssd1 vccd1 vccd1 _11234_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18830_ _19248_/CLK _18830_/D vssd1 vssd1 vccd1 vccd1 _18830_/Q sky130_fd_sc_hd__dfxtp_1
X_11165_ _19269_/Q _19107_/Q _18516_/Q _18286_/Q _10964_/S _11030_/X vssd1 vssd1 vccd1
+ vccd1 _11165_/X sky130_fd_sc_hd__mux4_1
XFILLER_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15475__A1 _19710_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10116_ _10115_/A _10113_/Y _10115_/Y _09890_/A vssd1 vssd1 vccd1 vccd1 _10116_/X
+ sky130_fd_sc_hd__o211a_1
X_15973_ _13579_/X _19318_/Q _15981_/S vssd1 vssd1 vccd1 vccd1 _15974_/A sky130_fd_sc_hd__mux2_1
XFILLER_122_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18761_ _19054_/CLK _18761_/D vssd1 vssd1 vccd1 vccd1 _18761_/Q sky130_fd_sc_hd__dfxtp_1
X_11096_ _11465_/A vssd1 vssd1 vccd1 vccd1 _11096_/Y sky130_fd_sc_hd__inv_2
XFILLER_121_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12004__B _17214_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17712_ _17709_/A _17709_/B _17589_/X _17711_/Y vssd1 vssd1 vccd1 vccd1 _17712_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_49_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10047_ _19293_/Q _19131_/Q _18540_/Q _18310_/Q _09981_/S _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10047_/X sky130_fd_sc_hd__mux4_1
X_14924_ _18908_/Q _14039_/X _14926_/S vssd1 vssd1 vccd1 vccd1 _14925_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18692_ _19086_/CLK _18692_/D vssd1 vssd1 vccd1 vccd1 _18692_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10395__S0 _10260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17643_ _17468_/A _17640_/Y _17642_/Y vssd1 vssd1 vccd1 vccd1 _17643_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11843__B _11950_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14855_ _14855_/A vssd1 vssd1 vccd1 vccd1 _18877_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16975__A1 _12669_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13806_ _13806_/A vssd1 vssd1 vccd1 vccd1 _18466_/D sky130_fd_sc_hd__clkbuf_1
X_17574_ _17574_/A vssd1 vssd1 vccd1 vccd1 _17574_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14786_ _14786_/A vssd1 vssd1 vccd1 vccd1 _18847_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10147__S0 _09930_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ _12020_/A _12461_/A _11997_/Y vssd1 vssd1 vccd1 vccd1 _17722_/A sky130_fd_sc_hd__a21oi_4
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16525_ _19489_/Q _16521_/C _16524_/Y vssd1 vssd1 vccd1 vccd1 _19489_/D sky130_fd_sc_hd__o21a_1
X_19313_ _19375_/CLK _19313_/D vssd1 vssd1 vccd1 vccd1 _19313_/Q sky130_fd_sc_hd__dfxtp_1
X_13737_ _13737_/A vssd1 vssd1 vccd1 vccd1 _18436_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__16727__A1 _19551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14646__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ _10949_/A _10949_/B _10949_/C vssd1 vssd1 vccd1 vccd1 _10949_/X sky130_fd_sc_hd__or3_2
XANTENNA__12955__A _13391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16456_ _16458_/A _16458_/C _16446_/X vssd1 vssd1 vccd1 vccd1 _16456_/Y sky130_fd_sc_hd__a21oi_1
X_19244_ _19247_/CLK _19244_/D vssd1 vssd1 vccd1 vccd1 _19244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13668_ _13668_/A vssd1 vssd1 vccd1 vccd1 _18405_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15407_ _19111_/Q _15022_/X _15411_/S vssd1 vssd1 vccd1 vccd1 _15408_/A sky130_fd_sc_hd__mux2_1
X_12619_ _12619_/A _16937_/C vssd1 vssd1 vccd1 vccd1 _12716_/S sky130_fd_sc_hd__nand2_2
XFILLER_129_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19175_ _19239_/CLK _19175_/D vssd1 vssd1 vccd1 vccd1 _19175_/Q sky130_fd_sc_hd__dfxtp_1
X_16387_ _19445_/Q _19444_/Q _16387_/C vssd1 vssd1 vccd1 vccd1 _16389_/B sky130_fd_sc_hd__and3_1
XFILLER_129_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13599_ _15083_/A vssd1 vssd1 vccd1 vccd1 _13599_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18126_ _09267_/B _18120_/X _18125_/X _18123_/X vssd1 vssd1 vccd1 vccd1 _19825_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15338_ _15338_/A vssd1 vssd1 vccd1 vccd1 _19080_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_117_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11972__B1 _16114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18057_ _19798_/Q _19419_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18058_/A sky130_fd_sc_hd__mux2_1
X_15269_ _15315_/S vssd1 vssd1 vccd1 vccd1 _15278_/S sky130_fd_sc_hd__buf_2
XANTENNA__10870__S1 _11174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17008_ _18097_/A vssd1 vssd1 vccd1 vccd1 _17008_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__09917__B1 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09830_ _09830_/A vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_99_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09761_/A vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__clkbuf_2
X_18959_ _19088_/CLK _18959_/D vssd1 vssd1 vccd1 vccd1 _18959_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18089__A _18089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13725__S _13725_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _10236_/A vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_172_clock_A clkbuf_4_3_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09504__A _10965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13229__A0 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16966__A1 _15515_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_148_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13026__A _13387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12584__B _12606_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_148_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_157_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17679__C1 _17466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09126_ _13114_/A vssd1 vssd1 vccd1 vccd1 _13132_/A sky130_fd_sc_hd__clkinv_2
XFILLER_163_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10766__A1 _09671_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15387__S _15387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_135_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11928__B _17201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11715__B1 _11674_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_150_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_150_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10613__S1 _09419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09959_ _18601_/Q _18872_/Q _19096_/Q _18840_/Q _10217_/S _09891_/A vssd1 vssd1 vccd1
+ vccd1 _09959_/X sky130_fd_sc_hd__mux4_1
XFILLER_106_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12970_ _16039_/A _12971_/B vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__nor2_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10377__S0 _10260_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09414__A _10764_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _19855_/Q _11920_/X _11943_/A vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__mux2_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11494__A2 _11481_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15850__S _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _16282_/A _18213_/B vssd1 vssd1 vccd1 vccd1 _14641_/A sky130_fd_sc_hd__and2_2
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _11791_/A _11790_/B _11824_/A _11851_/Y vssd1 vssd1 vccd1 vccd1 _11852_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _19178_/Q _18792_/Q _19242_/Q _18361_/Q _10872_/S _10802_/X vssd1 vssd1 vccd1
+ vccd1 _10804_/B sky130_fd_sc_hd__mux4_1
XFILLER_72_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _14569_/X _18762_/Q _14583_/S vssd1 vssd1 vccd1 vccd1 _14572_/A sky130_fd_sc_hd__mux2_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11842_/A _11842_/C _12050_/A vssd1 vssd1 vccd1 vccd1 _11784_/B sky130_fd_sc_hd__a21oi_1
XFILLER_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16310_ _19461_/Q _19460_/Q _19462_/Q _16426_/A vssd1 vssd1 vccd1 vccd1 _16435_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_159_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13522_ _15006_/A vssd1 vssd1 vccd1 vccd1 _13522_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17290_ _12358_/A _17492_/B _17293_/S vssd1 vssd1 vccd1 vccd1 _17290_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10734_ _18395_/Q _18656_/Q _18555_/Q _18890_/Q _10824_/S _09705_/A vssd1 vssd1 vccd1
+ vccd1 _10735_/B sky130_fd_sc_hd__mux4_1
XFILLER_41_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16241_ _16282_/A _16241_/B vssd1 vssd1 vccd1 vccd1 _16242_/A sky130_fd_sc_hd__and2_1
XFILLER_13_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13453_ _12924_/X _18327_/Q _13459_/S vssd1 vssd1 vccd1 vccd1 _13454_/A sky130_fd_sc_hd__mux2_1
X_10665_ _11313_/A _10665_/B vssd1 vssd1 vccd1 vccd1 _10665_/X sky130_fd_sc_hd__or2_1
X_12404_ _19801_/Q _11413_/A _12404_/S vssd1 vssd1 vccd1 vccd1 _12405_/A sky130_fd_sc_hd__mux2_4
XFILLER_173_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16172_ _13509_/X _19360_/Q _16180_/S vssd1 vssd1 vccd1 vccd1 _16173_/A sky130_fd_sc_hd__mux2_1
XANTENNA__17134__A1 _17114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13384_ _13051_/X _13382_/X _13383_/X vssd1 vssd1 vccd1 vccd1 _15098_/A sky130_fd_sc_hd__o21a_1
XANTENNA__17134__B2 _15612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10757__A1 _19113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10596_ _10597_/A _12461_/A vssd1 vssd1 vccd1 vccd1 _10598_/A sky130_fd_sc_hd__and2_1
XFILLER_126_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15123_ _18985_/Q _15028_/X _15123_/S vssd1 vssd1 vccd1 vccd1 _15124_/A sky130_fd_sc_hd__mux2_1
X_12335_ _12310_/A _17867_/B vssd1 vssd1 vccd1 vccd1 _12335_/X sky130_fd_sc_hd__and2b_1
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15054_ _15054_/A vssd1 vssd1 vccd1 vccd1 _15054_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_114_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12266_ _12223_/A _12224_/A _12223_/B _12249_/B _12221_/A vssd1 vssd1 vccd1 vccd1
+ _12267_/B sky130_fd_sc_hd__a311o_1
X_14005_ _18530_/Q _14004_/X _14011_/S vssd1 vssd1 vccd1 vccd1 _14006_/A sky130_fd_sc_hd__mux2_1
X_11217_ _18482_/Q _18977_/Q _18641_/Q vssd1 vssd1 vccd1 vccd1 _11218_/A sky130_fd_sc_hd__mux2_1
X_19862_ _19865_/CLK _19862_/D vssd1 vssd1 vccd1 vccd1 _19862_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_150_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12197_ _12223_/A _12197_/B vssd1 vssd1 vccd1 vccd1 _12199_/A sky130_fd_sc_hd__nand2_2
XFILLER_150_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11182__A1 _09431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput81 _12149_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[19] sky130_fd_sc_hd__buf_2
Xoutput92 _12389_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[29] sky130_fd_sc_hd__buf_2
X_18813_ _19389_/CLK _18813_/D vssd1 vssd1 vccd1 vccd1 _18813_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11148_ _18979_/Q vssd1 vssd1 vccd1 vccd1 _11148_/Y sky130_fd_sc_hd__inv_2
XFILLER_110_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19793_ _19793_/CLK _19793_/D vssd1 vssd1 vccd1 vccd1 _19793_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13545__S _13545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18744_ _19799_/CLK _18744_/D vssd1 vssd1 vccd1 vccd1 _18744_/Q sky130_fd_sc_hd__dfxtp_2
X_11079_ _18389_/Q _18650_/Q _18549_/Q _18884_/Q _09496_/A _11030_/X vssd1 vssd1 vccd1
+ vccd1 _11080_/B sky130_fd_sc_hd__mux4_1
X_15956_ _15956_/A vssd1 vssd1 vccd1 vccd1 _19310_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14907_ _18900_/Q _14013_/X _14915_/S vssd1 vssd1 vccd1 vccd1 _14908_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16948__A1 _13418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12682__A1 _19584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15887_ _19280_/Q _14566_/A _15887_/S vssd1 vssd1 vccd1 vccd1 _15888_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18675_ _19324_/CLK _18675_/D vssd1 vssd1 vccd1 vccd1 _18675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17626_ _17626_/A vssd1 vssd1 vccd1 vccd1 _17626_/X sky130_fd_sc_hd__clkbuf_2
X_14838_ _14838_/A vssd1 vssd1 vccd1 vccd1 _18869_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15620__A1 _15612_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14769_ _14769_/A vssd1 vssd1 vccd1 vccd1 _18839_/D sky130_fd_sc_hd__clkbuf_1
X_17557_ _17479_/X _17655_/B _17483_/X vssd1 vssd1 vccd1 vccd1 _17871_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__14376__S _14384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18165__A3 _18066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16508_ _19588_/Q _19589_/Q _19591_/Q _19590_/Q vssd1 vssd1 vccd1 vccd1 _16839_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_108_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17488_ _17584_/A vssd1 vssd1 vccd1 vccd1 _17898_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_149_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_149_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19227_ _19291_/CLK _19227_/D vssd1 vssd1 vccd1 vccd1 _19227_/Q sky130_fd_sc_hd__dfxtp_1
X_16439_ _16440_/A _16440_/C _16438_/Y vssd1 vssd1 vccd1 vccd1 _19463_/D sky130_fd_sc_hd__o21a_1
XFILLER_158_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_119_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_158_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19158_ _19162_/CLK _19158_/D vssd1 vssd1 vccd1 vccd1 _19158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18091__B _18091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10748__B2 _19717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18109_ _18109_/A _18128_/B vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__nand2_1
X_19089_ _19089_/CLK _19089_/D vssd1 vssd1 vccd1 vccd1 _19089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_117_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14124__B _14860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15935__S _15937_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _09813_/A vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__buf_2
XFILLER_99_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16100__A2 _15568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_140_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09744_ _19198_/Q _18812_/Q _19262_/Q _18381_/Q _11374_/S _09687_/A vssd1 vssd1 vccd1
+ vccd1 _09745_/B sky130_fd_sc_hd__mux4_1
XFILLER_101_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09675_ _09927_/A vssd1 vssd1 vccd1 vccd1 _09676_/A sky130_fd_sc_hd__buf_4
XFILLER_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18156__A3 _18066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__A1 _10895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10987__B2 _12449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11004__A _11171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_148_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10450_ _18625_/Q _18960_/Q _10450_/S vssd1 vssd1 vccd1 vccd1 _10450_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09109_ _19841_/Q vssd1 vssd1 vccd1 vccd1 _09182_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10381_ _18627_/Q _18962_/Q _10381_/S vssd1 vssd1 vccd1 vccd1 _10382_/B sky130_fd_sc_hd__mux2_1
XANTENNA__10203__A3 _10202_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12120_ _12120_/A _12120_/B vssd1 vssd1 vccd1 vccd1 _12120_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12051_ _12140_/A vssd1 vssd1 vccd1 vccd1 _17743_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ _11195_/A vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_120_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18092__A2 _12694_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10989__S _11241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15810_ _15810_/A vssd1 vssd1 vccd1 vccd1 _19245_/D sky130_fd_sc_hd__clkbuf_1
X_16790_ _19570_/Q _16790_/B _16790_/C vssd1 vssd1 vccd1 vccd1 _16791_/B sky130_fd_sc_hd__and3_1
XFILLER_120_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15741_ _13557_/X _19215_/Q _15743_/S vssd1 vssd1 vccd1 vccd1 _15742_/A sky130_fd_sc_hd__mux2_1
X_12953_ _12953_/A vssd1 vssd1 vccd1 vccd1 _12953_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11904_ _11904_/A vssd1 vssd1 vccd1 vccd1 _11904_/Y sky130_fd_sc_hd__inv_2
XANTENNA__10675__B1 _09374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _19309_/CLK _18460_/D vssd1 vssd1 vccd1 vccd1 _18460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15672_ _15672_/A vssd1 vssd1 vccd1 vccd1 _19184_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ input27/X _12781_/X _12883_/X _12798_/X vssd1 vssd1 vccd1 vccd1 _15012_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15602__A1 _15600_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14623_ _14623_/A vssd1 vssd1 vccd1 vccd1 _14623_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17907_/A _17407_/A _17724_/A _17410_/X vssd1 vssd1 vccd1 vccd1 _17411_/X
+ sky130_fd_sc_hd__o211a_1
X_11835_ _11887_/A vssd1 vssd1 vccd1 vccd1 _11835_/X sky130_fd_sc_hd__clkbuf_2
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _19308_/CLK _18391_/D vssd1 vssd1 vccd1 vccd1 _18391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output103_A _09096_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10427__B1 _09821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17342_ _17575_/S vssd1 vssd1 vccd1 vccd1 _17500_/S sky130_fd_sc_hd__clkbuf_2
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14621_/S vssd1 vssd1 vccd1 vccd1 _14567_/S sky130_fd_sc_hd__buf_2
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ _11859_/A vssd1 vssd1 vccd1 vccd1 _11766_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13505_ _13367_/X _18351_/Q _13507_/S vssd1 vssd1 vccd1 vccd1 _13506_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17273_ _17270_/X _17365_/B _17291_/S vssd1 vssd1 vccd1 vccd1 _17273_/X sky130_fd_sc_hd__mux2_1
X_10717_ _10773_/A _10717_/B vssd1 vssd1 vccd1 vccd1 _10717_/Y sky130_fd_sc_hd__nor2_1
X_14485_ _13896_/X _18727_/Q _14489_/S vssd1 vssd1 vccd1 vccd1 _14486_/A sky130_fd_sc_hd__mux2_1
X_11697_ _13430_/A _11551_/B _11695_/Y _11696_/Y vssd1 vssd1 vccd1 vccd1 _11706_/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA__14924__S _14926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16705__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16224_ _13592_/X _19384_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16225_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19012_ _19012_/CLK _19012_/D vssd1 vssd1 vccd1 vccd1 _19012_/Q sky130_fd_sc_hd__dfxtp_1
X_13436_ _18096_/A _14371_/B _14197_/C vssd1 vssd1 vccd1 vccd1 _15926_/B sky130_fd_sc_hd__nor3_4
XFILLER_174_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10648_ _10648_/A _12459_/A vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__or2_1
XFILLER_173_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_155_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16155_ _16159_/A _16159_/C vssd1 vssd1 vccd1 vccd1 _16155_/Y sky130_fd_sc_hd__xnor2_1
X_13367_ _14617_/A vssd1 vssd1 vccd1 vccd1 _13367_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_154_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10753__A _11309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10579_ _10579_/A vssd1 vssd1 vccd1 vccd1 _10579_/X sky130_fd_sc_hd__buf_4
XFILLER_170_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15106_ _18977_/Q _15003_/X _15112_/S vssd1 vssd1 vccd1 vccd1 _15107_/A sky130_fd_sc_hd__mux2_1
X_12318_ _19418_/Q vssd1 vssd1 vccd1 vccd1 _12321_/A sky130_fd_sc_hd__buf_2
X_16086_ _16086_/A vssd1 vssd1 vccd1 vccd1 _16156_/S sky130_fd_sc_hd__clkbuf_2
X_13298_ _19766_/Q vssd1 vssd1 vccd1 vccd1 _16142_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_142_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _15037_/A vssd1 vssd1 vccd1 vccd1 _18955_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_130_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12249_ _12348_/A _12249_/B vssd1 vssd1 vccd1 vccd1 _12251_/A sky130_fd_sc_hd__nor2_1
XFILLER_123_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10589__S0 _10017_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19845_ _19845_/CLK _19845_/D vssd1 vssd1 vccd1 vccd1 _19845_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_96_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10899__S _10964_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16094__A1 _12233_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A _18138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19776_ _19779_/CLK _19776_/D vssd1 vssd1 vccd1 vccd1 _19776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16988_ _12577_/B _16983_/X _16987_/X _16981_/X vssd1 vssd1 vccd1 vccd1 _19648_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_111_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18727_ _19377_/CLK _18727_/D vssd1 vssd1 vccd1 vccd1 _18727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_45_clock_A clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12655__A1 _16929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15939_ _15996_/S vssd1 vssd1 vccd1 vccd1 _15948_/S sky130_fd_sc_hd__buf_2
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13852__A0 _13851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12655__B2 _19584_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09460_ _19295_/Q _19133_/Q _18542_/Q _18312_/Q _09441_/X _10031_/A vssd1 vssd1 vccd1
+ vccd1 _09461_/B sky130_fd_sc_hd__mux4_1
X_18658_ _19310_/CLK _18658_/D vssd1 vssd1 vccd1 vccd1 _18658_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17594__A1 _11796_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10761__S0 _10660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17609_ _17609_/A _17609_/B vssd1 vssd1 vccd1 vccd1 _17609_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09391_ _18780_/Q vssd1 vssd1 vccd1 vccd1 _11242_/A sky130_fd_sc_hd__inv_2
X_18589_ _19086_/CLK _18589_/D vssd1 vssd1 vccd1 vccd1 _18589_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10513__S0 _09980_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10647__B _12459_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_138_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10139__S _10185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_164_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16306__C1 _16280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17649__A2 _17648_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_161_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_133_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15665__S _15671_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11146__A1 _09366_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11146__B2 _19709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_101_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17282__A0 _17856_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17821__A2 _17819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_170_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09727_ _09727_/A vssd1 vssd1 vccd1 vccd1 _09728_/A sky130_fd_sc_hd__buf_2
XFILLER_101_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13843__A0 _13837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09658_ _09658_/A vssd1 vssd1 vccd1 vccd1 _09658_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10752__S0 _10729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_169_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _09589_/A _09589_/B vssd1 vssd1 vccd1 vccd1 _09589_/X sky130_fd_sc_hd__and2_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11620_/A _18087_/A _17115_/A vssd1 vssd1 vccd1 vccd1 _11684_/D sky130_fd_sc_hd__or3b_1
XANTENNA__13214__A _13234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17337__A1 _17305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10504__S0 _09980_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _11551_/A _11551_/B vssd1 vssd1 vccd1 vccd1 _16000_/B sky130_fd_sc_hd__nor2_8
XFILLER_169_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14744__S _14748_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10502_ _10312_/A _10499_/X _10501_/X vssd1 vssd1 vccd1 vccd1 _10502_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09838__S _09840_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14270_ _17102_/A vssd1 vssd1 vccd1 vccd1 _18172_/A sky130_fd_sc_hd__buf_2
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11482_ _11491_/B _11646_/C _11481_/X vssd1 vssd1 vccd1 vccd1 _11495_/A sky130_fd_sc_hd__or3b_1
XFILLER_11_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13221_ _19542_/Q _12952_/X _12953_/X _19510_/Q _13220_/X vssd1 vssd1 vccd1 vccd1
+ _13221_/X sky130_fd_sc_hd__a221o_1
XANTENNA__13374__A2 _12603_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10433_ _18498_/Q _18993_/Q _10433_/S vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__mux2_1
XFILLER_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11669__A _11840_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input64_A io_ibus_inst[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ _19757_/Q _19758_/Q _13152_/C vssd1 vssd1 vccd1 vccd1 _13176_/B sky130_fd_sc_hd__and3_1
X_10364_ _10357_/X _10359_/X _10361_/X _10363_/X _09753_/A vssd1 vssd1 vccd1 vccd1
+ _10364_/X sky130_fd_sc_hd__a221o_4
XFILLER_151_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10593__C1 _09572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ _19345_/Q _11859_/X _12037_/X _12101_/X _12102_/X vssd1 vssd1 vccd1 vccd1
+ _12103_/X sky130_fd_sc_hd__o221a_1
XFILLER_97_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ _19753_/Q _13083_/B vssd1 vssd1 vccd1 vccd1 _13111_/C sky130_fd_sc_hd__and2_1
X_17960_ _13095_/A _19786_/Q _17968_/S vssd1 vssd1 vccd1 vccd1 _17961_/A sky130_fd_sc_hd__mux2_1
X_10295_ _19286_/Q _19124_/Q _18533_/Q _18303_/Q _10274_/X _10263_/X vssd1 vssd1 vccd1
+ vccd1 _10295_/X sky130_fd_sc_hd__mux4_1
XFILLER_151_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16911_ _16912_/B _16912_/C _16910_/Y vssd1 vssd1 vccd1 vccd1 _19616_/D sky130_fd_sc_hd__o21a_1
X_12034_ _12034_/A _12034_/B vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__xnor2_2
XFILLER_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17891_ _17888_/X _17890_/X _17542_/X vssd1 vssd1 vccd1 vccd1 _17891_/Y sky130_fd_sc_hd__a21oi_1
X_19630_ _19663_/CLK _19630_/D vssd1 vssd1 vccd1 vccd1 _19630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_144_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16842_ _16845_/B _16845_/C _16812_/X vssd1 vssd1 vccd1 vccd1 _16842_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_93_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19561_ _19564_/CLK _19561_/D vssd1 vssd1 vccd1 vccd1 _19561_/Q sky130_fd_sc_hd__dfxtp_2
X_16773_ _16840_/A _16782_/D vssd1 vssd1 vccd1 vccd1 _16773_/Y sky130_fd_sc_hd__nor2_1
X_13985_ _14557_/A vssd1 vssd1 vccd1 vccd1 _13985_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__13823__S _13831_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18512_ _19391_/CLK _18512_/D vssd1 vssd1 vccd1 vccd1 _18512_/Q sky130_fd_sc_hd__dfxtp_1
X_12936_ _16937_/A _19638_/Q _16937_/B _12935_/X vssd1 vssd1 vccd1 vccd1 _12936_/X
+ sky130_fd_sc_hd__a31o_2
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15724_ _13531_/X _19207_/Q _15732_/S vssd1 vssd1 vccd1 vccd1 _15725_/A sky130_fd_sc_hd__mux2_1
X_19492_ _19619_/CLK _19492_/D vssd1 vssd1 vccd1 vccd1 _19492_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _19387_/CLK _18443_/D vssd1 vssd1 vccd1 vccd1 _18443_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15655_ _15655_/A vssd1 vssd1 vccd1 vccd1 _19176_/D sky130_fd_sc_hd__clkbuf_1
X_12867_ _12867_/A vssd1 vssd1 vccd1 vccd1 _18286_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11818_ _19778_/Q _10895_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _17245_/A sky130_fd_sc_hd__mux2_4
X_14606_ _14605_/X _18773_/Q _14615_/S vssd1 vssd1 vccd1 vccd1 _14607_/A sky130_fd_sc_hd__mux2_1
X_18374_ _19502_/CLK _18374_/D vssd1 vssd1 vccd1 vccd1 _18374_/Q sky130_fd_sc_hd__dfxtp_1
X_15586_ _18273_/Q _15586_/B vssd1 vssd1 vccd1 vccd1 _15586_/X sky130_fd_sc_hd__or2_1
XANTENNA__13062__A1 _15534_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ _12976_/A vssd1 vssd1 vccd1 vccd1 _12798_/X sky130_fd_sc_hd__buf_4
XFILLER_15_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14537_ _14537_/A vssd1 vssd1 vccd1 vccd1 _14537_/X sky130_fd_sc_hd__clkbuf_2
X_17325_ _17432_/A _17432_/B _17190_/A vssd1 vssd1 vccd1 vccd1 _17771_/A sky130_fd_sc_hd__or3b_1
X_11749_ _11749_/A _11749_/B vssd1 vssd1 vccd1 vccd1 _11750_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14654__S _14654_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_105_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14468_ _14468_/A vssd1 vssd1 vccd1 vccd1 _18719_/D sky130_fd_sc_hd__clkbuf_1
X_17256_ _17256_/A vssd1 vssd1 vccd1 vccd1 _17572_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_128_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13419_ _13419_/A _13419_/B vssd1 vssd1 vccd1 vccd1 _13419_/Y sky130_fd_sc_hd__nand2_1
X_16207_ _13567_/X _19376_/Q _16213_/S vssd1 vssd1 vccd1 vccd1 _16208_/A sky130_fd_sc_hd__mux2_1
X_17187_ _17387_/B _17404_/C vssd1 vssd1 vccd1 vccd1 _17471_/A sky130_fd_sc_hd__or2_1
XFILLER_143_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14399_ _14399_/A vssd1 vssd1 vccd1 vccd1 _18688_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_127_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11376__A1 _10138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16138_ _16142_/A _16142_/C vssd1 vssd1 vccd1 vccd1 _16138_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_115_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_143_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16069_ _16069_/A _16073_/C vssd1 vssd1 vccd1 vccd1 _16069_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_130_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_130_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16067__A1 _19341_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17264__A0 _17790_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19828_ _19828_/CLK _19828_/D vssd1 vssd1 vccd1 vccd1 _19828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10982__S0 _09625_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12628__A1 _16929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19759_ _19759_/CLK _19759_/D vssd1 vssd1 vccd1 vccd1 _19759_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18097__A _18097_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09512_ _09512_/A vssd1 vssd1 vccd1 vccd1 _09513_/A sky130_fd_sc_hd__buf_2
XFILLER_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11300__A1 _09394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10734__S0 _10824_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11761__B _17250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__A _09512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ _09443_/A vssd1 vssd1 vccd1 vccd1 _09443_/X sky130_fd_sc_hd__buf_4
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09374_ _09374_/A vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14564__S _14567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09655__S1 _10586_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15502__A0 _19714_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10080_ _10080_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10327__C1 _09857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_99_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12113__A _17779_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_101_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13816__A0 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15424__A _15446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__A _17696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13770_ _12828_/X _18450_/Q _13776_/S vssd1 vssd1 vccd1 vccd1 _13771_/A sky130_fd_sc_hd__mux2_1
X_10982_ _19272_/Q _19110_/Q _18519_/Q _18289_/Q _09625_/A _10910_/X vssd1 vssd1 vccd1
+ vccd1 _10982_/X sky130_fd_sc_hd__mux4_1
XFILLER_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15569__A0 _19726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12721_ _17937_/A vssd1 vssd1 vccd1 vccd1 _17520_/S sky130_fd_sc_hd__buf_2
XFILLER_83_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15440_ _19126_/Q _15070_/X _15444_/S vssd1 vssd1 vccd1 vccd1 _15441_/A sky130_fd_sc_hd__mux2_1
X_12652_ _15632_/S _12652_/B vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09141__B _19864_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11603_ _11840_/A _17207_/A _17438_/S vssd1 vssd1 vccd1 vccd1 _11607_/A sky130_fd_sc_hd__a21oi_1
XFILLER_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15371_ _15371_/A vssd1 vssd1 vccd1 vccd1 _19095_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_168_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _12782_/A vssd1 vssd1 vccd1 vccd1 _12583_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14474__S _14478_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_156_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ _14322_/A vssd1 vssd1 vccd1 vccd1 _18655_/D sky130_fd_sc_hd__clkbuf_1
X_17110_ _17110_/A _17169_/B vssd1 vssd1 vccd1 vccd1 _17131_/C sky130_fd_sc_hd__or2_1
X_18090_ _19843_/Q _12694_/X _18089_/Y _18084_/X vssd1 vssd1 vccd1 vccd1 _19811_/D
+ sky130_fd_sc_hd__o211a_1
X_11534_ _11721_/S _17145_/C _11514_/X _11533_/X vssd1 vssd1 vccd1 vccd1 _11534_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_157_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11070__A3 _11069_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17041_ _17098_/S vssd1 vssd1 vccd1 vccd1 _17050_/S sky130_fd_sc_hd__clkbuf_4
X_14253_ _18633_/Q _14026_/X _14253_/S vssd1 vssd1 vccd1 vccd1 _14254_/A sky130_fd_sc_hd__mux2_1
XFILLER_8_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11465_ _11465_/A _11465_/B _11465_/C _11465_/D vssd1 vssd1 vccd1 vccd1 _11470_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_143_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_109_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13204_ _19728_/Q _15580_/B _13306_/A vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__mux2_1
XFILLER_87_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _09674_/A _10415_/X _10250_/A vssd1 vssd1 vccd1 vccd1 _10416_/X sky130_fd_sc_hd__a21o_1
XFILLER_125_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14184_ _14184_/A vssd1 vssd1 vccd1 vccd1 _18602_/D sky130_fd_sc_hd__clkbuf_1
X_11396_ _11402_/A _11395_/X _09767_/X vssd1 vssd1 vccd1 vccd1 _11396_/X sky130_fd_sc_hd__o21a_1
XANTENNA__16297__A1 _19416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13818__S _13820_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13135_ input9/X _13134_/X _13120_/X vssd1 vssd1 vccd1 vccd1 _13135_/X sky130_fd_sc_hd__a21o_1
XFILLER_174_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10347_ _10347_/A vssd1 vssd1 vccd1 vccd1 _10348_/A sky130_fd_sc_hd__buf_2
XFILLER_151_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18992_ _19120_/CLK _18992_/D vssd1 vssd1 vccd1 vccd1 _18992_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11846__B _17198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17943_ _17943_/A vssd1 vssd1 vccd1 vccd1 _19746_/D sky130_fd_sc_hd__clkbuf_1
X_13066_ _13153_/A _13062_/X _13065_/X vssd1 vssd1 vccd1 vccd1 _13066_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__10318__C1 _09728_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10278_ _10531_/A vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__buf_2
XANTENNA__11205__S1 _11177_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__A1 _15998_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16049__A1 _19338_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10750__B _12455_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _16978_/A _12044_/C vssd1 vssd1 vccd1 vccd1 _12017_/Y sky130_fd_sc_hd__nand2_1
XFILLER_120_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17874_ _17874_/A vssd1 vssd1 vccd1 vccd1 _19733_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_66_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17797__A1 _19726_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19613_ _19618_/CLK _19613_/D vssd1 vssd1 vccd1 vccd1 _19613_/Q sky130_fd_sc_hd__dfxtp_1
X_16825_ _16838_/A _16825_/B _16827_/B vssd1 vssd1 vccd1 vccd1 _19581_/D sky130_fd_sc_hd__nor3_1
XFILLER_94_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19544_ _19549_/CLK _19544_/D vssd1 vssd1 vccd1 vccd1 _19544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16756_ _16760_/B _16758_/C _16755_/Y vssd1 vssd1 vccd1 vccd1 _19560_/D sky130_fd_sc_hd__o21a_1
XFILLER_93_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13968_ _13968_/A vssd1 vssd1 vccd1 vccd1 _18518_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__S0 _09645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09332__A _19855_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15707_ _15707_/A vssd1 vssd1 vccd1 vccd1 _19200_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_80_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12919_ _19594_/Q _12560_/X _12562_/X _19462_/Q _12918_/X vssd1 vssd1 vccd1 vccd1
+ _15493_/B sky130_fd_sc_hd__a221o_2
X_19475_ _19610_/CLK _19475_/D vssd1 vssd1 vccd1 vccd1 _19475_/Q sky130_fd_sc_hd__dfxtp_1
X_16687_ _19538_/Q _19537_/Q _19536_/Q _16687_/D vssd1 vssd1 vccd1 vccd1 _16695_/D
+ sky130_fd_sc_hd__and4_1
X_13899_ _14579_/A vssd1 vssd1 vccd1 vccd1 _13899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18426_ _19180_/CLK _18426_/D vssd1 vssd1 vccd1 vccd1 _18426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15638_ _15926_/A _15782_/B vssd1 vssd1 vccd1 vccd1 _15695_/A sky130_fd_sc_hd__nand2_4
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13035__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13789__A _13835_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18357_ _19302_/CLK _18357_/D vssd1 vssd1 vccd1 vccd1 _18357_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14384__S _14384_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15569_ _19726_/Q _15568_/X _15569_/S vssd1 vssd1 vccd1 vccd1 _15569_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11141__S0 _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16165__A _19770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_159_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_148_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17308_ _17404_/A _11842_/A _17234_/Y vssd1 vssd1 vccd1 vccd1 _17309_/B sky130_fd_sc_hd__o21ai_1
X_09090_ _19847_/Q vssd1 vssd1 vccd1 vccd1 _09186_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_174_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18288_ _19271_/CLK _18288_/D vssd1 vssd1 vccd1 vccd1 _18288_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15732__A0 _13544_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239_ _17239_/A vssd1 vssd1 vccd1 vccd1 _17463_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_174_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_116_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13728__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09992_ _19196_/Q _18810_/Q _19260_/Q _18379_/Q _09850_/A _09977_/X vssd1 vssd1 vccd1
+ vccd1 _09993_/B sky130_fd_sc_hd__mux4_1
XFILLER_171_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09507__A _09507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12849__B2 _12781_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10955__S0 _11196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10183__S1 _09676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09426_ _11305_/A vssd1 vssd1 vccd1 vccd1 _10667_/A sky130_fd_sc_hd__buf_2
XFILLER_53_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09357_ _17102_/A _17133_/B vssd1 vssd1 vccd1 vccd1 _12751_/A sky130_fd_sc_hd__nand2_4
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12785__B1 _12704_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09288_ _19820_/Q _19818_/Q _09288_/C vssd1 vssd1 vccd1 vccd1 _16624_/A sky130_fd_sc_hd__or3_2
XFILLER_21_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_167_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11012__A _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11250_ _10943_/X _11245_/X _11249_/X _11001_/A vssd1 vssd1 vccd1 vccd1 _11250_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_106_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10201_ _10195_/A _10198_/X _10200_/X _09740_/A vssd1 vssd1 vccd1 vccd1 _10201_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17768__A_N _17215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11181_ _11188_/A _11178_/X _11180_/X _10883_/X vssd1 vssd1 vccd1 vccd1 _11181_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__16014__S _16024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14323__A _14369_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10851__A _10962_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_79_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_161_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10132_ _10125_/Y _10127_/Y _10129_/Y _10131_/Y _09831_/X vssd1 vssd1 vccd1 vccd1
+ _10132_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09417__A _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14940_ _18916_/Q vssd1 vssd1 vccd1 vccd1 _14941_/A sky130_fd_sc_hd__clkbuf_1
X_10063_ _10680_/A _10062_/X _09640_/X vssd1 vssd1 vccd1 vccd1 _10063_/X sky130_fd_sc_hd__o21a_1
XFILLER_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10946__S0 _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input27_A io_dbus_rdata[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ _18884_/Q _13962_/X _14871_/S vssd1 vssd1 vccd1 vccd1 _14872_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16610_ _16610_/A _16613_/B vssd1 vssd1 vccd1 vccd1 _16610_/Y sky130_fd_sc_hd__nor2_1
X_13822_ _13822_/A vssd1 vssd1 vccd1 vccd1 _13831_/S sky130_fd_sc_hd__buf_4
X_17590_ _17537_/X _17585_/X _17588_/Y _17589_/X vssd1 vssd1 vccd1 vccd1 _17590_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_141_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16541_ _16541_/A _16541_/B _16541_/C vssd1 vssd1 vccd1 vccd1 _19494_/D sky130_fd_sc_hd__nor3_1
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11276__B1 _11022_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13753_ _13753_/A vssd1 vssd1 vccd1 vccd1 _18443_/D sky130_fd_sc_hd__clkbuf_1
X_10965_ _10965_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10965_/Y sky130_fd_sc_hd__nand2_1
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12704_ _13009_/A vssd1 vssd1 vccd1 vccd1 _12704_/X sky130_fd_sc_hd__buf_2
XFILLER_16_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19260_ _19386_/CLK _19260_/D vssd1 vssd1 vccd1 vccd1 _19260_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__13017__A1 _15520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16472_ _16474_/A _16474_/C _16446_/X vssd1 vssd1 vccd1 vccd1 _16472_/Y sky130_fd_sc_hd__a21oi_1
X_13684_ _13330_/X _18413_/Q _13686_/S vssd1 vssd1 vccd1 vccd1 _13685_/A sky130_fd_sc_hd__mux2_1
X_10896_ _18488_/Q _18983_/Q _11071_/S vssd1 vssd1 vccd1 vccd1 _10897_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17951__A1 _19782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18211_ _18213_/A _18211_/B vssd1 vssd1 vccd1 vccd1 _18212_/A sky130_fd_sc_hd__and2_1
XANTENNA__11028__B1 _09481_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ _13054_/A vssd1 vssd1 vccd1 vccd1 _12635_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_184_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19306_/CLK sky130_fd_sc_hd__clkbuf_16
X_15423_ _15423_/A vssd1 vssd1 vccd1 vccd1 _19118_/D sky130_fd_sc_hd__clkbuf_1
X_19191_ _19502_/CLK _19191_/D vssd1 vssd1 vccd1 vccd1 _19191_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11579__A1 _19842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12776__B1 _11413_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18142_ _18142_/A _18142_/B vssd1 vssd1 vccd1 vccd1 _18142_/Y sky130_fd_sc_hd__nand2_1
X_15354_ _15354_/A vssd1 vssd1 vccd1 vccd1 _19087_/D sky130_fd_sc_hd__clkbuf_1
X_12566_ _12958_/A vssd1 vssd1 vccd1 vccd1 _12566_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_129_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09641__B1 _09640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10787__C1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14305_ _14305_/A vssd1 vssd1 vccd1 vccd1 _18647_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_8_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11517_ _17175_/A _17168_/A _17145_/A _11516_/X vssd1 vssd1 vccd1 vccd1 _11533_/B
+ sky130_fd_sc_hd__or4bb_1
X_15285_ _14576_/X _19057_/Q _15289_/S vssd1 vssd1 vccd1 vccd1 _15286_/A sky130_fd_sc_hd__mux2_1
X_18073_ _18073_/A vssd1 vssd1 vccd1 vccd1 _19804_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_117_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12497_ _12553_/C vssd1 vssd1 vccd1 vccd1 _17026_/S sky130_fd_sc_hd__buf_2
XFILLER_145_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16713__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17024_ _19662_/Q _17024_/B vssd1 vssd1 vccd1 vccd1 _17024_/X sky130_fd_sc_hd__or2_1
X_14236_ _18625_/Q _14001_/X _14242_/S vssd1 vssd1 vccd1 vccd1 _14237_/A sky130_fd_sc_hd__mux2_1
XANTENNA_output95_A _12432_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11448_ _11448_/A _11451_/A _11448_/C vssd1 vssd1 vccd1 vccd1 _11448_/Y sky130_fd_sc_hd__nand3_1
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_153_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11857__A _11879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ _18595_/Q _14007_/X _14169_/S vssd1 vssd1 vccd1 vccd1 _14168_/A sky130_fd_sc_hd__mux2_1
XFILLER_152_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11379_ _18416_/Q _18677_/Q _18576_/Q _18911_/Q _09743_/A _09733_/A vssd1 vssd1 vccd1
+ vccd1 _11380_/B sky130_fd_sc_hd__mux4_1
XFILLER_153_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_140_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _12975_/A _12975_/B _09305_/A input7/X _12976_/B vssd1 vssd1 vccd1 vccd1
+ _13254_/A sky130_fd_sc_hd__a41o_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_122_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19802_/CLK sky130_fd_sc_hd__clkbuf_16
X_14098_ _14109_/A vssd1 vssd1 vccd1 vccd1 _14107_/S sky130_fd_sc_hd__buf_2
X_18975_ _18975_/CLK _18975_/D vssd1 vssd1 vccd1 vccd1 _18975_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15763__S _15765_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _13048_/X _18295_/Q _13091_/S vssd1 vssd1 vccd1 vccd1 _13050_/A sky130_fd_sc_hd__mux2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _17937_/A vssd1 vssd1 vccd1 vccd1 _17935_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11503__A1 _11557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17857_ _17586_/X _17854_/Y _17856_/Y vssd1 vssd1 vccd1 vccd1 _17857_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15064__A _15080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16808_ _19576_/Q _16816_/D vssd1 vssd1 vccd1 vccd1 _16810_/B sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_137_clock clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 _19724_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17788_ _17790_/A _17790_/B vssd1 vssd1 vccd1 vccd1 _17788_/Y sky130_fd_sc_hd__nand2_1
XFILLER_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19527_ _19529_/CLK _19527_/D vssd1 vssd1 vccd1 vccd1 _19527_/Q sky130_fd_sc_hd__dfxtp_1
X_16739_ _16762_/A _16739_/B vssd1 vssd1 vccd1 vccd1 _16739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_81_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19458_ _19594_/CLK _19458_/D vssd1 vssd1 vccd1 vccd1 _19458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09211_ _09211_/A _09211_/B vssd1 vssd1 vccd1 vccd1 _09211_/Y sky130_fd_sc_hd__nand2_1
X_18409_ _19096_/CLK _18409_/D vssd1 vssd1 vccd1 vccd1 _18409_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10490__A1 _09764_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19389_ _19389_/CLK _19389_/D vssd1 vssd1 vccd1 vccd1 _19389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12767__B1 _11357_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09142_ _09142_/A _09167_/C _09175_/C vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__or3_1
XFILLER_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_163_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11767__A _19397_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _09975_/A _12474_/B vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__nor2_1
XFILLER_131_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13982__A _14049_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13193__S _13252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_93_clock_A clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13247__A1 _12712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12110__B _17768_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10750_ _10749_/B _12455_/B vssd1 vssd1 vccd1 vccd1 _10751_/B sky130_fd_sc_hd__and2b_1
XFILLER_53_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09700__A _09700_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ _11065_/A vssd1 vssd1 vccd1 vccd1 _09410_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_13_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15944__A0 _13538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10681_ _18460_/Q _19051_/Q _19213_/Q _18428_/Q _10566_/X _10586_/X vssd1 vssd1 vccd1
+ vccd1 _10682_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11105__S0 _09624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12758__B1 _11445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12420_ _12388_/A _12388_/B _12387_/A _12386_/A _12408_/A vssd1 vssd1 vccd1 vccd1
+ _12430_/B sky130_fd_sc_hd__a311o_1
XFILLER_166_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15848__S _15848_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _12351_/A _17878_/B vssd1 vssd1 vccd1 vccd1 _12351_/Y sky130_fd_sc_hd__nand2_1
XFILLER_154_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _11298_/X _11300_/X _11301_/X _10617_/A _09608_/A vssd1 vssd1 vccd1 vccd1
+ _11307_/B sky130_fd_sc_hd__o221a_1
XANTENNA__11981__A1 _11342_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15070_ _15070_/A vssd1 vssd1 vccd1 vccd1 _15070_/X sky130_fd_sc_hd__clkbuf_2
X_12282_ _12305_/A _17845_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12283_/B sky130_fd_sc_hd__a21boi_1
XFILLER_154_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14021_ _18535_/Q _14020_/X _14027_/S vssd1 vssd1 vccd1 vccd1 _14022_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13368__S _13387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _18450_/Q _19041_/Q _19203_/Q _18418_/Q _11074_/S _09511_/A vssd1 vssd1 vccd1
+ vccd1 _11233_/X sky130_fd_sc_hd__mux4_1
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_122_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11164_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15475__A2 _16024_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10115_ _10115_/A _10115_/B vssd1 vssd1 vccd1 vccd1 _10115_/Y sky130_fd_sc_hd__nand2_1
XFILLER_150_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18760_ _19247_/CLK _18760_/D vssd1 vssd1 vccd1 vccd1 _18760_/Q sky130_fd_sc_hd__dfxtp_1
X_15972_ _15983_/A vssd1 vssd1 vccd1 vccd1 _15981_/S sky130_fd_sc_hd__buf_4
X_11095_ _11016_/X _12448_/B _11070_/X _12447_/B vssd1 vssd1 vccd1 vccd1 _11465_/A
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_54_clock clkbuf_opt_1_0_clock/X vssd1 vssd1 vccd1 vccd1 _19379_/CLK sky130_fd_sc_hd__clkbuf_16
X_17711_ _17910_/A _17711_/B vssd1 vssd1 vccd1 vccd1 _17711_/Y sky130_fd_sc_hd__nand2_1
X_14923_ _14923_/A vssd1 vssd1 vccd1 vccd1 _18907_/D sky130_fd_sc_hd__clkbuf_1
X_10046_ _10046_/A _10046_/B vssd1 vssd1 vccd1 vccd1 _10046_/X sky130_fd_sc_hd__or2_1
X_18691_ _19373_/CLK _18691_/D vssd1 vssd1 vccd1 vccd1 _18691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_152_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10395__S1 _10436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17642_ _17642_/A _17642_/B vssd1 vssd1 vccd1 vccd1 _17642_/Y sky130_fd_sc_hd__nor2_1
X_14854_ _18877_/Q _14042_/X _14854_/S vssd1 vssd1 vccd1 vccd1 _14855_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13805_ _13138_/X _18466_/Q _13809_/S vssd1 vssd1 vccd1 vccd1 _13806_/A sky130_fd_sc_hd__mux2_1
X_17573_ _17398_/X _17572_/X _17573_/S vssd1 vssd1 vccd1 vccd1 _17574_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_69_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19223_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11997_ _11566_/A _12021_/A _12022_/A vssd1 vssd1 vccd1 vccd1 _11997_/Y sky130_fd_sc_hd__a21oi_1
X_14785_ _14620_/X _18847_/Q _14785_/S vssd1 vssd1 vccd1 vccd1 _14786_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10147__S1 _09871_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13831__S _13831_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19312_ _19312_/CLK _19312_/D vssd1 vssd1 vccd1 vccd1 _19312_/Q sky130_fd_sc_hd__dfxtp_1
X_16524_ _16524_/A _16529_/C vssd1 vssd1 vccd1 vccd1 _16524_/Y sky130_fd_sc_hd__nor2_1
XFILLER_44_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13736_ _13171_/X _18436_/Q _13736_/S vssd1 vssd1 vccd1 vccd1 _13737_/A sky130_fd_sc_hd__mux2_1
X_10948_ _10889_/A _10945_/X _10947_/X _10883_/X vssd1 vssd1 vccd1 vccd1 _10949_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16727__A2 _16750_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17924__A1 _12432_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15935__A0 _13525_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19243_ _19243_/CLK _19243_/D vssd1 vssd1 vccd1 vccd1 _19243_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16455_ _19468_/Q _16452_/B _16454_/Y vssd1 vssd1 vccd1 vccd1 _19468_/D sky130_fd_sc_hd__o21a_1
X_13667_ _13191_/X _18405_/Q _13675_/S vssd1 vssd1 vccd1 vccd1 _13668_/A sky130_fd_sc_hd__mux2_1
X_10879_ _18584_/Q _18855_/Q _19079_/Q _18823_/Q _11172_/S _10817_/X vssd1 vssd1 vccd1
+ vccd1 _10879_/X sky130_fd_sc_hd__mux4_1
XANTENNA__13132__A _13132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15406_ _15406_/A vssd1 vssd1 vccd1 vccd1 _19110_/D sky130_fd_sc_hd__clkbuf_1
X_12618_ _13422_/B vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__buf_2
X_19174_ _19237_/CLK _19174_/D vssd1 vssd1 vccd1 vccd1 _19174_/Q sky130_fd_sc_hd__dfxtp_1
X_16386_ _19444_/Q _16387_/C _19445_/Q vssd1 vssd1 vccd1 vccd1 _16388_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11016__A3 _11015_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ _13598_/A vssd1 vssd1 vccd1 vccd1 _18378_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__13410__B2 _18252_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10224__A1 _09909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18125_ _18125_/A _18135_/B vssd1 vssd1 vccd1 vccd1 _18125_/X sky130_fd_sc_hd__or2_1
XFILLER_145_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12549_ _12714_/A vssd1 vssd1 vccd1 vccd1 _12549_/X sky130_fd_sc_hd__buf_2
X_15337_ _19080_/Q _15025_/X _15339_/S vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__mux2_1
XANTENNA__11972__A1 _19340_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18056_ _18056_/A vssd1 vssd1 vccd1 vccd1 _19797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_145_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15268_ _15268_/A vssd1 vssd1 vccd1 vccd1 _19049_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_126_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17007_ _19656_/Q _17011_/B vssd1 vssd1 vccd1 vccd1 _17007_/X sky130_fd_sc_hd__or2_1
XANTENNA__09917__A1 _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14219_ _14219_/A vssd1 vssd1 vccd1 vccd1 _18617_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_160_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10491__A _19723_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15199_ _15199_/A vssd1 vssd1 vccd1 vccd1 _19018_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_99_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_98_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09760_ _09760_/A vssd1 vssd1 vccd1 vccd1 _09761_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_112_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_98_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18958_ _19098_/CLK _18958_/D vssd1 vssd1 vccd1 vccd1 _18958_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18089__B _18091_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_115_clock_A clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _17406_/X _17910_/B _17908_/X _17659_/X vssd1 vssd1 vccd1 vccd1 _17909_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11814__A1_N _11890_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ _18509_/Q _19004_/Q _11375_/S vssd1 vssd1 vccd1 vccd1 _09691_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18889_ _19081_/CLK _18889_/D vssd1 vssd1 vccd1 vccd1 _18889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14426__A0 _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_clock_A clkbuf_4_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14837__S _14843_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13741__S _13747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17915__A1 _12408_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14138__A _14195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _18745_/Q vssd1 vssd1 vccd1 vccd1 _13114_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_157_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_163_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_163_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_163_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_173_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17851__B1 _17850_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _18409_/Q _18670_/Q _18569_/Q _18904_/Q _10168_/S _09773_/A vssd1 vssd1 vccd1
+ vccd1 _09958_/X sky130_fd_sc_hd__mux4_1
XFILLER_44_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09889_ _18937_/Q _18703_/Q _19385_/Q _19033_/Q _10114_/S _09888_/X vssd1 vssd1 vccd1
+ vccd1 _09890_/B sky130_fd_sc_hd__mux4_1
XANTENNA__10377__S1 _10436_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11920_ _11919_/Y _19842_/Q _17183_/A vssd1 vssd1 vccd1 vccd1 _11920_/X sky130_fd_sc_hd__mux2_1
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_174_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ _11822_/X _11850_/Y _11821_/B vssd1 vssd1 vccd1 vccd1 _11851_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13651__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ _11174_/A vssd1 vssd1 vccd1 vccd1 _10802_/X sky130_fd_sc_hd__buf_2
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _14602_/A vssd1 vssd1 vccd1 vccd1 _14583_/S sky130_fd_sc_hd__clkbuf_8
X_11782_ _17563_/A _11782_/B vssd1 vssd1 vccd1 vccd1 _11842_/C sky130_fd_sc_hd__and2b_1
XFILLER_82_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13521_ _13521_/A vssd1 vssd1 vccd1 vccd1 _18354_/D sky130_fd_sc_hd__clkbuf_1
X_10733_ _18587_/Q _18858_/Q _19082_/Q _18826_/Q _11299_/S _09590_/A vssd1 vssd1 vccd1
+ vccd1 _10733_/X sky130_fd_sc_hd__mux4_1
XANTENNA__10576__A _10631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13452_ _13452_/A vssd1 vssd1 vccd1 vccd1 _18326_/D sky130_fd_sc_hd__clkbuf_1
X_16240_ _16240_/A vssd1 vssd1 vccd1 vccd1 _19391_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_174_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10664_ _18588_/Q _18859_/Q _19083_/Q _18827_/Q _10650_/X _09380_/A vssd1 vssd1 vccd1
+ vccd1 _10665_/B sky130_fd_sc_hd__mux4_1
XFILLER_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12403_ _17907_/B _12403_/B vssd1 vssd1 vccd1 vccd1 _12419_/A sky130_fd_sc_hd__xnor2_4
XFILLER_12_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16171_ _16239_/S vssd1 vssd1 vccd1 vccd1 _16180_/S sky130_fd_sc_hd__clkbuf_4
X_13383_ input25/X _13117_/X _13120_/X vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__a21o_1
XFILLER_139_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10595_ _09617_/X _10583_/X _10593_/X _09579_/A _10594_/Y vssd1 vssd1 vccd1 vccd1
+ _12461_/A sky130_fd_sc_hd__o32a_4
XFILLER_127_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15122_ _15122_/A vssd1 vssd1 vccd1 vccd1 _18984_/D sky130_fd_sc_hd__clkbuf_1
X_12334_ _12351_/A _12349_/A vssd1 vssd1 vccd1 vccd1 _12347_/B sky130_fd_sc_hd__xor2_4
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15053_ _15053_/A vssd1 vssd1 vccd1 vccd1 _18960_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_108_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12265_ _12265_/A _12289_/A vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__xnor2_4
XFILLER_142_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14004_ _14576_/A vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_123_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11216_ _11228_/A _11216_/B vssd1 vssd1 vccd1 vccd1 _11216_/Y sky130_fd_sc_hd__nor2_1
XFILLER_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_122_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19861_ _19866_/CLK _19861_/D vssd1 vssd1 vccd1 vccd1 _19861_/Q sky130_fd_sc_hd__dfxtp_1
X_12196_ _12196_/A _17810_/B vssd1 vssd1 vccd1 vccd1 _12197_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11557__D _11557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput71 _12488_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[0] sky130_fd_sc_hd__buf_2
XFILLER_123_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput82 _11612_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[1] sky130_fd_sc_hd__buf_2
X_18812_ _19388_/CLK _18812_/D vssd1 vssd1 vccd1 vccd1 _18812_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput93 _11644_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[2] sky130_fd_sc_hd__buf_2
X_11147_ _18915_/Q _18681_/Q _19363_/Q _19011_/Q _10962_/S _11075_/A vssd1 vssd1 vccd1
+ vccd1 _11147_/X sky130_fd_sc_hd__mux4_1
XFILLER_110_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16202__S _16202_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19792_ _19796_/CLK _19792_/D vssd1 vssd1 vccd1 vccd1 _19792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11854__B _11854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18743_ _19799_/CLK _18743_/D vssd1 vssd1 vccd1 vccd1 _18743_/Q sky130_fd_sc_hd__dfxtp_1
X_15955_ _13554_/X _19310_/Q _15959_/S vssd1 vssd1 vccd1 vccd1 _15956_/A sky130_fd_sc_hd__mux2_1
X_11078_ _11262_/A _11072_/Y _11075_/X _11077_/Y vssd1 vssd1 vccd1 vccd1 _11078_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_76_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14906_ _14917_/A vssd1 vssd1 vccd1 vccd1 _14915_/S sky130_fd_sc_hd__buf_2
XFILLER_64_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10029_ _10082_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _11426_/A sky130_fd_sc_hd__and2_1
XFILLER_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18674_ _19326_/CLK _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12682__A2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15886_ _15886_/A vssd1 vssd1 vccd1 vccd1 _19279_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17070__A1 _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17625_ _17457_/B _17612_/Y _17625_/S vssd1 vssd1 vccd1 vccd1 _17625_/X sky130_fd_sc_hd__mux2_1
X_14837_ _18869_/Q _14017_/X _14843_/S vssd1 vssd1 vccd1 vccd1 _14838_/A sky130_fd_sc_hd__mux2_1
XFILLER_17_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13561__S _13561_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11870__A _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17556_ _17550_/S _17437_/X _17399_/Y vssd1 vssd1 vccd1 vccd1 _17655_/B sky130_fd_sc_hd__a21o_1
X_14768_ _14595_/X _18839_/Q _14770_/S vssd1 vssd1 vccd1 vccd1 _14769_/A sky130_fd_sc_hd__mux2_1
X_16507_ _16321_/B _16504_/B _16506_/Y vssd1 vssd1 vccd1 vccd1 _19487_/D sky130_fd_sc_hd__o21a_1
XFILLER_108_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13719_ _13038_/X _18428_/Q _13725_/S vssd1 vssd1 vccd1 vccd1 _13720_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17487_ _17731_/S _17492_/B vssd1 vssd1 vccd1 vccd1 _17487_/Y sky130_fd_sc_hd__nand2_1
X_14699_ _14699_/A vssd1 vssd1 vccd1 vccd1 _18808_/D sky130_fd_sc_hd__clkbuf_1
X_19226_ _19471_/CLK _19226_/D vssd1 vssd1 vccd1 vccd1 _19226_/Q sky130_fd_sc_hd__dfxtp_1
X_16438_ _16440_/A _16440_/C _16402_/X vssd1 vssd1 vccd1 vccd1 _16438_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19157_ _19688_/CLK _19157_/D vssd1 vssd1 vccd1 vccd1 _19157_/Q sky130_fd_sc_hd__dfxtp_1
X_16369_ _19438_/Q _16371_/C _16368_/Y vssd1 vssd1 vccd1 vccd1 _19438_/D sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_41_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10748__A2 _10737_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18108_ _19818_/Q _18106_/X _18107_/X _18097_/X vssd1 vssd1 vccd1 vccd1 _19818_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088_ _19088_/CLK _19088_/D vssd1 vssd1 vccd1 vccd1 _19088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_172_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_173_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18039_ _18039_/A vssd1 vssd1 vccd1 vccd1 _19790_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11158__C1 _09553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09997__S0 _09850_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13736__S _13736_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _09812_/A vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__buf_4
XFILLER_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09515__A _10623_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ _09743_/A vssd1 vssd1 vccd1 vccd1 _11374_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_28_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15951__S _15959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13037__A _15035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ _09674_/A vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__buf_2
XFILLER_27_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17061__A1 _15542_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14567__S _14567_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16348__A _16890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11308__S0 _10729_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09921__S0 _09904_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11633__B1 _11632_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_167_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_161_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10987__A2 _12450_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15398__S _15400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11936__A1 _19339_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09108_ _09154_/A vssd1 vssd1 vccd1 vccd1 _09171_/B sky130_fd_sc_hd__clkbuf_2
XANTENNA__10295__S0 _10274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _10380_/A vssd1 vssd1 vccd1 vccd1 _10380_/Y sky130_fd_sc_hd__inv_2
XFILLER_124_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17907__A _17907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_163_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_105_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12050_ _12050_/A vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10047__S0 _09981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_132_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11001_ _11001_/A _11001_/B _11001_/C vssd1 vssd1 vccd1 vccd1 _11001_/X sky130_fd_sc_hd__or3_1
XFILLER_81_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_132_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09425__A _10823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15861__S _15865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ _15740_/A vssd1 vssd1 vccd1 vccd1 _19214_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__17642__A _17642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12952_ _13004_/A vssd1 vssd1 vccd1 vccd1 _12952_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10675__A1 _09989_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ _11903_/A _11903_/B vssd1 vssd1 vccd1 vccd1 _11904_/A sky130_fd_sc_hd__xnor2_4
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15671_ _14566_/X _19184_/Q _15671_/S vssd1 vssd1 vccd1 vccd1 _15672_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _12869_/X _12882_/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12883_/X sky130_fd_sc_hd__mux2_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17410_ _17534_/A _17410_/B vssd1 vssd1 vccd1 vccd1 _17410_/X sky130_fd_sc_hd__or2_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14622_/A vssd1 vssd1 vccd1 vccd1 _18778_/D sky130_fd_sc_hd__clkbuf_1
X_11834_ _19638_/Q _11832_/B _16086_/A vssd1 vssd1 vccd1 vccd1 _11834_/Y sky130_fd_sc_hd__o21ai_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _19305_/CLK _18390_/D vssd1 vssd1 vccd1 vccd1 _18390_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17341_ _17337_/Y _17340_/Y _17396_/A vssd1 vssd1 vccd1 vccd1 _17341_/X sky130_fd_sc_hd__mux2_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11624__B1 _19393_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11765_ _11765_/A vssd1 vssd1 vccd1 vccd1 _11765_/Y sky130_fd_sc_hd__clkinv_4
X_14553_ _14553_/A vssd1 vssd1 vccd1 vccd1 _14553_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _19276_/Q _19114_/Q _18523_/Q _18293_/Q _09645_/S _09541_/A vssd1 vssd1 vccd1
+ vccd1 _10717_/B sky130_fd_sc_hd__mux4_1
X_13504_ _13504_/A vssd1 vssd1 vccd1 vccd1 _18350_/D sky130_fd_sc_hd__clkbuf_1
X_17272_ _17367_/S vssd1 vssd1 vccd1 vccd1 _17291_/S sky130_fd_sc_hd__clkbuf_2
X_11696_ _11698_/B _11696_/B vssd1 vssd1 vccd1 vccd1 _11696_/Y sky130_fd_sc_hd__nand2_1
X_14484_ _14484_/A vssd1 vssd1 vccd1 vccd1 _18726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19011_ _19012_/CLK _19011_/D vssd1 vssd1 vccd1 vccd1 _19011_/Q sky130_fd_sc_hd__dfxtp_1
X_16223_ _16223_/A vssd1 vssd1 vccd1 vccd1 _19383_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_173_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13435_ _16619_/D _13435_/B vssd1 vssd1 vccd1 vccd1 _14197_/C sky130_fd_sc_hd__nand2_2
X_10647_ _10648_/A _12459_/A vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__nand2_1
XFILLER_158_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_173_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_155_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16154_ _16154_/A vssd1 vssd1 vccd1 vccd1 _19356_/D sky130_fd_sc_hd__clkbuf_1
X_13366_ _15095_/A vssd1 vssd1 vccd1 vccd1 _14617_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_10578_ _18399_/Q _18660_/Q _18559_/Q _18894_/Q _10576_/X _10577_/X vssd1 vssd1 vccd1
+ vccd1 _10578_/X sky130_fd_sc_hd__mux4_1
XFILLER_170_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15105_ _15105_/A vssd1 vssd1 vccd1 vccd1 _18976_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_154_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12317_ _12317_/A vssd1 vssd1 vccd1 vccd1 _12317_/Y sky130_fd_sc_hd__inv_4
XFILLER_127_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13297_ input20/X _13117_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _13297_/Y sky130_fd_sc_hd__a21oi_1
X_16085_ _16091_/A _16091_/C vssd1 vssd1 vccd1 vccd1 _16085_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_108_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_170_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15036_ _18955_/Q _15035_/X _15045_/S vssd1 vssd1 vccd1 vccd1 _15037_/A sky130_fd_sc_hd__mux2_1
X_12248_ _12248_/A _17835_/B vssd1 vssd1 vccd1 vccd1 _12249_/B sky130_fd_sc_hd__and2_1
XANTENNA__10589__S1 _10577_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19844_ _19846_/CLK _19844_/D vssd1 vssd1 vccd1 vccd1 _19844_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_111_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12179_ _12201_/B _12179_/B _12178_/X vssd1 vssd1 vccd1 vccd1 _12179_/X sky130_fd_sc_hd__or3b_1
XFILLER_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16094__A2 _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19775_ _19775_/CLK _19775_/D vssd1 vssd1 vccd1 vccd1 _19775_/Q sky130_fd_sc_hd__dfxtp_1
X_16987_ _19648_/Q _16998_/B vssd1 vssd1 vccd1 vccd1 _16987_/X sky130_fd_sc_hd__or2_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18726_ _19250_/CLK _18726_/D vssd1 vssd1 vccd1 vccd1 _18726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_97_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15938_ _15938_/A vssd1 vssd1 vccd1 vccd1 _19302_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__12655__A2 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10210__S0 _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18657_ _19310_/CLK _18657_/D vssd1 vssd1 vccd1 vccd1 _18657_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12696__A _12696_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15869_ _15869_/A vssd1 vssd1 vccd1 vccd1 _19271_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14387__S _14395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17608_ _17597_/X _17599_/Y _17607_/X _17333_/X vssd1 vssd1 vccd1 vccd1 _17608_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__10761__S1 _10655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09390_ _09390_/A _09390_/B vssd1 vssd1 vccd1 vccd1 _09390_/X sky130_fd_sc_hd__and2_1
XFILLER_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18588_ _18987_/CLK _18588_/D vssd1 vssd1 vccd1 vccd1 _18588_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17539_ _17252_/X _17732_/S vssd1 vssd1 vccd1 vccd1 _17539_/X sky130_fd_sc_hd__and2b_1
XANTENNA__10513__S1 _10310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19209_ _19241_/CLK _19209_/D vssd1 vssd1 vccd1 vccd1 _19209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_149_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_158_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_138_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14850__S _14854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13466__S _13470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15247__A _15315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input1_A io_dbus_rdata[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09726_ _09726_/A vssd1 vssd1 vccd1 vccd1 _09727_/A sky130_fd_sc_hd__buf_2
XANTENNA__10657__A1 _11313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09657_ _10680_/A _09654_/X _09656_/X vssd1 vssd1 vccd1 vccd1 _09657_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_83_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10752__S1 _11298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15596__A1 _19162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ _18511_/Q _19006_/Q _10542_/A vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__mux2_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11606__B1 _17230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16806__A _16806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10504__S1 _10310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _12179_/B vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_168_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10501_ _10414_/A _10500_/X _10236_/A vssd1 vssd1 vccd1 vccd1 _10501_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ _09664_/Y _11362_/X _11415_/X _11492_/D _11480_/X vssd1 vssd1 vccd1 vccd1
+ _11481_/X sky130_fd_sc_hd__a221o_2
XFILLER_137_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11909__A1 _11904_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13220_ _19446_/Q _13005_/X _13219_/X vssd1 vssd1 vccd1 vccd1 _13220_/X sky130_fd_sc_hd__o21a_1
XFILLER_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10432_ _10425_/Y _10427_/Y _10429_/Y _10431_/Y _09830_/A vssd1 vssd1 vccd1 vccd1
+ _10432_/X sky130_fd_sc_hd__o221a_4
X_13151_ _16091_/B _13152_/C _19758_/Q vssd1 vssd1 vccd1 vccd1 _13153_/B sky130_fd_sc_hd__a21oi_1
XFILLER_136_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ _10323_/A _10362_/X _10243_/X vssd1 vssd1 vccd1 vccd1 _10363_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_109_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12102_ _12654_/B vssd1 vssd1 vccd1 vccd1 _12102_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13082_ _19721_/Q _15540_/B _13143_/S vssd1 vssd1 vccd1 vccd1 _13082_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input57_A io_ibus_inst[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10294_ _10335_/A _10294_/B vssd1 vssd1 vccd1 vccd1 _10294_/Y sky130_fd_sc_hd__nor2_1
X_16910_ _16912_/B _16912_/C _16344_/A vssd1 vssd1 vccd1 vccd1 _16910_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_111_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12033_ _12008_/A _12008_/B _12005_/A vssd1 vssd1 vccd1 vccd1 _12034_/B sky130_fd_sc_hd__a21bo_1
XFILLER_2_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17890_ _17886_/B _17885_/B _17494_/X _17889_/Y vssd1 vssd1 vccd1 vccd1 _17890_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16841_ _19591_/Q _16838_/B _16840_/Y vssd1 vssd1 vccd1 vccd1 _19591_/D sky130_fd_sc_hd__o21a_1
XANTENNA__10440__S0 _10341_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19560_ _19564_/CLK _19560_/D vssd1 vssd1 vccd1 vccd1 _19560_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_9_clock_A clkbuf_4_1_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16772_ _19565_/Q _16778_/C _16772_/C _16772_/D vssd1 vssd1 vccd1 vccd1 _16782_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_65_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_93_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13984_ _13984_/A vssd1 vssd1 vccd1 vccd1 _18523_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18511_ _19006_/CLK _18511_/D vssd1 vssd1 vccd1 vccd1 _18511_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15723_ _15780_/S vssd1 vssd1 vccd1 vccd1 _15732_/S sky130_fd_sc_hd__buf_2
X_12935_ _19625_/Q _12605_/Y _12933_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _12935_/X
+ sky130_fd_sc_hd__a211o_1
X_19491_ _19491_/CLK _19491_/D vssd1 vssd1 vccd1 vccd1 _19491_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09271__A_N _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18442_ _19291_/CLK _18442_/D vssd1 vssd1 vccd1 vccd1 _18442_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15654_ _14541_/X _19176_/Q _15660_/S vssd1 vssd1 vccd1 vccd1 _15655_/A sky130_fd_sc_hd__mux2_1
XFILLER_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12865_/X _18286_/Q _12887_/S vssd1 vssd1 vccd1 vccd1 _12867_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14605_ _14605_/A vssd1 vssd1 vccd1 vccd1 _14605_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18373_ _19380_/CLK _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11817_ _17605_/A _11817_/B vssd1 vssd1 vccd1 vccd1 _11850_/A sky130_fd_sc_hd__xnor2_1
X_15585_ _15585_/A vssd1 vssd1 vccd1 vccd1 _19159_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16716__A _16762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _13119_/A vssd1 vssd1 vccd1 vccd1 _12976_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17309_/Y _17321_/X _17419_/A vssd1 vssd1 vccd1 vccd1 _17324_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12270__B1 _19416_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14536_ _14536_/A vssd1 vssd1 vccd1 vccd1 _18751_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11748_ _13419_/A _16951_/A vssd1 vssd1 vccd1 vccd1 _11749_/B sky130_fd_sc_hd__or2b_1
XFILLER_30_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17255_ _17249_/X _17435_/B _17446_/S vssd1 vssd1 vccd1 vccd1 _17255_/X sky130_fd_sc_hd__mux2_1
XFILLER_146_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14467_ _13870_/X _18719_/Q _14467_/S vssd1 vssd1 vccd1 vccd1 _14468_/A sky130_fd_sc_hd__mux2_1
X_11679_ _19774_/Q _11677_/X _11818_/S vssd1 vssd1 vccd1 vccd1 _17237_/A sky130_fd_sc_hd__mux2_8
XFILLER_146_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16206_ _16206_/A vssd1 vssd1 vccd1 vccd1 _19375_/D sky130_fd_sc_hd__clkbuf_1
X_13418_ _13418_/A _13418_/B vssd1 vssd1 vccd1 vccd1 _13419_/B sky130_fd_sc_hd__nand2_4
XFILLER_155_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17186_ _17190_/A _17432_/B vssd1 vssd1 vccd1 vccd1 _17404_/C sky130_fd_sc_hd__or2b_2
XFILLER_128_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14398_ _13873_/X _18688_/Q _14406_/S vssd1 vssd1 vccd1 vccd1 _14399_/A sky130_fd_sc_hd__mux2_1
XFILLER_155_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10179__A3 _10177_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16137_ _16137_/A vssd1 vssd1 vccd1 vccd1 _19353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14670__S _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13349_ _14614_/A vssd1 vssd1 vccd1 vccd1 _13349_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_170_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15511__A1 _19146_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16068_ _16068_/A vssd1 vssd1 vccd1 vccd1 _19341_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_97_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15067__A _15067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15019_ _15019_/A vssd1 vssd1 vccd1 vccd1 _15019_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_97_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12876__A2 _12784_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17264__A1 _17696_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_151_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19827_ _19828_/CLK _19827_/D vssd1 vssd1 vccd1 vccd1 _19827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10982__S1 _10910_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10004__A _10014_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ _19793_/CLK _19758_/D vssd1 vssd1 vccd1 vccd1 _19758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09511_ _09511_/A vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__buf_4
X_18709_ _18975_/CLK _18709_/D vssd1 vssd1 vccd1 vccd1 _18709_/Q sky130_fd_sc_hd__dfxtp_1
X_19689_ _19693_/CLK _19689_/D vssd1 vssd1 vccd1 vccd1 _19689_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15514__B hold18/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10939__A _11241_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10734__S1 _09705_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ _09442_/A vssd1 vssd1 vccd1 vccd1 _09443_/A sky130_fd_sc_hd__buf_2
XANTENNA__15578__A1 _19158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _11307_/A vssd1 vssd1 vccd1 vccd1 _09374_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_21_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_149_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_165_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_146_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15676__S _15682_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14580__S _14583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_133_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_133_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15502__A1 _16919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_133_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_163_clock_A clkbuf_4_9_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ _10310_/A vssd1 vssd1 vccd1 vccd1 _09710_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09703__A _10094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ _10981_/A _10981_/B vssd1 vssd1 vccd1 vccd1 _10981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12720_ _12720_/A vssd1 vssd1 vccd1 vccd1 _17937_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_128_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15569__A1 _15568_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_128_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12651_ _12557_/X _12649_/X _12650_/Y _12549_/X _18262_/Q vssd1 vssd1 vccd1 vccd1
+ _12651_/X sky130_fd_sc_hd__a32o_4
XANTENNA__09141__C _19863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14755__S _14759_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11602_ _11716_/D vssd1 vssd1 vccd1 vccd1 _17438_/S sky130_fd_sc_hd__clkbuf_2
X_12582_ _19570_/Q _12518_/X _12581_/X vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__a21o_1
X_15370_ _19095_/Q _15073_/X _15372_/S vssd1 vssd1 vccd1 vccd1 _15371_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14321_ _13870_/X _18655_/Q _14321_/S vssd1 vssd1 vccd1 vccd1 _14322_/A sky130_fd_sc_hd__mux2_1
X_11533_ _11562_/A _11533_/B _17110_/A _11533_/D vssd1 vssd1 vccd1 vccd1 _11533_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_128_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17040_ _17040_/A vssd1 vssd1 vccd1 vccd1 _19668_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14252_ _14252_/A vssd1 vssd1 vccd1 vccd1 _18632_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11464_ _11464_/A vssd1 vssd1 vccd1 vccd1 _11465_/C sky130_fd_sc_hd__clkinv_2
XFILLER_137_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13203_ _19609_/Q _12501_/X _12503_/X _19477_/Q _13202_/X vssd1 vssd1 vccd1 vccd1
+ _15580_/B sky130_fd_sc_hd__a221o_2
X_10415_ _18626_/Q _18961_/Q _10450_/S vssd1 vssd1 vccd1 vccd1 _10415_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_88_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11395_ _18608_/Q _18879_/Q _19103_/Q _18847_/Q _11388_/S _09788_/A vssd1 vssd1 vccd1
+ vccd1 _11395_/X sky130_fd_sc_hd__mux4_1
X_14183_ _18602_/Q _14029_/X _14191_/S vssd1 vssd1 vccd1 vccd1 _14184_/A sky130_fd_sc_hd__mux2_1
XFILLER_164_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16271__A _16890_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_99_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10346_ _18404_/Q _18665_/Q _18564_/Q _18899_/Q _10215_/S _10272_/A vssd1 vssd1 vccd1
+ vccd1 _10346_/X sky130_fd_sc_hd__mux4_1
X_13134_ _13166_/A vssd1 vssd1 vccd1 vccd1 _13134_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18991_ _19088_/CLK _18991_/D vssd1 vssd1 vccd1 vccd1 _18991_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10661__S0 _10660_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output163_A _12397_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _19746_/Q _19778_/Q _17946_/S vssd1 vssd1 vccd1 vccd1 _17943_/A sky130_fd_sc_hd__mux2_1
X_13065_ _13065_/A _13065_/B _13083_/B vssd1 vssd1 vccd1 vccd1 _13065_/X sky130_fd_sc_hd__or3_1
X_10277_ _10277_/A vssd1 vssd1 vccd1 vccd1 _10531_/A sky130_fd_sc_hd__clkbuf_2
X_12016_ _16978_/A _12044_/C vssd1 vssd1 vccd1 vccd1 _12016_/X sky130_fd_sc_hd__or2_1
XANTENNA__17246__A1 _12289_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_120_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17873_ _19733_/Q _17872_/X _17873_/S vssd1 vssd1 vccd1 vccd1 _17874_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13119__B _13254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16824_ _19581_/Q _16824_/B vssd1 vssd1 vccd1 vccd1 _16827_/B sky130_fd_sc_hd__and2_1
X_19612_ _19618_/CLK _19612_/D vssd1 vssd1 vccd1 vccd1 _19612_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_171_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19543_ _19543_/CLK _19543_/D vssd1 vssd1 vccd1 vccd1 _19543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16755_ _16760_/B _16760_/C _16718_/X vssd1 vssd1 vccd1 vccd1 _16755_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13967_ _18518_/Q _13965_/X _13979_/S vssd1 vssd1 vccd1 vccd1 _13968_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15706_ _14617_/X _19200_/Q _15708_/S vssd1 vssd1 vccd1 vccd1 _15707_/A sky130_fd_sc_hd__mux2_1
X_12918_ _19526_/Q _12939_/S _12699_/X _19494_/Q _12917_/X vssd1 vssd1 vccd1 vccd1
+ _12918_/X sky130_fd_sc_hd__a221o_1
X_19474_ _19610_/CLK _19474_/D vssd1 vssd1 vccd1 vccd1 _19474_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_94_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16757__B1 _19561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16686_ _16689_/C _16689_/D _19538_/Q vssd1 vssd1 vccd1 vccd1 _16688_/B sky130_fd_sc_hd__a21oi_1
X_13898_ _13898_/A vssd1 vssd1 vccd1 vccd1 _18498_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_94_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18425_ _19306_/CLK _18425_/D vssd1 vssd1 vccd1 vccd1 _18425_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15637_ _15637_/A vssd1 vssd1 vccd1 vccd1 _19169_/D sky130_fd_sc_hd__clkbuf_1
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ _12831_/X _12845_/X _12848_/Y input23/X _12781_/X vssd1 vssd1 vccd1 vccd1
+ _15006_/A sky130_fd_sc_hd__a32o_2
XANTENNA__16446__A _16546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12974__A _12974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__A1 _09477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18356_ _19237_/CLK _18356_/D vssd1 vssd1 vccd1 vccd1 _18356_/Q sky130_fd_sc_hd__dfxtp_1
X_15568_ _15565_/X _15566_/X _15567_/Y _15549_/X _18270_/Q vssd1 vssd1 vccd1 vccd1
+ _15568_/X sky130_fd_sc_hd__a32o_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17307_ _17391_/A _17457_/B vssd1 vssd1 vccd1 vccd1 _17483_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11141__S1 _10934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14519_ _14519_/A vssd1 vssd1 vccd1 vccd1 _14519_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_18287_ _19237_/CLK _18287_/D vssd1 vssd1 vccd1 vccd1 _18287_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10494__A _10494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15499_ _18258_/Q _15499_/B vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__or2_1
XFILLER_147_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17238_ _17492_/B _12358_/A _17274_/A vssd1 vssd1 vccd1 vccd1 _17238_/X sky130_fd_sc_hd__mux2_1
XFILLER_128_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13743__A0 _13228_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_156_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17169_ _17169_/A _17169_/B _17185_/A _17169_/D vssd1 vssd1 vccd1 vccd1 _17319_/B
+ sky130_fd_sc_hd__nor4_4
XFILLER_116_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_131_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10652__S0 _10650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15496__A0 _19713_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ _09726_/A _09979_/X _09984_/X _09990_/X _10040_/A vssd1 vssd1 vccd1 vccd1
+ _09991_/X sky130_fd_sc_hd__a311o_4
XFILLER_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10433__S _10433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12214__A _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_130_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10955__S1 _10934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15525__A _15636_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10669__A _10669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09425_ _10823_/A vssd1 vssd1 vccd1 vccd1 _11305_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09356_ _16937_/D vssd1 vssd1 vccd1 vccd1 _17133_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__11037__B2 _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_139_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_138_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10245__C1 _09670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09287_ _19822_/Q _19821_/Q _19819_/Q vssd1 vssd1 vccd1 vccd1 _09288_/C sky130_fd_sc_hd__or3_1
XFILLER_100_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_165_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17712__A2 _17709_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10891__S0 _10878_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_147_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10548__B1 _11313_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10200_/X sky130_fd_sc_hd__or2_1
XFILLER_107_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17476__A1 _19709_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11180_ _11195_/A _11180_/B vssd1 vssd1 vccd1 vccd1 _11180_/X sky130_fd_sc_hd__or2_1
XFILLER_161_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_122_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10131_ _11390_/A _10130_/X _09767_/A vssd1 vssd1 vccd1 vccd1 _10131_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_133_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_121_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10062_ _18412_/Q _18673_/Q _18572_/Q _18907_/Q _09538_/A _09542_/A vssd1 vssd1 vccd1
+ vccd1 _10062_/X sky130_fd_sc_hd__mux4_1
XFILLER_134_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15435__A _15446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__S1 _10934_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14870_ _14870_/A vssd1 vssd1 vccd1 vccd1 _18883_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_85_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13821_ _13821_/A vssd1 vssd1 vccd1 vccd1 _18473_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16540_ _19494_/Q _16540_/B _16540_/C vssd1 vssd1 vccd1 vccd1 _16541_/C sky130_fd_sc_hd__and3_1
XFILLER_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13752_ _13294_/X _18443_/Q _13758_/S vssd1 vssd1 vccd1 vccd1 _13753_/A sky130_fd_sc_hd__mux2_1
X_10964_ _18615_/Q _18950_/Q _10964_/S vssd1 vssd1 vccd1 vccd1 _10965_/B sky130_fd_sc_hd__mux2_1
XFILLER_44_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12703_ _13008_/A vssd1 vssd1 vccd1 vccd1 _12703_/X sky130_fd_sc_hd__clkbuf_2
X_16471_ _19474_/Q _16468_/B _16470_/Y vssd1 vssd1 vccd1 vccd1 _19474_/D sky130_fd_sc_hd__o21a_1
XANTENNA__14485__S _14489_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15411__A0 _19113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13683_ _13683_/A vssd1 vssd1 vccd1 vccd1 _18412_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10895_ _09367_/A _10885_/X _10894_/X _09470_/A _19714_/Q vssd1 vssd1 vccd1 vccd1
+ _10895_/X sky130_fd_sc_hd__a32o_2
X_18210_ _18210_/A vssd1 vssd1 vccd1 vccd1 _19852_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_31_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11028__A1 _11111_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15422_ _19118_/Q _15044_/X _15422_/S vssd1 vssd1 vccd1 vccd1 _15423_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19190_ _19319_/CLK _19190_/D vssd1 vssd1 vccd1 vccd1 _19190_/Q sky130_fd_sc_hd__dfxtp_1
X_12634_ _13261_/A vssd1 vssd1 vccd1 vccd1 _12634_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11579__A2 _11542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12776__A1 hold7/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18141_ _16619_/B _18134_/X _18140_/X _18136_/X vssd1 vssd1 vccd1 vccd1 _19831_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_129_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15353_ _19087_/Q _15047_/X _15361_/S vssd1 vssd1 vccd1 vccd1 _15354_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13402__B hold21/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12565_ _12565_/A vssd1 vssd1 vccd1 vccd1 _12565_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_141_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10518__S _10518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09641__A1 _11331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_145_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14304_ _13845_/X _18647_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _14305_/A sky130_fd_sc_hd__mux2_1
XFILLER_157_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18072_ _18150_/A _18072_/B vssd1 vssd1 vccd1 vccd1 _18073_/A sky130_fd_sc_hd__or2_1
X_11516_ _11516_/A vssd1 vssd1 vccd1 vccd1 _11516_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_156_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15284_ _15284_/A vssd1 vssd1 vccd1 vccd1 _19056_/D sky130_fd_sc_hd__clkbuf_1
X_12496_ _17133_/B _17028_/C _12496_/C vssd1 vssd1 vccd1 vccd1 _12553_/C sky130_fd_sc_hd__and3_1
XFILLER_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17023_ _17023_/A vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__inv_2
XFILLER_116_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13829__S _13831_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14235_ _14235_/A vssd1 vssd1 vccd1 vccd1 _18624_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_171_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11447_ _11451_/A _11448_/C _11448_/A vssd1 vssd1 vccd1 vccd1 _11447_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16205__S _16213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_125_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14166_ _14166_/A vssd1 vssd1 vccd1 vccd1 _18594_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_98_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11378_ _18608_/Q _18879_/Q _19103_/Q _18847_/Q _11375_/S _09715_/X vssd1 vssd1 vccd1
+ vccd1 _11378_/X sky130_fd_sc_hd__mux4_1
XANTENNA_output88_A _12291_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10329_ _09667_/A _10319_/X _10328_/X _09758_/A _19726_/Q vssd1 vssd1 vccd1 vccd1
+ _11351_/A sky130_fd_sc_hd__a32o_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ _13166_/A vssd1 vssd1 vccd1 vccd1 _13117_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _14097_/A vssd1 vssd1 vccd1 vccd1 _18564_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _18974_/CLK _18974_/D vssd1 vssd1 vccd1 vccd1 _18974_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13048_ _14560_/A vssd1 vssd1 vccd1 vccd1 _13048_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _19738_/Q _17430_/X _17924_/X vssd1 vssd1 vccd1 vccd1 _19738_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17856_ _17856_/A _17856_/B vssd1 vssd1 vccd1 vccd1 _17856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_78_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_1_0_clock_A clkbuf_3_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ _19575_/Q _19574_/Q _16807_/C vssd1 vssd1 vccd1 vccd1 _16816_/D sky130_fd_sc_hd__and3_1
XANTENNA__09343__A _19845_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17787_ _17790_/A _17790_/B _17832_/S vssd1 vssd1 vccd1 vccd1 _17787_/X sky130_fd_sc_hd__mux2_1
X_14999_ _15080_/A vssd1 vssd1 vccd1 vccd1 _15099_/S sky130_fd_sc_hd__buf_4
XFILLER_81_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11267__A1 _11033_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16738_ _16752_/D _16741_/C vssd1 vssd1 vccd1 vccd1 _16739_/B sky130_fd_sc_hd__and2_1
X_19526_ _19550_/CLK _19526_/D vssd1 vssd1 vccd1 vccd1 _19526_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19457_ _19529_/CLK _19457_/D vssd1 vssd1 vccd1 vccd1 _19457_/Q sky130_fd_sc_hd__dfxtp_1
X_16669_ _19532_/Q _19531_/Q _19530_/Q _16669_/D vssd1 vssd1 vccd1 vccd1 _16679_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_35_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14395__S _14395_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15080__A _15080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ _11513_/C vssd1 vssd1 vccd1 vccd1 _09210_/X sky130_fd_sc_hd__buf_2
X_18408_ _19127_/CLK _18408_/D vssd1 vssd1 vccd1 vccd1 _18408_/Q sky130_fd_sc_hd__dfxtp_1
X_19388_ _19388_/CLK _19388_/D vssd1 vssd1 vccd1 vccd1 _19388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09141_ _19865_/Q _19864_/Q _19863_/Q vssd1 vssd1 vccd1 vccd1 _09175_/C sky130_fd_sc_hd__or3_1
X_18339_ _19058_/CLK _18339_/D vssd1 vssd1 vccd1 vccd1 _18339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_111_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13739__S _13747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_116_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09518__A _11318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_116_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_144_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_103_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16130__A1 _19352_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09237__B _11569_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _10087_/A _12473_/B vssd1 vssd1 vccd1 vccd1 _10088_/A sky130_fd_sc_hd__nand2_1
XFILLER_131_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_130_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_130_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12598__B _16245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_clock_A clkbuf_4_4_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19586__CLK _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16086__A _16086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09408_ _18779_/Q vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_71_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10680_ _10680_/A _10680_/B vssd1 vssd1 vccd1 vccd1 _10680_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11105__S1 _11020_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_166_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09339_ _18122_/A _17126_/B _11584_/B _17126_/C vssd1 vssd1 vccd1 vccd1 _09339_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _12351_/A _17878_/B _12335_/X vssd1 vssd1 vccd1 vccd1 _12350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_166_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_138_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13649__S _13653_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11301_ _18925_/Q _18691_/Q _19373_/Q _19021_/Q _10542_/A _09443_/A vssd1 vssd1 vccd1
+ vccd1 _11301_/X sky130_fd_sc_hd__mux4_1
XFILLER_138_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12281_ _12301_/A _12474_/B _12280_/Y vssd1 vssd1 vccd1 vccd1 _17856_/A sky130_fd_sc_hd__o21ai_4
XFILLER_119_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10862__A _11071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14020_ _14592_/A vssd1 vssd1 vccd1 vccd1 _14020_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_11232_ _11232_/A _11232_/B vssd1 vssd1 vccd1 vccd1 _11232_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14380__A0 _13848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10616__S0 _10670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09428__A _10042_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_150_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ _18452_/Q _19043_/Q _19205_/Q _18420_/Q _10904_/X _11072_/A vssd1 vssd1 vccd1
+ vccd1 _11164_/B sky130_fd_sc_hd__mux4_2
XFILLER_84_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_121_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_96_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10941__B1 _10807_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _18632_/Q _18967_/Q _10114_/S vssd1 vssd1 vccd1 vccd1 _10115_/B sky130_fd_sc_hd__mux2_1
XFILLER_122_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15971_ _15971_/A vssd1 vssd1 vccd1 vccd1 _19317_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11094_ _09477_/A _11083_/X _11092_/X _09577_/A _11093_/Y vssd1 vssd1 vccd1 vccd1
+ _12447_/B sky130_fd_sc_hd__o32a_4
XFILLER_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17710_ _17708_/X _17711_/B _17710_/S vssd1 vssd1 vccd1 vccd1 _17710_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14922_ _18907_/Q _14036_/X _14926_/S vssd1 vssd1 vccd1 vccd1 _14923_/A sky130_fd_sc_hd__mux2_1
X_10045_ _18476_/Q _19067_/Q _19229_/Q _18444_/Q _09441_/X _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10046_/B sky130_fd_sc_hd__mux4_1
XFILLER_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18690_ _19086_/CLK _18690_/D vssd1 vssd1 vccd1 vccd1 _18690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_102_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17641_ _17639_/X _17640_/Y _17710_/S vssd1 vssd1 vccd1 vccd1 _17641_/X sky130_fd_sc_hd__mux2_1
XANTENNA__17621__A1 _19714_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14853_ _14853_/A vssd1 vssd1 vccd1 vccd1 _18876_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15632__A0 _19737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13804_ _13804_/A vssd1 vssd1 vccd1 vccd1 _18465_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__11249__A1 _11254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17572_ _17436_/Y _17441_/Y _17572_/S vssd1 vssd1 vccd1 vccd1 _17572_/X sky130_fd_sc_hd__mux2_1
X_14784_ _14784_/A vssd1 vssd1 vccd1 vccd1 _18846_/D sky130_fd_sc_hd__clkbuf_1
X_11996_ _12011_/A _11665_/X _11992_/X _11995_/Y vssd1 vssd1 vccd1 vccd1 _16272_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_16_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19311_ _19311_/CLK _19311_/D vssd1 vssd1 vccd1 vccd1 _19311_/Q sky130_fd_sc_hd__dfxtp_1
X_16523_ _16533_/D vssd1 vssd1 vccd1 vccd1 _16529_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13735_ _13735_/A vssd1 vssd1 vccd1 vccd1 _18435_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10947_ _11048_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _10947_/X sky130_fd_sc_hd__or2_1
XFILLER_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19242_ _19243_/CLK _19242_/D vssd1 vssd1 vccd1 vccd1 _19242_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15104__S _15112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16454_ _16470_/A _16458_/C vssd1 vssd1 vccd1 vccd1 _16454_/Y sky130_fd_sc_hd__nor2_1
X_13666_ _13677_/A vssd1 vssd1 vccd1 vccd1 _13675_/S sky130_fd_sc_hd__clkbuf_4
X_10878_ _10878_/A vssd1 vssd1 vccd1 vccd1 _11172_/S sky130_fd_sc_hd__buf_4
XANTENNA__12749__A1 _18262_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15405_ _19110_/Q _15019_/X _15411_/S vssd1 vssd1 vccd1 vccd1 _15406_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13132__B _13132_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12617_ _18254_/Q _12614_/Y _12616_/X vssd1 vssd1 vccd1 vccd1 _13422_/B sky130_fd_sc_hd__o21a_2
X_19173_ _19237_/CLK _19173_/D vssd1 vssd1 vccd1 vccd1 _19173_/Q sky130_fd_sc_hd__dfxtp_1
X_16385_ _19444_/Q _16387_/C _16384_/Y vssd1 vssd1 vccd1 vccd1 _19444_/D sky130_fd_sc_hd__o21a_1
XANTENNA__17137__B1 _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ _18378_/Q _13595_/X _13609_/S vssd1 vssd1 vccd1 vccd1 _13598_/A sky130_fd_sc_hd__mux2_1
XANTENNA__16724__A _19551_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18124_ _13391_/A _18120_/X _18122_/X _18123_/X vssd1 vssd1 vccd1 vccd1 _19824_/D
+ sky130_fd_sc_hd__o211a_1
X_15336_ _15336_/A vssd1 vssd1 vccd1 vccd1 _19079_/D sky130_fd_sc_hd__clkbuf_1
X_12548_ _12548_/A vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__17688__B2 _11932_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_129_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18055_ _19797_/Q _12321_/A _18061_/S vssd1 vssd1 vccd1 vccd1 _18056_/A sky130_fd_sc_hd__mux2_1
X_15267_ _14550_/X _19049_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15268_/A sky130_fd_sc_hd__mux2_1
X_12479_ _12480_/A _12479_/B vssd1 vssd1 vccd1 vccd1 _12479_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_160_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17006_ _12715_/X _16997_/X _17005_/X _16995_/X vssd1 vssd1 vccd1 vccd1 _19655_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09338__A _18130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10607__S0 _10670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14218_ _18617_/Q _13975_/X _14220_/S vssd1 vssd1 vccd1 vccd1 _14219_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_172_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_126_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15198_ _19018_/Q _15031_/X _15206_/S vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__mux2_1
XANTENNA__18101__A2 _18086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15774__S _15776_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16112__A1 _19349_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_113_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14149_ _14195_/S vssd1 vssd1 vccd1 vccd1 _14158_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_141_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_141_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18957_ _19006_/CLK _18957_/D vssd1 vssd1 vccd1 vccd1 _18957_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_140_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _11512_/B _17906_/B _17462_/X _17907_/X vssd1 vssd1 vccd1 vccd1 _17908_/X
+ sky130_fd_sc_hd__o211a_1
X_09690_ _09690_/A vssd1 vssd1 vccd1 vccd1 _10138_/A sky130_fd_sc_hd__buf_2
XFILLER_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18888_ _19081_/CLK _18888_/D vssd1 vssd1 vccd1 vccd1 _18888_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17839_ _17571_/X _17625_/X _17838_/X _17592_/X vssd1 vssd1 vccd1 vccd1 _17839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_82_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__A1 _19561_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19509_ _19540_/CLK _19509_/D vssd1 vssd1 vccd1 vccd1 _19509_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_5_0_clock_A clkbuf_4_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10947__A _11048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_109_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09124_ _09124_/A _09124_/B vssd1 vssd1 vccd1 vccd1 _17166_/A sky130_fd_sc_hd__nand2_8
XFILLER_109_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_148_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10682__A _10682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_144_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11715__A2 _12445_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_132_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _09905_/X _09953_/Y _09956_/Y _10205_/A vssd1 vssd1 vccd1 vccd1 _09957_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_131_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_183_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19241_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_131_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09888_ _09954_/A vssd1 vssd1 vccd1 vccd1 _09888_/X sky130_fd_sc_hd__clkbuf_4
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15614__A0 _13306_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13932__S _13935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11850_ _11850_/A _17245_/A vssd1 vssd1 vccd1 vccd1 _11850_/Y sky130_fd_sc_hd__nand2_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__12979__A1 _11538_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09711__A _10238_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _10801_/A vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__buf_4
XFILLER_82_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _11670_/A _12449_/B _11813_/A _18135_/A vssd1 vssd1 vccd1 vccd1 _17587_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13520_ _18354_/Q _13519_/X _13529_/S vssd1 vssd1 vccd1 vccd1 _13521_/A sky130_fd_sc_hd__mux2_1
XFILLER_159_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10732_ _10031_/A _10729_/X _10731_/X vssd1 vssd1 vccd1 vccd1 _10732_/X sky130_fd_sc_hd__a21o_1
XFILLER_158_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_121_clock clkbuf_4_14_0_clock/X vssd1 vssd1 vccd1 vccd1 _19854_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__15859__S _15865_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13451_ _12907_/X _18326_/Q _13459_/S vssd1 vssd1 vccd1 vccd1 _13452_/A sky130_fd_sc_hd__mux2_1
X_10663_ _10653_/X _10657_/X _10659_/X _10662_/X _09614_/X vssd1 vssd1 vccd1 vccd1
+ _10663_/X sky130_fd_sc_hd__a221o_4
XANTENNA__17119__B1 _17907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12402_ _17387_/B _12401_/Y _12381_/B vssd1 vssd1 vccd1 vccd1 _12403_/B sky130_fd_sc_hd__o21a_1
X_16170_ _16226_/A vssd1 vssd1 vccd1 vccd1 _16239_/S sky130_fd_sc_hd__buf_4
XFILLER_127_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10594_ _19721_/Q vssd1 vssd1 vccd1 vccd1 _10594_/Y sky130_fd_sc_hd__inv_2
X_13382_ _13370_/Y _13371_/X _13381_/X _12848_/A vssd1 vssd1 vccd1 vccd1 _13382_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_154_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17134__A3 _17149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15121_ _18984_/Q _15025_/X _15123_/S vssd1 vssd1 vccd1 vccd1 _15122_/A sky130_fd_sc_hd__mux2_1
X_12333_ _19798_/Q _10080_/A _12404_/S vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__mux2_8
XFILLER_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_136_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19780_/CLK sky130_fd_sc_hd__clkbuf_16
X_15052_ _18960_/Q _15051_/X _15061_/S vssd1 vssd1 vccd1 vccd1 _15053_/A sky130_fd_sc_hd__mux2_1
XFILLER_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12264_ _19795_/Q _10087_/A _12357_/S vssd1 vssd1 vccd1 vccd1 _12289_/A sky130_fd_sc_hd__mux2_8
XFILLER_107_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_108_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14999__A _15080_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14003_ _14003_/A vssd1 vssd1 vccd1 vccd1 _18529_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18095__A1 _14860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ _18913_/Q _18679_/Q _19361_/Q _19009_/Q _10969_/A _09511_/A vssd1 vssd1 vccd1
+ vccd1 _11216_/B sky130_fd_sc_hd__mux4_1
X_19860_ _19866_/CLK _19860_/D vssd1 vssd1 vccd1 vccd1 _19860_/Q sky130_fd_sc_hd__dfxtp_1
X_12195_ _12195_/A vssd1 vssd1 vccd1 vccd1 _17810_/B sky130_fd_sc_hd__buf_2
XANTENNA__14105__A0 _13915_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput72 _11904_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[10] sky130_fd_sc_hd__buf_2
X_18811_ _19197_/CLK _18811_/D vssd1 vssd1 vccd1 vccd1 _18811_/Q sky130_fd_sc_hd__dfxtp_1
X_11146_ _09366_/A _11136_/X _11145_/X _09469_/A _19709_/Q vssd1 vssd1 vccd1 vccd1
+ _11284_/A sky130_fd_sc_hd__a32o_4
Xoutput83 _12175_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[20] sky130_fd_sc_hd__buf_2
XFILLER_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput94 _12408_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[30] sky130_fd_sc_hd__buf_2
XFILLER_96_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19791_ _19802_/CLK _19791_/D vssd1 vssd1 vccd1 vccd1 _19791_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_49_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_95_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13408__A _18252_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15954_ _15954_/A vssd1 vssd1 vccd1 vccd1 _19309_/D sky130_fd_sc_hd__clkbuf_1
X_11077_ _11232_/A _11077_/B vssd1 vssd1 vccd1 vccd1 _11077_/Y sky130_fd_sc_hd__nor2_1
X_18742_ _19706_/CLK _18742_/D vssd1 vssd1 vccd1 vccd1 _18742_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_163_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14905_ _14905_/A vssd1 vssd1 vccd1 vccd1 _18899_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10028_ _09760_/A _10012_/X _10026_/X _09833_/A _10027_/Y vssd1 vssd1 vccd1 vccd1
+ _12476_/B sky130_fd_sc_hd__o32a_4
XFILLER_49_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18673_ _19006_/CLK _18673_/D vssd1 vssd1 vccd1 vccd1 _18673_/Q sky130_fd_sc_hd__dfxtp_1
X_15885_ _19279_/Q _14563_/A _15887_/S vssd1 vssd1 vccd1 vccd1 _15886_/A sky130_fd_sc_hd__mux2_1
XFILLER_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12031__B _17211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14836_ _14836_/A vssd1 vssd1 vccd1 vccd1 _18868_/D sky130_fd_sc_hd__clkbuf_1
X_17624_ _17622_/Y _17623_/X _17739_/S vssd1 vssd1 vccd1 vccd1 _17624_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_91_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15620__A3 _09234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17555_ _17657_/A _17554_/X _17732_/S vssd1 vssd1 vccd1 vccd1 _17555_/X sky130_fd_sc_hd__mux2_2
XFILLER_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_91_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _14767_/A vssd1 vssd1 vccd1 vccd1 _18838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11979_ _12025_/A _12025_/B _12111_/A vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__o21ai_1
XFILLER_17_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16506_ _16321_/B _16504_/B _16489_/X vssd1 vssd1 vccd1 vccd1 _16506_/Y sky130_fd_sc_hd__a21oi_1
X_13718_ _13718_/A vssd1 vssd1 vccd1 vccd1 _18427_/D sky130_fd_sc_hd__clkbuf_1
X_17486_ _17504_/S _17492_/B _17896_/S vssd1 vssd1 vccd1 vccd1 _17486_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14698_ _14598_/X _18808_/Q _14698_/S vssd1 vssd1 vccd1 vccd1 _14699_/A sky130_fd_sc_hd__mux2_1
XANTENNA__13919__A0 _13918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16437_ _19462_/Q _16433_/B _16436_/Y vssd1 vssd1 vccd1 vccd1 _19462_/D sky130_fd_sc_hd__o21a_1
X_19225_ _19382_/CLK _19225_/D vssd1 vssd1 vccd1 vccd1 _19225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_108_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13649_ _13048_/X _18397_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13650_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_164_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19156_ _19694_/CLK _19156_/D vssd1 vssd1 vccd1 vccd1 _19156_/Q sky130_fd_sc_hd__dfxtp_1
X_16368_ _19438_/Q _16371_/C _16359_/X vssd1 vssd1 vccd1 vccd1 _16368_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_9_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10828__S0 _09598_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18107_ _18107_/A _18116_/B vssd1 vssd1 vccd1 vccd1 _18107_/X sky130_fd_sc_hd__or2_1
XFILLER_9_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15319_ _15387_/S vssd1 vssd1 vccd1 vccd1 _15328_/S sky130_fd_sc_hd__buf_4
XANTENNA__10748__A3 _10747_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19087_ _19119_/CLK _19087_/D vssd1 vssd1 vccd1 vccd1 _19087_/Q sky130_fd_sc_hd__dfxtp_1
X_16299_ _16299_/A vssd1 vssd1 vccd1 vccd1 _19417_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_133_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18038_ _19790_/Q _19411_/Q _18038_/S vssd1 vssd1 vccd1 vccd1 _18039_/A sky130_fd_sc_hd__mux2_1
XFILLER_132_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11253__S0 _09410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ _09811_/A vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__buf_4
XFILLER_140_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09742_ _09859_/A _09742_/B _09742_/C vssd1 vssd1 vccd1 vccd1 _09742_/X sky130_fd_sc_hd__or3_1
XFILLER_101_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09749__S1 _09715_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09673_ _10229_/A vssd1 vssd1 vccd1 vccd1 _09674_/A sky130_fd_sc_hd__buf_2
XFILLER_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14848__S _14854_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13752__S _13758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11881__A1 _11877_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__S1 _10655_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14149__A _14195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18010__A1 _11826_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09921__S1 _09888_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13988__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_168_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__14583__S _14583_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12189__A2 _12470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_53_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19378_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09107_ _09328_/A _09325_/A vssd1 vssd1 vccd1 vccd1 _09154_/A sky130_fd_sc_hd__nor2_1
XANTENNA__10295__S1 _10263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_108_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_123_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17907__B _17907_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12116__B _17219_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_68_clock clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 _19384_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17195__A _17195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10047__S1 _09708_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11000_ _10807_/A _10996_/X _10999_/X _09447_/A vssd1 vssd1 vccd1 vccd1 _11001_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17824__A1 _17820_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _13261_/A vssd1 vssd1 vccd1 vccd1 _12951_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13662__S _13664_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11854_/A _11854_/B _11876_/A _11901_/X vssd1 vssd1 vccd1 vccd1 _11903_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_93_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15670_ _15670_/A vssd1 vssd1 vccd1 vccd1 _19183_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _19711_/Q _15479_/B _13103_/S vssd1 vssd1 vccd1 vccd1 _12882_/X sky130_fd_sc_hd__mux2_1
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09441__A _10670_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14621_ _14620_/X _18778_/Q _14621_/S vssd1 vssd1 vccd1 vccd1 _14622_/A sky130_fd_sc_hd__mux2_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _15474_/A vssd1 vssd1 vccd1 vccd1 _16086_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17340_ _17340_/A vssd1 vssd1 vccd1 vccd1 _17340_/Y sky130_fd_sc_hd__inv_2
XANTENNA__18001__A1 _19394_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14552_/A vssd1 vssd1 vccd1 vccd1 _18756_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _11788_/C _11764_/B vssd1 vssd1 vccd1 vccd1 _11765_/A sky130_fd_sc_hd__xnor2_4
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_159_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13349_/X _18350_/Q _13503_/S vssd1 vssd1 vccd1 vccd1 _13504_/A sky130_fd_sc_hd__mux2_1
X_17271_ _17819_/B _17642_/B _17286_/S vssd1 vssd1 vccd1 vccd1 _17365_/B sky130_fd_sc_hd__mux2_1
X_10715_ _09630_/A _10712_/Y _10714_/Y _09658_/A vssd1 vssd1 vccd1 vccd1 _10715_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__10832__C1 _11307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14483_ _13893_/X _18726_/Q _14489_/S vssd1 vssd1 vccd1 vccd1 _14484_/A sky130_fd_sc_hd__mux2_1
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11695_ _11803_/A _19584_/Q _11805_/C vssd1 vssd1 vccd1 vccd1 _11695_/Y sky130_fd_sc_hd__o21ai_1
X_19010_ _19736_/CLK _19010_/D vssd1 vssd1 vccd1 vccd1 _19010_/Q sky130_fd_sc_hd__dfxtp_1
X_16222_ _13589_/X _19383_/Q _16224_/S vssd1 vssd1 vccd1 vccd1 _16223_/A sky130_fd_sc_hd__mux2_1
XFILLER_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13434_ _14197_/B vssd1 vssd1 vccd1 vccd1 _14371_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_174_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10646_ _09617_/X _10630_/X _10644_/X _09579_/A _10645_/Y vssd1 vssd1 vccd1 vccd1
+ _12459_/A sky130_fd_sc_hd__o32a_4
XANTENNA_clkbuf_leaf_5_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16153_ _16152_/X _19356_/Q _16167_/S vssd1 vssd1 vccd1 vccd1 _16154_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_158_clock_A clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13365_ _13365_/A _13365_/B vssd1 vssd1 vccd1 vccd1 _15095_/A sky130_fd_sc_hd__nor2_4
XFILLER_6_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10577_ _10586_/A vssd1 vssd1 vccd1 vccd1 _10577_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15104_ _18976_/Q _14996_/X _15112_/S vssd1 vssd1 vccd1 vccd1 _15105_/A sky130_fd_sc_hd__mux2_1
XFILLER_170_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12316_ _12347_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12317_/A sky130_fd_sc_hd__xnor2_1
X_16084_ _16084_/A vssd1 vssd1 vccd1 vccd1 _19344_/D sky130_fd_sc_hd__clkbuf_1
X_13296_ _13296_/A vssd1 vssd1 vccd1 vccd1 _18309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_154_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15035_ _15035_/A vssd1 vssd1 vccd1 vccd1 _15035_/X sky130_fd_sc_hd__clkbuf_2
X_12247_ _12267_/A vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__inv_2
XANTENNA__16213__S _16213_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14522__A _14621_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19843_ _19846_/CLK _19843_/D vssd1 vssd1 vccd1 vccd1 _19843_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_122_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10363__A1 _10323_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_110_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ _19412_/Q _12226_/C vssd1 vssd1 vccd1 vccd1 _12178_/X sky130_fd_sc_hd__or2_1
XFILLER_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_111_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_95_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11129_ _09393_/A _11128_/X _11208_/A vssd1 vssd1 vccd1 vccd1 _11129_/X sky130_fd_sc_hd__a21o_1
X_19774_ _19786_/CLK _19774_/D vssd1 vssd1 vccd1 vccd1 _19774_/Q sky130_fd_sc_hd__dfxtp_1
X_16986_ _17013_/A vssd1 vssd1 vccd1 vccd1 _16998_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_77_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13301__B2 _19355_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18725_ _19249_/CLK _18725_/D vssd1 vssd1 vccd1 vccd1 _18725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15937_ _13528_/X _19302_/Q _15937_/S vssd1 vssd1 vccd1 vccd1 _15938_/A sky130_fd_sc_hd__mux2_1
XFILLER_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14668__S _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16449__A _16549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17044__S _17050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10210__S1 _09954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15868_ _19271_/Q _14537_/A _15876_/S vssd1 vssd1 vccd1 vccd1 _15869_/A sky130_fd_sc_hd__mux2_1
X_18656_ _19370_/CLK _18656_/D vssd1 vssd1 vccd1 vccd1 _18656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12696__B input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09351__A _09351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17607_ _17413_/X _17602_/X _17606_/Y _17532_/X vssd1 vssd1 vccd1 vccd1 _17607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_36_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14819_ _18861_/Q _13991_/X _14821_/S vssd1 vssd1 vccd1 vccd1 _14820_/A sky130_fd_sc_hd__mux2_1
X_15799_ _15799_/A vssd1 vssd1 vccd1 vccd1 _19240_/D sky130_fd_sc_hd__clkbuf_1
X_18587_ _18974_/CLK _18587_/D vssd1 vssd1 vccd1 vccd1 _18587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17538_ _17406_/X _17533_/X _17536_/X _17537_/X vssd1 vssd1 vccd1 vccd1 _17538_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_33_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17469_ _17461_/A _17463_/B _17419_/X _17467_/X _17468_/Y vssd1 vssd1 vccd1 vccd1
+ _17469_/X sky130_fd_sc_hd__o2111a_1
XANTENNA__17751__B1 _17750_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_149_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19208_ _19306_/CLK _19208_/D vssd1 vssd1 vccd1 vccd1 _19208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19139_ _19668_/CLK _19139_/D vssd1 vssd1 vccd1 vccd1 _19139_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16306__A1 _12391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14317__A0 _13864_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_145_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_160_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13747__S _13747_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18059__A1 _19420_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_154_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__17806__A1 _17733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_114_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15962__S _15970_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13048__A _14560_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09725_ _11380_/A vssd1 vssd1 vccd1 vccd1 _11373_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16359__A _16546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_103_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09656_ _09632_/A _09655_/X _10073_/A vssd1 vssd1 vccd1 vccd1 _09656_/X sky130_fd_sc_hd__o21a_1
XFILLER_83_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _10660_/A vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__buf_4
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10200__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_168_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16545__A1 _19495_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10500_ _18496_/Q _18991_/Q _10500_/S vssd1 vssd1 vccd1 vccd1 _10500_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13511__A _16619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15202__S _15206_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_168_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_149_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ _11417_/A _11415_/A _11428_/X _11478_/X _11479_/Y vssd1 vssd1 vccd1 vccd1
+ _11480_/X sky130_fd_sc_hd__a2111o_1
XFILLER_149_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10431_ _10394_/A _10430_/X _09764_/A vssd1 vssd1 vccd1 vccd1 _10431_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16822__A _16838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14308__A0 _13851_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13150_ _13150_/A vssd1 vssd1 vccd1 vccd1 _18301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_163_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10362_ _18467_/Q _19058_/Q _19220_/Q _18435_/Q _10247_/X _10238_/X vssd1 vssd1 vccd1
+ vccd1 _10362_/X sky130_fd_sc_hd__mux4_2
XFILLER_163_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12101_ _12099_/Y _12092_/Y _12341_/S vssd1 vssd1 vccd1 vccd1 _12101_/X sky130_fd_sc_hd__mux2_1
X_10293_ _18469_/Q _19060_/Q _19222_/Q _18437_/Q _10286_/X _10275_/X vssd1 vssd1 vccd1
+ vccd1 _10294_/B sky130_fd_sc_hd__mux4_1
X_13081_ _19602_/Q _12633_/X _12634_/X _19470_/Q _13080_/X vssd1 vssd1 vccd1 vccd1
+ _15540_/B sky130_fd_sc_hd__a221o_2
XFILLER_105_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09436__A _09596_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ _12032_/A _12032_/B vssd1 vssd1 vccd1 vccd1 _12034_/A sky130_fd_sc_hd__nor2_1
XFILLER_104_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16840_ _16840_/A _16845_/C vssd1 vssd1 vccd1 vccd1 _16840_/Y sky130_fd_sc_hd__nor2_1
XFILLER_144_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16771_ _16848_/A vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__clkbuf_4
X_13983_ _18523_/Q _13981_/X _13995_/S vssd1 vssd1 vccd1 vccd1 _13984_/A sky130_fd_sc_hd__mux2_1
XFILLER_101_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15722_ _15722_/A vssd1 vssd1 vccd1 vccd1 _19206_/D sky130_fd_sc_hd__clkbuf_1
X_18510_ _19292_/CLK _18510_/D vssd1 vssd1 vccd1 vccd1 _18510_/Q sky130_fd_sc_hd__dfxtp_1
X_12934_ _19335_/Q _12600_/Y _13179_/A _19145_/Q vssd1 vssd1 vccd1 vccd1 _12934_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11845__A1 _11291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19490_ _19619_/CLK _19490_/D vssd1 vssd1 vccd1 vccd1 _19490_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_84_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _19384_/CLK _18441_/D vssd1 vssd1 vccd1 vccd1 _18441_/Q sky130_fd_sc_hd__dfxtp_1
X_15653_ _15653_/A vssd1 vssd1 vccd1 vccd1 _19175_/D sky130_fd_sc_hd__clkbuf_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _14531_/A vssd1 vssd1 vccd1 vccd1 _12865_/X sky130_fd_sc_hd__clkbuf_1
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14604_ _14604_/A vssd1 vssd1 vccd1 vccd1 _18772_/D sky130_fd_sc_hd__clkbuf_1
X_18372_ _19379_/CLK _18372_/D vssd1 vssd1 vccd1 vccd1 _18372_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11816_ _11842_/A _11842_/B _11842_/C _12050_/A vssd1 vssd1 vccd1 vccd1 _11817_/B
+ sky130_fd_sc_hd__a31o_1
X_15584_ _15583_/X _19159_/Q _15596_/S vssd1 vssd1 vccd1 vccd1 _15585_/A sky130_fd_sc_hd__mux2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12796_ _18744_/Q vssd1 vssd1 vccd1 vccd1 _13119_/A sky130_fd_sc_hd__inv_2
XFILLER_144_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17323_ _17530_/A vssd1 vssd1 vccd1 vccd1 _17419_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535_ _14534_/X _18751_/Q _14535_/S vssd1 vssd1 vccd1 vccd1 _14536_/A sky130_fd_sc_hd__mux2_1
XFILLER_30_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ _19635_/Q _13419_/A vssd1 vssd1 vccd1 vccd1 _11749_/A sky130_fd_sc_hd__or2b_1
XANTENNA__12270__A1 _19415_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14517__A _18163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15112__S _15112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_169_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17254_ _17251_/X _17344_/B _17336_/A vssd1 vssd1 vccd1 vccd1 _17435_/B sky130_fd_sc_hd__mux2_1
XFILLER_147_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14466_ _14466_/A vssd1 vssd1 vccd1 vccd1 _18718_/D sky130_fd_sc_hd__clkbuf_1
X_11678_ _11678_/A vssd1 vssd1 vccd1 vccd1 _11818_/S sky130_fd_sc_hd__buf_2
X_16205_ _13563_/X _19375_/Q _16213_/S vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__mux2_1
X_13417_ _12557_/X _13415_/X _13416_/Y _12575_/X _18253_/Q vssd1 vssd1 vccd1 vccd1
+ _13418_/B sky130_fd_sc_hd__a32o_4
XFILLER_139_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10629_ _10680_/A _10628_/X _09640_/X vssd1 vssd1 vccd1 vccd1 _10629_/Y sky130_fd_sc_hd__o21ai_1
X_17185_ _17185_/A _17185_/B vssd1 vssd1 vccd1 vccd1 _17432_/B sky130_fd_sc_hd__nor2_4
X_14397_ _14443_/S vssd1 vssd1 vccd1 vccd1 _14406_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__16732__A _16737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10033__B1 _09982_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16136_ _16135_/X _19353_/Q _16140_/S vssd1 vssd1 vccd1 vccd1 _16137_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13348_ _15092_/A vssd1 vssd1 vccd1 vccd1 _14614_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11781__B1 _11813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_154_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _16066_/X _19341_/Q _16083_/S vssd1 vssd1 vccd1 vccd1 _16068_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_13279_ _19765_/Q _13281_/B vssd1 vssd1 vccd1 vccd1 _13315_/C sky130_fd_sc_hd__and2_1
XFILLER_142_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_170_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09346__A _11618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ _15018_/A vssd1 vssd1 vccd1 vccd1 _18949_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_170_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_123_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19826_ _19830_/CLK _19826_/D vssd1 vssd1 vccd1 vccd1 _19826_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_111_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13286__B1 _13285_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19757_ _19793_/CLK _19757_/D vssd1 vssd1 vccd1 vccd1 _19757_/Q sky130_fd_sc_hd__dfxtp_1
X_16969_ _15522_/X _16956_/X _16967_/X _16968_/X vssd1 vssd1 vccd1 vccd1 _19641_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_110_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14398__S _14406_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09510_ _18642_/Q vssd1 vssd1 vccd1 vccd1 _09511_/A sky130_fd_sc_hd__buf_2
XANTENNA__15083__A _15083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18708_ _19006_/CLK _18708_/D vssd1 vssd1 vccd1 vccd1 _18708_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12500__A _12697_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19688_ _19688_/CLK _19688_/D vssd1 vssd1 vccd1 vccd1 _19688_/Q sky130_fd_sc_hd__dfxtp_1
X_09441_ _10670_/S vssd1 vssd1 vccd1 vccd1 _09441_/X sky130_fd_sc_hd__buf_4
X_18639_ _19296_/CLK _18639_/D vssd1 vssd1 vccd1 vccd1 _18639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11116__A _11116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_80_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _10949_/A vssd1 vssd1 vccd1 vccd1 _11307_/A sky130_fd_sc_hd__buf_2
XFILLER_21_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15957__S _15959_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10166__S _10166_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__A1 _19342_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_118_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_146_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09955__S _09955_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__B1 _09640_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_165_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_118_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_118_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13477__S _13481_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15258__A _15315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_161_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_88_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10327__A1 _09866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_88_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_102_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_106_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_87_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_114_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09708_ _09708_/A vssd1 vssd1 vccd1 vccd1 _10310_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14101__S _14107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10980_ _18455_/Q _19046_/Q _19208_/Q _18423_/Q _10862_/X _09513_/A vssd1 vssd1 vccd1
+ vccd1 _10981_/B sky130_fd_sc_hd__mux4_1
XFILLER_74_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _19296_/Q _19134_/Q _18543_/Q _18313_/Q _10572_/S _09542_/A vssd1 vssd1 vccd1
+ vccd1 _09639_/X sky130_fd_sc_hd__mux4_1
XANTENNA__16766__A1 _16772_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16817__A _16838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_71_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_128_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12650_ _12713_/A _18262_/Q vssd1 vssd1 vccd1 vccd1 _12650_/Y sky130_fd_sc_hd__nand2_1
XFILLER_70_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_169_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11601_ _11723_/S _12443_/B _11600_/Y vssd1 vssd1 vccd1 vccd1 _11716_/D sky130_fd_sc_hd__o21a_1
XFILLER_12_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _19621_/Q _12496_/C _12565_/X _16989_/A _12580_/X vssd1 vssd1 vccd1 vccd1
+ _12581_/X sky130_fd_sc_hd__a221o_1
XFILLER_12_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09653__C1 _10575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_168_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14320_ _14320_/A vssd1 vssd1 vccd1 vccd1 _18654_/D sky130_fd_sc_hd__clkbuf_1
X_11532_ _17183_/A _11564_/C _17174_/B _11532_/D vssd1 vssd1 vccd1 vccd1 _11533_/D
+ sky130_fd_sc_hd__or4_1
XFILLER_156_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_139_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14251_ _18632_/Q _14023_/X _14253_/S vssd1 vssd1 vccd1 vccd1 _14252_/A sky130_fd_sc_hd__mux2_1
X_11463_ _11463_/A _11463_/B _11463_/C vssd1 vssd1 vccd1 vccd1 _11463_/Y sky130_fd_sc_hd__nand3_1
XFILLER_87_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ _19541_/Q _12952_/X _12953_/X _19509_/Q _13201_/X vssd1 vssd1 vccd1 vccd1
+ _13202_/X sky130_fd_sc_hd__a221o_1
XFILLER_109_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_opt_4_0_clock clkbuf_4_13_0_clock/X vssd1 vssd1 vccd1 vccd1 clkbuf_opt_4_0_clock/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10414_ _10414_/A _10414_/B vssd1 vssd1 vccd1 vccd1 _10414_/X sky130_fd_sc_hd__and2_1
XFILLER_99_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_171_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14182_ _14182_/A vssd1 vssd1 vccd1 vccd1 _14191_/S sky130_fd_sc_hd__buf_4
X_11394_ _18416_/Q _18677_/Q _18576_/Q _18911_/Q _11388_/S _11389_/A vssd1 vssd1 vccd1
+ vccd1 _11394_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13387__S _13387_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_136_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _13360_/S _19724_/Q _13154_/A _13132_/X vssd1 vssd1 vccd1 vccd1 _13133_/X
+ sky130_fd_sc_hd__o211a_1
X_10345_ _10345_/A _10345_/B vssd1 vssd1 vccd1 vccd1 _10345_/Y sky130_fd_sc_hd__nor2_1
XFILLER_125_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10661__S1 _09707_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18990_ _18990_/CLK _18990_/D vssd1 vssd1 vccd1 vccd1 _18990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _17941_/A vssd1 vssd1 vccd1 vccd1 _19745_/D sky130_fd_sc_hd__clkbuf_1
X_13064_ _19751_/Q _19752_/Q _13064_/C vssd1 vssd1 vccd1 vccd1 _13083_/B sky130_fd_sc_hd__and3_1
XFILLER_79_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10276_ _18597_/Q _18868_/Q _19092_/Q _18836_/Q _10274_/X _10275_/X vssd1 vssd1 vccd1
+ vccd1 _10276_/X sky130_fd_sc_hd__mux4_1
XANTENNA_output156_A _12237_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_155_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10318__B2 _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12015_ _19645_/Q vssd1 vssd1 vccd1 vccd1 _16978_/A sky130_fd_sc_hd__clkbuf_2
X_17872_ _17592_/A _17870_/X _17871_/X _17596_/A _12317_/Y vssd1 vssd1 vccd1 vccd1
+ _17872_/X sky130_fd_sc_hd__a32o_2
XFILLER_79_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_2_1_0_clock_A clkbuf_2_1_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19611_ _19618_/CLK _19611_/D vssd1 vssd1 vccd1 vccd1 _19611_/Q sky130_fd_sc_hd__dfxtp_1
X_16823_ _19581_/Q _16824_/B vssd1 vssd1 vccd1 vccd1 _16825_/B sky130_fd_sc_hd__nor2_1
XFILLER_78_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11635__S _11678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19542_ _19543_/CLK _19542_/D vssd1 vssd1 vccd1 vccd1 _19542_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11818__A1 _10895_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16754_ _19553_/Q _19552_/Q _16754_/C _16754_/D vssd1 vssd1 vccd1 vccd1 _16760_/C
+ sky130_fd_sc_hd__and4_1
XANTENNA__14011__S _14011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13966_ _14049_/S vssd1 vssd1 vccd1 vccd1 _13979_/S sky130_fd_sc_hd__buf_2
XANTENNA__12320__A _12321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12917_ _19430_/Q _12700_/X _12916_/X vssd1 vssd1 vccd1 vccd1 _12917_/X sky130_fd_sc_hd__o21a_1
X_15705_ _15705_/A vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_74_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16685_ _16689_/C _16689_/D _16684_/Y vssd1 vssd1 vccd1 vccd1 _19537_/D sky130_fd_sc_hd__o21a_1
X_19473_ _19610_/CLK _19473_/D vssd1 vssd1 vccd1 vccd1 _19473_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16757__A1 _16760_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ _13896_/X _18498_/Q _13903_/S vssd1 vssd1 vccd1 vccd1 _13898_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18424_ _19241_/CLK _18424_/D vssd1 vssd1 vccd1 vccd1 _18424_/Q sky130_fd_sc_hd__dfxtp_1
X_15636_ _15635_/X _19169_/Q _15636_/S vssd1 vssd1 vccd1 vccd1 _15637_/A sky130_fd_sc_hd__mux2_1
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ _12848_/A _15998_/A vssd1 vssd1 vccd1 vccd1 _12848_/Y sky130_fd_sc_hd__nand2_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15567_ _15607_/A _18270_/Q vssd1 vssd1 vccd1 vccd1 _15567_/Y sky130_fd_sc_hd__nand2_1
X_18355_ _19300_/CLK _18355_/D vssd1 vssd1 vccd1 vccd1 _18355_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12779_ _12975_/B vssd1 vssd1 vccd1 vccd1 _12779_/Y sky130_fd_sc_hd__inv_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14518_ _16833_/A _14518_/B vssd1 vssd1 vccd1 vccd1 _18746_/D sky130_fd_sc_hd__nor2_1
X_17306_ _17396_/B vssd1 vssd1 vccd1 vccd1 _17457_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15498_ _15498_/A vssd1 vssd1 vccd1 vccd1 _19144_/D sky130_fd_sc_hd__clkbuf_1
X_18286_ _19237_/CLK _18286_/D vssd1 vssd1 vccd1 vccd1 _18286_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17182__A1 _11566_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10494__B _12464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14449_ _14449_/A vssd1 vssd1 vccd1 vccd1 _18710_/D sky130_fd_sc_hd__clkbuf_1
X_17237_ _17237_/A vssd1 vssd1 vccd1 vccd1 _17492_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14681__S _14687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_156_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11203__C1 _18782_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17168_ _17168_/A _17168_/B _17167_/X vssd1 vssd1 vccd1 vccd1 _17169_/D sky130_fd_sc_hd__or3b_1
XFILLER_127_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16119_ _16119_/A vssd1 vssd1 vccd1 vccd1 _16140_/S sky130_fd_sc_hd__clkbuf_2
X_17099_ _17099_/A vssd1 vssd1 vccd1 vccd1 _19695_/D sky130_fd_sc_hd__clkbuf_1
X_09990_ _09998_/A _09985_/X _09988_/X _09989_/X vssd1 vssd1 vccd1 vccd1 _09990_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10652__S1 _11298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15496__A1 _15495_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_170_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_142_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_124_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15806__A _15852_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_96_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19809_ _19838_/CLK _19809_/D vssd1 vssd1 vccd1 vccd1 _19809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16996__A1 _15574_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_111_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12230__A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14856__S _14858_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13760__S _13762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09424_ _10951_/A vssd1 vssd1 vccd1 vccd1 _10823_/A sky130_fd_sc_hd__buf_2
XFILLER_53_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ _12672_/A _13391_/C vssd1 vssd1 vccd1 vccd1 _16937_/D sky130_fd_sc_hd__nor2_1
XFILLER_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12785__A2 _12703_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_100_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09286_ _12543_/B _13400_/A _09285_/X vssd1 vssd1 vccd1 vccd1 _09301_/A sky130_fd_sc_hd__o21a_1
XFILLER_138_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_100_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_166_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15687__S _15693_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10891__S1 _10817_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16920__B2 _16932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_clock_A clkbuf_4_7_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_165_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_158_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10548__A1 _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_162_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17476__A2 _17430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12405__A _12405_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15487__B2 hold19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ _19289_/Q _19127_/Q _18536_/Q _18306_/Q _09918_/X _09900_/A vssd1 vssd1 vccd1
+ vccd1 _10130_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__13935__S _13935_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10061_ _18604_/Q _18875_/Q _19099_/Q _18843_/Q _09500_/A _10693_/A vssd1 vssd1 vccd1
+ vccd1 _10061_/X sky130_fd_sc_hd__mux4_1
XFILLER_88_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09714__A _09714_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13820_ _13251_/X _18473_/Q _13820_/S vssd1 vssd1 vccd1 vccd1 _13821_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ _13751_/A vssd1 vssd1 vccd1 vccd1 _18442_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14766__S _14770_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10963_ _10963_/A vssd1 vssd1 vccd1 vccd1 _10963_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ _19162_/Q _12895_/A _12640_/X _19352_/Q vssd1 vssd1 vccd1 vccd1 _12702_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16470_ _16470_/A _16474_/C vssd1 vssd1 vccd1 vccd1 _16470_/Y sky130_fd_sc_hd__nor2_1
X_13682_ _13311_/X _18412_/Q _13686_/S vssd1 vssd1 vccd1 vccd1 _13683_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10894_ _09431_/A _10887_/X _10889_/X _10893_/X _09614_/A vssd1 vssd1 vccd1 vccd1
+ _10894_/X sky130_fd_sc_hd__a311o_2
XFILLER_44_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15421_ _15421_/A vssd1 vssd1 vccd1 vccd1 _19117_/D sky130_fd_sc_hd__clkbuf_1
X_12633_ _13260_/A vssd1 vssd1 vccd1 vccd1 _12633_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_157_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18140_ _18140_/A _18146_/B vssd1 vssd1 vccd1 vccd1 _18140_/X sky130_fd_sc_hd__or2_1
X_15352_ _15374_/A vssd1 vssd1 vccd1 vccd1 _15361_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12776__A2 _12773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12564_ _19569_/Q vssd1 vssd1 vccd1 vccd1 _16790_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_12_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_169_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10787__A1 _09651_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14303_ _14303_/A vssd1 vssd1 vccd1 vccd1 _18646_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_12_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18071_ _09236_/C _19804_/Q _18071_/S vssd1 vssd1 vccd1 vccd1 _18072_/B sky130_fd_sc_hd__mux2_1
X_11515_ _11530_/A _17108_/B _17108_/A vssd1 vssd1 vccd1 vccd1 _11562_/A sky130_fd_sc_hd__a21oi_1
X_15283_ _14573_/X _19056_/Q _15289_/S vssd1 vssd1 vccd1 vccd1 _15284_/A sky130_fd_sc_hd__mux2_1
X_12495_ _16937_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _12496_/C sky130_fd_sc_hd__nor2_2
X_17022_ _15631_/X _17010_/X _17020_/X _17021_/X vssd1 vssd1 vccd1 vccd1 _19661_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_156_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14234_ _18624_/Q _13997_/X _14242_/S vssd1 vssd1 vccd1 vccd1 _14235_/A sky130_fd_sc_hd__mux2_1
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11446_ _11446_/A _11446_/B vssd1 vssd1 vccd1 vccd1 _11446_/Y sky130_fd_sc_hd__nand2_1
XFILLER_109_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_109_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14165_ _18594_/Q _14004_/X _14169_/S vssd1 vssd1 vccd1 vccd1 _14166_/A sky130_fd_sc_hd__mux2_1
XFILLER_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11377_ _09687_/A _11374_/X _11376_/X vssd1 vssd1 vccd1 vccd1 _11377_/X sky130_fd_sc_hd__a21o_1
XFILLER_153_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_152_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_140_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _13132_/A _12542_/B _12542_/C _13115_/X _13234_/A vssd1 vssd1 vccd1 vccd1
+ _13116_/X sky130_fd_sc_hd__o311a_1
X_10328_ _09844_/A _10321_/X _10323_/X _10327_/X _09754_/A vssd1 vssd1 vccd1 vccd1
+ _10328_/X sky130_fd_sc_hd__a311o_4
XFILLER_125_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_124_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _13902_/X _18564_/Q _14096_/S vssd1 vssd1 vccd1 vccd1 _14097_/A sky130_fd_sc_hd__mux2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _19292_/CLK _18973_/D vssd1 vssd1 vccd1 vccd1 _18973_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _15038_/A vssd1 vssd1 vccd1 vccd1 _14560_/A sky130_fd_sc_hd__clkbuf_2
X_17924_ _12432_/Y _17786_/A _17923_/X _12744_/A vssd1 vssd1 vccd1 vccd1 _17924_/X
+ sky130_fd_sc_hd__a211o_1
X_10259_ _10485_/A vssd1 vssd1 vccd1 vccd1 _10378_/A sky130_fd_sc_hd__buf_2
XFILLER_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09624__A _09624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11873__B _17195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17855_ _17853_/X _17854_/Y _17855_/S vssd1 vssd1 vccd1 vccd1 _17855_/X sky130_fd_sc_hd__mux2_1
XFILLER_94_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16806_ _16806_/A vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__buf_2
XANTENNA__09343__B _19844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12050__A _12050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17786_ _17786_/A vssd1 vssd1 vccd1 vccd1 _17786_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14998_ _14998_/A _14998_/B vssd1 vssd1 vccd1 vccd1 _15080_/A sky130_fd_sc_hd__and2_2
XFILLER_19_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19525_ _19529_/CLK _19525_/D vssd1 vssd1 vccd1 vccd1 _19525_/Q sky130_fd_sc_hd__dfxtp_1
X_16737_ _16737_/A _16737_/B _16741_/C vssd1 vssd1 vccd1 vccd1 _19555_/D sky130_fd_sc_hd__nor3_1
XANTENNA__14676__S _14676_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13949_ _14030_/A vssd1 vssd1 vccd1 vccd1 _14049_/S sky130_fd_sc_hd__buf_8
XFILLER_19_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_clock_A clkbuf_3_5_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19456_ _19594_/CLK _19456_/D vssd1 vssd1 vccd1 vccd1 _19456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16668_ _19532_/Q _16668_/B vssd1 vssd1 vccd1 vccd1 _16670_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18407_ _18902_/CLK _18407_/D vssd1 vssd1 vccd1 vccd1 _18407_/Q sky130_fd_sc_hd__dfxtp_1
X_15619_ _13325_/X _15613_/Y _18279_/Q vssd1 vssd1 vccd1 vccd1 _15619_/X sky130_fd_sc_hd__mux2_1
X_19387_ _19387_/CLK _19387_/D vssd1 vssd1 vccd1 vccd1 _19387_/Q sky130_fd_sc_hd__dfxtp_1
X_16599_ _16610_/A _16604_/C vssd1 vssd1 vccd1 vccd1 _16599_/Y sky130_fd_sc_hd__nor2_1
X_09140_ _09142_/A _09167_/B _09338_/C vssd1 vssd1 vccd1 vccd1 _11589_/A sky130_fd_sc_hd__or3_2
X_18338_ _19284_/CLK _18338_/D vssd1 vssd1 vccd1 vccd1 _18338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_148_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10322__S0 _09682_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__A1 _19113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18269_ _19162_/CLK _18269_/D vssd1 vssd1 vccd1 vccd1 _18269_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15300__S _15300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_129_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_147_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_116_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_104_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_115_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09973_ _09762_/A _09962_/X _09971_/X _09835_/A _09972_/Y vssd1 vssd1 vccd1 vccd1
+ _12473_/B sky130_fd_sc_hd__o32a_4
XFILLER_131_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_162_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10389__S0 _10274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_112_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09534__A _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16969__A1 _15522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15970__S _15970_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13490__S _13492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_164_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10561__S0 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09407_ _09688_/A _09400_/X _10046_/A vssd1 vssd1 vccd1 vccd1 _09407_/X sky130_fd_sc_hd__a21o_1
XFILLER_164_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12207__A1 _19413_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12758__A2 _12752_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ _18130_/A _11522_/A _09338_/C _11522_/C vssd1 vssd1 vccd1 vccd1 _17126_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA__17146__A1 _19701_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_139_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11966__B1 _16114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17146__B2 _18099_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17198__A _17198_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ _12584_/A _12605_/A vssd1 vssd1 vccd1 vccd1 _12956_/A sky130_fd_sc_hd__or2_2
XFILLER_154_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_126_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _09394_/A _11299_/X _10547_/A vssd1 vssd1 vccd1 vccd1 _11300_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09709__A _10310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _18132_/A _11516_/A _12302_/A vssd1 vssd1 vccd1 vccd1 _12280_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_101_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_119_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11231_ _19267_/Q _19105_/Q _18514_/Q _18284_/Q _11265_/S _10971_/A vssd1 vssd1 vccd1
+ vccd1 _11232_/B sky130_fd_sc_hd__mux4_1
XFILLER_134_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_150_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11162_ _11164_/A _11161_/X _09561_/A vssd1 vssd1 vccd1 vccd1 _11162_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_171_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_161_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10941__A1 _09393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_171_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10113_ _10113_/A vssd1 vssd1 vccd1 vccd1 _10113_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15446__A _15446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15970_ _13576_/X _19317_/Q _15970_/S vssd1 vssd1 vccd1 vccd1 _15971_/A sky130_fd_sc_hd__mux2_1
XFILLER_121_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11093_ _19711_/Q vssd1 vssd1 vccd1 vccd1 _11093_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12143__A0 _19790_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input32_A io_dbus_rdata[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_121_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14921_ _14921_/A vssd1 vssd1 vccd1 vccd1 _18906_/D sky130_fd_sc_hd__clkbuf_1
X_10044_ _10046_/A _10043_/X _09434_/A vssd1 vssd1 vccd1 vccd1 _10044_/X sky130_fd_sc_hd__o21a_1
XFILLER_102_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_130_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_102_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17640_ _17642_/A _17642_/B vssd1 vssd1 vccd1 vccd1 _17640_/Y sky130_fd_sc_hd__nand2_1
XFILLER_36_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14852_ _18876_/Q _14039_/X _14854_/S vssd1 vssd1 vccd1 vccd1 _14853_/A sky130_fd_sc_hd__mux2_1
XANTENNA__15632__A1 _15631_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13803_ _13124_/X _18465_/Q _13809_/S vssd1 vssd1 vccd1 vccd1 _13804_/A sky130_fd_sc_hd__mux2_1
XANTENNA__14496__S _14500_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17571_ _17571_/A vssd1 vssd1 vccd1 vccd1 _17571_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_14783_ _14617_/X _18846_/Q _14785_/S vssd1 vssd1 vccd1 vccd1 _14784_/A sky130_fd_sc_hd__mux2_1
X_11995_ _12230_/A _11993_/Y _12044_/C _11962_/A vssd1 vssd1 vccd1 vccd1 _11995_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_44_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_91_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19310_ _19310_/CLK _19310_/D vssd1 vssd1 vccd1 vccd1 _19310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13734_ _13148_/X _18435_/Q _13736_/S vssd1 vssd1 vccd1 vccd1 _13735_/A sky130_fd_sc_hd__mux2_1
X_16522_ _19489_/Q _19488_/Q _19619_/Q _16522_/D vssd1 vssd1 vccd1 vccd1 _16533_/D
+ sky130_fd_sc_hd__and4_1
X_10946_ _18391_/Q _18652_/Q _18551_/Q _18886_/Q _11050_/S _10934_/A vssd1 vssd1 vccd1
+ vccd1 _10947_/B sky130_fd_sc_hd__mux4_1
XFILLER_90_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10552__S0 _10542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_91_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19241_ _19241_/CLK _19241_/D vssd1 vssd1 vccd1 vccd1 _19241_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ _13665_/A vssd1 vssd1 vccd1 vccd1 _18404_/D sky130_fd_sc_hd__clkbuf_1
X_16453_ _16453_/A vssd1 vssd1 vccd1 vccd1 _16458_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_10877_ _09705_/A _10872_/X _10876_/X vssd1 vssd1 vccd1 vccd1 _10877_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13946__A1 _16619_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12616_ _13397_/A _12615_/Y _12714_/A vssd1 vssd1 vccd1 vccd1 _12616_/X sky130_fd_sc_hd__a21o_1
X_15404_ _15404_/A vssd1 vssd1 vccd1 vccd1 _19109_/D sky130_fd_sc_hd__clkbuf_1
X_16384_ _19444_/Q _16387_/C _16359_/X vssd1 vssd1 vccd1 vccd1 _16384_/Y sky130_fd_sc_hd__a21oi_1
X_19172_ _19202_/CLK _19172_/D vssd1 vssd1 vccd1 vccd1 _19172_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__17137__A1 _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13596_ _13596_/A vssd1 vssd1 vccd1 vccd1 _13609_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__17137__B2 _12543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12029__B _17211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18123_ _18136_/A vssd1 vssd1 vccd1 vccd1 _18123_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15335_ _19079_/Q _15022_/X _15339_/S vssd1 vssd1 vccd1 vccd1 _15336_/A sky130_fd_sc_hd__mux2_1
X_12547_ _12713_/A hold8/A vssd1 vssd1 vccd1 vccd1 _12547_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16216__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_118_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15266_ _15266_/A vssd1 vssd1 vccd1 vccd1 _19048_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09619__A _09644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18054_ _18054_/A vssd1 vssd1 vccd1 vccd1 _19796_/D sky130_fd_sc_hd__clkbuf_1
X_12478_ _12480_/A _12478_/B vssd1 vssd1 vccd1 vccd1 _12478_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_126_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17005_ _17005_/A _17011_/B vssd1 vssd1 vccd1 vccd1 _17005_/X sky130_fd_sc_hd__or2_1
X_14217_ _14217_/A vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__18098__C1 _18097_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_11429_ _11431_/A _11433_/A _11431_/C _12473_/B _10087_/A vssd1 vssd1 vccd1 vccd1
+ _11429_/X sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_4_12_0_clock_A clkbuf_3_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10607__S1 _09590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15197_ _15243_/S vssd1 vssd1 vccd1 vccd1 _15206_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_99_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_153_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _14148_/A vssd1 vssd1 vccd1 vccd1 _18586_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10932__A1 _09477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_113_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14079_ _13877_/X _18556_/Q _14085_/S vssd1 vssd1 vccd1 vccd1 _14080_/A sky130_fd_sc_hd__mux2_1
X_18956_ _19098_/CLK _18956_/D vssd1 vssd1 vccd1 vccd1 _18956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_67_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09354__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ _17907_/A _17907_/B vssd1 vssd1 vccd1 vccd1 _17907_/X sky130_fd_sc_hd__or2_1
XFILLER_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18887_ _19365_/CLK _18887_/D vssd1 vssd1 vccd1 vccd1 _18887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09550__A1 _09803_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17838_ _17390_/A _17624_/X _17837_/X _17633_/X vssd1 vssd1 vccd1 vccd1 _17838_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_67_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12437__A1 _11686_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17769_ _17920_/B _17764_/X _17768_/X _17478_/A vssd1 vssd1 vccd1 vccd1 _17769_/X
+ sky130_fd_sc_hd__a211o_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19508_ _19540_/CLK _19508_/D vssd1 vssd1 vccd1 vccd1 _19508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10543__S0 _10763_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19439_ _19583_/CLK _19439_/D vssd1 vssd1 vccd1 vccd1 _19439_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16915__A _16915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17128__A1 _17114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_9_0_clock_A clkbuf_4_9_0_clock/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ _09325_/A _11528_/A _09146_/C _11646_/B vssd1 vssd1 vccd1 vccd1 _09124_/B
+ sky130_fd_sc_hd__or4_4
XFILLER_163_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_132_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12373__B1 _15632_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_173_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_106_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09956_ _09956_/A _09956_/B vssd1 vssd1 vccd1 vccd1 _09956_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17851__A2 _12727_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09887_ _10342_/A vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__buf_2
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_100_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_100_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12829__S _12887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18159__A3 _18066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ _11124_/A vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__buf_2
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _19397_/Q _11640_/X _11772_/X _11779_/X vssd1 vssd1 vccd1 vccd1 _16253_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10534__S0 _10433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _09394_/A _10730_/X _09596_/A vssd1 vssd1 vccd1 vccd1 _10731_/X sky130_fd_sc_hd__a21o_1
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16825__A _16838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13450_ _13507_/S vssd1 vssd1 vccd1 vccd1 _13459_/S sky130_fd_sc_hd__buf_2
XFILLER_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10662_ _09597_/X _10661_/X _09602_/X vssd1 vssd1 vccd1 vccd1 _10662_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17119__A1 _17114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_167_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_167_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12401_ _17899_/A vssd1 vssd1 vccd1 vccd1 _12401_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11969__A _19402_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13381_ _19738_/Q _13380_/X _13381_/S vssd1 vssd1 vccd1 vccd1 _13381_/X sky130_fd_sc_hd__mux2_1
X_10593_ _10585_/Y _10588_/Y _10590_/Y _10592_/Y _09572_/A vssd1 vssd1 vccd1 vccd1
+ _10593_/X sky130_fd_sc_hd__o221a_4
XFILLER_51_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_139_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _15120_/A vssd1 vssd1 vccd1 vccd1 _18983_/D sky130_fd_sc_hd__clkbuf_1
X_12332_ _17878_/A _12332_/B vssd1 vssd1 vccd1 vccd1 _12351_/A sky130_fd_sc_hd__xnor2_4
XFILLER_126_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_127_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15051_ _15051_/A vssd1 vssd1 vccd1 vccd1 _15051_/X sky130_fd_sc_hd__clkbuf_2
X_12263_ _17845_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12265_/A sky130_fd_sc_hd__xnor2_4
XFILLER_142_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14002_ _18529_/Q _14001_/X _14011_/S vssd1 vssd1 vccd1 vccd1 _14003_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09455__S1 _09390_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_135_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11214_ _09366_/A _11204_/X _11213_/X _09469_/A _19708_/Q vssd1 vssd1 vccd1 vccd1
+ _11239_/A sky130_fd_sc_hd__a32o_2
XANTENNA__18095__A2 _18086_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12194_ _12196_/A _12195_/A vssd1 vssd1 vccd1 vccd1 _12223_/A sky130_fd_sc_hd__or2_1
XANTENNA__10375__C1 _09669_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_150_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18810_ _19386_/CLK _18810_/D vssd1 vssd1 vccd1 vccd1 _18810_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_122_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11145_ _10943_/X _11138_/X _11140_/X _11144_/X _09465_/A vssd1 vssd1 vccd1 vccd1
+ _11145_/X sky130_fd_sc_hd__a311o_1
Xoutput73 _11932_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[11] sky130_fd_sc_hd__buf_2
Xoutput84 _12200_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[21] sky130_fd_sc_hd__buf_2
X_19790_ _19800_/CLK _19790_/D vssd1 vssd1 vccd1 vccd1 _19790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_123_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput95 _12432_/Y vssd1 vssd1 vccd1 vccd1 io_dbus_addr[31] sky130_fd_sc_hd__buf_2
X_18741_ _19071_/CLK _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13408__B _13408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15953_ _13551_/X _19309_/Q _15959_/S vssd1 vssd1 vccd1 vccd1 _15954_/A sky130_fd_sc_hd__mux2_1
X_11076_ _18916_/Q _18682_/Q _19364_/Q _19012_/Q _11265_/S _11033_/A vssd1 vssd1 vccd1
+ vccd1 _11077_/B sky130_fd_sc_hd__mux4_1
XFILLER_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14904_ _18899_/Q _14010_/X _14904_/S vssd1 vssd1 vccd1 vccd1 _14905_/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_1_clock_A clkbuf_4_0_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ _19733_/Q vssd1 vssd1 vccd1 vccd1 _10027_/Y sky130_fd_sc_hd__inv_2
XFILLER_64_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18672_ _18990_/CLK _18672_/D vssd1 vssd1 vccd1 vccd1 _18672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15884_ _15884_/A vssd1 vssd1 vccd1 vccd1 _19278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_76_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_91_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17623_ _17281_/X _17229_/X _17738_/S vssd1 vssd1 vccd1 vccd1 _17623_/X sky130_fd_sc_hd__mux2_1
X_14835_ _18868_/Q _14013_/X _14843_/S vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17554_ _17653_/A _17551_/X _17553_/X vssd1 vssd1 vccd1 vccd1 _17554_/X sky130_fd_sc_hd__o21ba_1
XFILLER_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14766_ _14592_/X _18838_/Q _14770_/S vssd1 vssd1 vccd1 vccd1 _14767_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11978_ _12025_/C vssd1 vssd1 vccd1 vccd1 _17709_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__10525__S0 _10433_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ _19486_/Q _16503_/B _16504_/Y vssd1 vssd1 vccd1 vccd1 _19486_/D sky130_fd_sc_hd__o21a_1
XFILLER_16_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13717_ _13025_/X _18427_/Q _13725_/S vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__mux2_1
X_10929_ _10929_/A vssd1 vssd1 vccd1 vccd1 _11044_/A sky130_fd_sc_hd__clkbuf_2
X_14697_ _14697_/A vssd1 vssd1 vccd1 vccd1 _18807_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17485_ _17485_/A vssd1 vssd1 vccd1 vccd1 _17896_/S sky130_fd_sc_hd__buf_2
X_19224_ _19471_/CLK _19224_/D vssd1 vssd1 vccd1 vccd1 _19224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16436_ _16470_/A _16440_/C vssd1 vssd1 vccd1 vccd1 _16436_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13648_ _13648_/A vssd1 vssd1 vccd1 vccd1 _18396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11879__A _11879_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _19688_/CLK _19155_/D vssd1 vssd1 vccd1 vccd1 _19155_/Q sky130_fd_sc_hd__dfxtp_1
X_16367_ _19437_/Q _16365_/B _16366_/Y vssd1 vssd1 vccd1 vccd1 _19437_/D sky130_fd_sc_hd__o21a_1
X_13579_ _15063_/A vssd1 vssd1 vccd1 vccd1 _13579_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__10828__S1 _10802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_173_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18106_ _18134_/A vssd1 vssd1 vccd1 vccd1 _18106_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_118_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09349__A _19863_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15318_ _15374_/A vssd1 vssd1 vccd1 vccd1 _15387_/S sky130_fd_sc_hd__buf_6
XFILLER_157_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16298_ _16298_/A _16298_/B vssd1 vssd1 vccd1 vccd1 _16299_/A sky130_fd_sc_hd__and2_1
X_19086_ _19086_/CLK _19086_/D vssd1 vssd1 vccd1 vccd1 _19086_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_173_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_172_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__15785__S _15793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18037_ _18037_/A vssd1 vssd1 vccd1 vccd1 _19789_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_172_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15249_ _15249_/A vssd1 vssd1 vccd1 vccd1 _19040_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_114_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_99_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09783__S _09786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_125_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_114_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09810_ _09817_/A _09802_/X _09809_/X vssd1 vssd1 vccd1 vccd1 _09810_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15086__A _15086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_141_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09741_ _11368_/A _09734_/X _09736_/X _09740_/X vssd1 vssd1 vccd1 vccd1 _09742_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_101_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13855__A0 _13854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18939_ _18987_/CLK _18939_/D vssd1 vssd1 vccd1 vccd1 _18939_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_95_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09672_ _09672_/A vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__buf_2
XFILLER_95_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09812__A _09812_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_168_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11633__A2 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_74_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15780__A0 _13614_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_109_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10693__A _10693_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_148_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _09174_/B vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_164_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18071__S _18071_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_104_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12897__A1 _19143_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__B2 _19333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_132_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_105_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17285__A0 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_89_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14099__A0 _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17824__A2 _17819_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_131_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09939_ _09844_/X _09929_/X _09933_/X _09938_/X _09670_/A vssd1 vssd1 vccd1 vccd1
+ _09939_/X sky130_fd_sc_hd__a311o_2
XANTENNA__10109__C1 _09740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13846__A0 _13845_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _13260_/A vssd1 vssd1 vccd1 vccd1 _12950_/X sky130_fd_sc_hd__clkbuf_2
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18100__A _18100_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_93_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _11848_/A _11872_/X _11874_/B vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__o21a_1
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09722__A _10200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12881_ _13114_/A vssd1 vssd1 vccd1 vccd1 _13103_/S sky130_fd_sc_hd__clkbuf_2
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11832_ _19638_/Q _11832_/B vssd1 vssd1 vccd1 vccd1 _11886_/C sky130_fd_sc_hd__and2_1
X_14620_ _14620_/A vssd1 vssd1 vccd1 vccd1 _14620_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_73_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14551_ _14550_/X _18756_/Q _14551_/S vssd1 vssd1 vccd1 vccd1 _14552_/A sky130_fd_sc_hd__mux2_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ _11788_/A _11788_/B _11729_/A vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__a21bo_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _10719_/A _10714_/B vssd1 vssd1 vccd1 vccd1 _10714_/Y sky130_fd_sc_hd__nor2_1
X_13502_ _13502_/A vssd1 vssd1 vccd1 vccd1 _18349_/D sky130_fd_sc_hd__clkbuf_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14482_ _14482_/A vssd1 vssd1 vccd1 vccd1 _18725_/D sky130_fd_sc_hd__clkbuf_1
X_17270_ _12245_/A _17630_/B _17283_/S vssd1 vssd1 vccd1 vccd1 _17270_/X sky130_fd_sc_hd__mux2_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ _19633_/Q vssd1 vssd1 vccd1 vccd1 _16947_/A sky130_fd_sc_hd__inv_2
XFILLER_14_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16221_ _16221_/A vssd1 vssd1 vccd1 vccd1 _19382_/D sky130_fd_sc_hd__clkbuf_1
X_13433_ _13619_/A vssd1 vssd1 vccd1 vccd1 _18096_/A sky130_fd_sc_hd__buf_6
XFILLER_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10645_ _19719_/Q vssd1 vssd1 vccd1 vccd1 _10645_/Y sky130_fd_sc_hd__inv_2
X_16152_ _16114_/X _15620_/X _16151_/Y vssd1 vssd1 vccd1 vccd1 _16152_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13364_ _13154_/X _13360_/X _13363_/X vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__a21oi_1
X_10576_ _10631_/S vssd1 vssd1 vccd1 vccd1 _10576_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_154_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_80_clock_A _19161_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15103_ _15171_/S vssd1 vssd1 vccd1 vccd1 _15112_/S sky130_fd_sc_hd__clkbuf_4
X_12315_ _12267_/A _12267_/B _12312_/Y _12314_/Y vssd1 vssd1 vccd1 vccd1 _12316_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_154_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16083_ _16082_/X _19344_/Q _16083_/S vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_115_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13295_ _13294_/X _18309_/Q _13350_/S vssd1 vssd1 vccd1 vccd1 _13296_/A sky130_fd_sc_hd__mux2_1
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15034_ _15034_/A vssd1 vssd1 vccd1 vccd1 _18954_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12246_ _12248_/A _17835_/B vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__or2_1
XFILLER_142_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17276__A0 _17802_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_123_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_122_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19842_ _19865_/CLK _19842_/D vssd1 vssd1 vccd1 vccd1 _19842_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12177_ _19410_/Q _19411_/Q _19412_/Q _12177_/D vssd1 vssd1 vccd1 vccd1 _12201_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_111_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10994__S0 _11050_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11128_ _18483_/Q _18978_/Q _11128_/S vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__mux2_1
XFILLER_68_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19773_ _19786_/CLK _19773_/D vssd1 vssd1 vccd1 vccd1 _19773_/Q sky130_fd_sc_hd__dfxtp_1
X_16985_ _12550_/X _16983_/X _16984_/X _16981_/X vssd1 vssd1 vccd1 vccd1 _19647_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_95_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_110_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18724_ _19312_/CLK _18724_/D vssd1 vssd1 vccd1 vccd1 _18724_/Q sky130_fd_sc_hd__dfxtp_1
X_11059_ _11171_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11059_/X sky130_fd_sc_hd__or2_1
X_15936_ _15936_/A vssd1 vssd1 vccd1 vccd1 _19301_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_97_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09632__A _09632_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18655_ _19308_/CLK _18655_/D vssd1 vssd1 vccd1 vccd1 _18655_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15867_ _15924_/S vssd1 vssd1 vccd1 vccd1 _15876_/S sky130_fd_sc_hd__buf_2
XFILLER_36_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17606_ _17910_/A _17601_/Y _17605_/Y vssd1 vssd1 vccd1 vccd1 _17606_/Y sky130_fd_sc_hd__a21oi_1
X_14818_ _14818_/A vssd1 vssd1 vccd1 vccd1 _18860_/D sky130_fd_sc_hd__clkbuf_1
X_18586_ _19081_/CLK _18586_/D vssd1 vssd1 vccd1 vccd1 _18586_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_91_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15798_ _13535_/X _19240_/Q _15804_/S vssd1 vssd1 vccd1 vccd1 _15799_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17537_ _17626_/A vssd1 vssd1 vccd1 vccd1 _17537_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14749_ _14749_/A vssd1 vssd1 vccd1 vccd1 _18830_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17468_ _17468_/A _17468_/B vssd1 vssd1 vccd1 vccd1 _17468_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_149_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19207_ _19239_/CLK _19207_/D vssd1 vssd1 vccd1 vccd1 _19207_/Q sky130_fd_sc_hd__dfxtp_1
X_16419_ _19456_/Q vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_182_clock clkbuf_4_2_0_clock/X vssd1 vssd1 vccd1 vccd1 _19239_/CLK sky130_fd_sc_hd__clkbuf_16
X_17399_ _17573_/S _17457_/B vssd1 vssd1 vccd1 vccd1 _17399_/Y sky130_fd_sc_hd__nor2_2
XFILLER_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19138_ _19667_/CLK _19138_/D vssd1 vssd1 vccd1 vccd1 _19138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09079__A _09166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_157_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_145_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_146_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_118_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19069_ _19375_/CLK _19069_/D vssd1 vssd1 vccd1 vccd1 _19069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_146_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10018__A _10261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_173_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_161_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09807__A _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_172_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13329__A _15089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12233__A _16114_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10354__A2 _10338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_120_clock clkbuf_opt_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19865_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__17743__B _17743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09724_ _10108_/A vssd1 vssd1 vccd1 vccd1 _11380_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_101_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_170_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09542__A _09542_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_67_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09655_ _18607_/Q _18878_/Q _19102_/Q _18846_/Q _10785_/S _10586_/A vssd1 vssd1 vccd1
+ vccd1 _09655_/X sky130_fd_sc_hd__mux4_1
XFILLER_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_135_clock clkbuf_4_11_0_clock/X vssd1 vssd1 vccd1 vccd1 _19779_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _18942_/Q _18708_/Q _19390_/Q _19038_/Q _10030_/S _10669_/A vssd1 vssd1 vccd1
+ vccd1 _09586_/X sky130_fd_sc_hd__mux4_1
XFILLER_83_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18066__S _18066_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_169_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17742__A1 _17743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_102_clock_A _19586_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ _18466_/Q _19057_/Q _19219_/Q _18434_/Q _10339_/S _10270_/A vssd1 vssd1 vccd1
+ vccd1 _10430_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13938__S _13941_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09983__A1 _09688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _10361_/A _10361_/B vssd1 vssd1 vccd1 vccd1 _10361_/X sky130_fd_sc_hd__or2_1
XFILLER_136_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_164_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_152_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_151_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12100_ _12100_/A vssd1 vssd1 vccd1 vccd1 _12341_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13080_ _16681_/C _12782_/X _12635_/X hold1/A _13079_/X vssd1 vssd1 vccd1 vccd1 _13080_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_152_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10292_ _10394_/A _10291_/X _09822_/A vssd1 vssd1 vccd1 vccd1 _10292_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_151_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11781__A2_N _12449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12031_ _12031_/A _17211_/A vssd1 vssd1 vccd1 vccd1 _12032_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13239__A _15073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_160_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10976__S0 _10862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_77_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_1_1_0_clock_A clkbuf_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13673__S _13675_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16770_ _16799_/A _16770_/B _16770_/C vssd1 vssd1 vccd1 vccd1 _19564_/D sky130_fd_sc_hd__nor3_1
XANTENNA__14492__A0 _13905_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13982_ _14049_/S vssd1 vssd1 vccd1 vccd1 _13995_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_19_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_74_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ _13528_/X _19206_/Q _15721_/S vssd1 vssd1 vccd1 vccd1 _15722_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09594__S0 _10603_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09452__A _10040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_92_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12933_ _19671_/Q _13008_/A _12660_/B _19624_/Q _12932_/X vssd1 vssd1 vccd1 vccd1
+ _12933_/X sky130_fd_sc_hd__a221o_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_27_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _19382_/CLK _18440_/D vssd1 vssd1 vccd1 vccd1 _18440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15652_ _14537_/X _19175_/Q _15660_/S vssd1 vssd1 vccd1 vccd1 _15653_/A sky130_fd_sc_hd__mux2_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _15009_/A vssd1 vssd1 vccd1 vccd1 _14531_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14603_ _14601_/X _18772_/Q _14615_/S vssd1 vssd1 vccd1 vccd1 _14604_/A sky130_fd_sc_hd__mux2_1
X_18371_ _19378_/CLK _18371_/D vssd1 vssd1 vccd1 vccd1 _18371_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _17587_/A vssd1 vssd1 vccd1 vccd1 _11842_/B sky130_fd_sc_hd__inv_2
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15583_ _19728_/Q _15582_/X _15595_/S vssd1 vssd1 vccd1 vccd1 _15583_/X sky130_fd_sc_hd__mux2_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output101_A _11855_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12795_ _19739_/Q _12792_/X _13144_/S vssd1 vssd1 vccd1 vccd1 _12795_/X sky130_fd_sc_hd__mux2_2
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16285__A _16301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17322_ _17404_/C _17404_/A _17319_/B vssd1 vssd1 vccd1 vccd1 _17530_/A sky130_fd_sc_hd__or3b_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ _11746_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _13419_/A sky130_fd_sc_hd__nor2_1
XFILLER_144_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14534_ _14534_/A vssd1 vssd1 vccd1 vccd1 _14534_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_42_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_147_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17253_ _17252_/X _12349_/A _17261_/S vssd1 vssd1 vccd1 vccd1 _17344_/B sky130_fd_sc_hd__mux2_1
XFILLER_174_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14465_ _13867_/X _18718_/Q _14467_/S vssd1 vssd1 vccd1 vccd1 _14466_/A sky130_fd_sc_hd__mux2_1
X_11677_ _09665_/A _11182_/X _11191_/X _09756_/A _19710_/Q vssd1 vssd1 vccd1 vccd1
+ _11677_/X sky130_fd_sc_hd__a32o_2
XFILLER_169_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_146_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ _16226_/A vssd1 vssd1 vccd1 vccd1 _16213_/S sky130_fd_sc_hd__buf_4
X_13416_ _15599_/A _18253_/Q vssd1 vssd1 vccd1 vccd1 _13416_/Y sky130_fd_sc_hd__nand2_1
X_10628_ _19278_/Q _19116_/Q _18525_/Q _18295_/Q _10055_/S _11321_/A vssd1 vssd1 vccd1
+ vccd1 _10628_/X sky130_fd_sc_hd__mux4_1
XFILLER_174_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14396_ _14396_/A vssd1 vssd1 vccd1 vccd1 _18687_/D sky130_fd_sc_hd__clkbuf_1
X_17184_ _17184_/A _17184_/B _17184_/C _11542_/A vssd1 vssd1 vccd1 vccd1 _17185_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_139_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_127_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16135_ _16114_/X _15600_/X _16134_/Y vssd1 vssd1 vccd1 vccd1 _16135_/X sky130_fd_sc_hd__a21o_1
X_13347_ _12855_/X _13333_/X _13337_/Y _13346_/X vssd1 vssd1 vccd1 vccd1 _15092_/A
+ sky130_fd_sc_hd__a22o_4
XFILLER_154_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10559_ _10559_/A _10559_/B vssd1 vssd1 vccd1 vccd1 _10559_/X sky130_fd_sc_hd__or2_1
XANTENNA__16224__S _16224_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11781__B2 _18135_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09627__A _09645_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16066_ _15536_/X _16065_/Y _16082_/S vssd1 vssd1 vccd1 vccd1 _16066_/X sky130_fd_sc_hd__mux2_1
X_13278_ input19/X _13134_/X _13254_/X vssd1 vssd1 vccd1 vccd1 _13278_/X sky130_fd_sc_hd__a21o_1
XFILLER_64_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_97_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12229_ _12392_/S _12229_/B _12271_/C vssd1 vssd1 vccd1 vccd1 _12229_/X sky130_fd_sc_hd__or3_1
X_15017_ _18949_/Q _15015_/X _15029_/S vssd1 vssd1 vccd1 vccd1 _15018_/A sky130_fd_sc_hd__mux2_1
XANTENNA__09346__B _11619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__10967__S0 _10862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19825_ _19828_/CLK _19825_/D vssd1 vssd1 vccd1 vccd1 _19825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_151_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14679__S _14687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19756_ _19756_/CLK _19756_/D vssd1 vssd1 vccd1 vccd1 _19756_/Q sky130_fd_sc_hd__dfxtp_1
X_16968_ _16981_/A vssd1 vssd1 vccd1 vccd1 _16968_/X sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_52_clock clkbuf_4_5_0_clock/X vssd1 vssd1 vccd1 vccd1 _19058_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18707_ _19389_/CLK _18707_/D vssd1 vssd1 vccd1 vccd1 _18707_/Q sky130_fd_sc_hd__dfxtp_1
X_15919_ _15919_/A vssd1 vssd1 vccd1 vccd1 _19294_/D sky130_fd_sc_hd__clkbuf_1
X_19687_ _19687_/CLK _19687_/D vssd1 vssd1 vccd1 vccd1 _19687_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16899_ _16899_/A vssd1 vssd1 vccd1 vccd1 _16904_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_09440_ _10824_/S vssd1 vssd1 vccd1 vccd1 _10670_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18638_ _19292_/CLK _18638_/D vssd1 vssd1 vccd1 vccd1 _18638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09371_ _11001_/A vssd1 vssd1 vccd1 vccd1 _10949_/A sky130_fd_sc_hd__buf_2
X_18569_ _18569_/CLK _18569_/D vssd1 vssd1 vccd1 vccd1 _18569_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_67_clock _19161_/CLK vssd1 vssd1 vccd1 vccd1 _19610_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15303__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12261__A2 _12473_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_165_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_119_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12228__A _19414_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_159_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_165_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_119_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_174_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10024__A1 _10590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13758__S _13758_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_174_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_119_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10971__A _10971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__A1 _19333_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09537__A _10631_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_161_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15973__S _15981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_160_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_141_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_102_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09272__A _16622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ _09707_/A vssd1 vssd1 vccd1 vccd1 _09708_/A sky130_fd_sc_hd__buf_2
XFILLER_114_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_167_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11307__A _11307_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _10704_/S vssd1 vssd1 vccd1 vccd1 _10572_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13514__A_N _14860_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09569_ _18645_/Q vssd1 vssd1 vccd1 vccd1 _10929_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15213__S _15217_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11600_ _09207_/X _11598_/X _11599_/X vssd1 vssd1 vccd1 vccd1 _11600_/Y sky130_fd_sc_hd__o21ai_4
XANTENNA__13522__A _15006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_90_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12580_ _19626_/Q _16931_/A _12526_/X _19156_/Q _12579_/X vssd1 vssd1 vccd1 vccd1
+ _12580_/X sky130_fd_sc_hd__a221o_1
XFILLER_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_142_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_130_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_157_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_129_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15726__A0 _13535_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _11531_/A _11577_/B _17166_/C _09168_/X vssd1 vssd1 vccd1 vccd1 _11532_/D
+ sky130_fd_sc_hd__or4b_1
XFILLER_169_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_168_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_157_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16833__A _16833_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14250_ _14250_/A vssd1 vssd1 vccd1 vccd1 _18631_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_156_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11462_ _11462_/A _11462_/B vssd1 vssd1 vccd1 vccd1 _11462_/Y sky130_fd_sc_hd__nand2_1
XFILLER_165_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13201_ _19445_/Q _13005_/X _13200_/X vssd1 vssd1 vccd1 vccd1 _13201_/X sky130_fd_sc_hd__o21a_1
XFILLER_99_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10413_ _18498_/Q _18993_/Q _10413_/S vssd1 vssd1 vccd1 vccd1 _10414_/B sky130_fd_sc_hd__mux2_1
X_14181_ _14181_/A vssd1 vssd1 vccd1 vccd1 _18601_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ _11404_/A _11393_/B vssd1 vssd1 vccd1 vccd1 _11393_/Y sky130_fd_sc_hd__nor2_1
XFILLER_165_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_124_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_152_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13132_ _13132_/A _13132_/B _13132_/C _12571_/Y vssd1 vssd1 vccd1 vccd1 _13132_/X
+ sky130_fd_sc_hd__or4b_2
XFILLER_99_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_151_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10344_ _18931_/Q _18697_/Q _19379_/Q _19027_/Q _10215_/S _10272_/A vssd1 vssd1 vccd1
+ vccd1 _10345_/B sky130_fd_sc_hd__mux4_1
XANTENNA_input62_A io_ibus_inst[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16151__B1 _15482_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_124_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15883__S _15887_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17940_ _16021_/B _19777_/Q _17946_/S vssd1 vssd1 vccd1 vccd1 _17941_/A sky130_fd_sc_hd__mux2_1
X_13063_ _16055_/B _13064_/C _19752_/Q vssd1 vssd1 vccd1 vccd1 _13065_/B sky130_fd_sc_hd__a21oi_1
XFILLER_79_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10275_ _10482_/A vssd1 vssd1 vccd1 vccd1 _10275_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__09166__B _09166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_140_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12014_ _12009_/Y _12012_/X _12013_/Y vssd1 vssd1 vccd1 vccd1 _12014_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_151_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_105_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_120_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_17871_ _17871_/A _17871_/B vssd1 vssd1 vccd1 vccd1 _17871_/X sky130_fd_sc_hd__or2_1
XFILLER_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output149_A _12080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19610_ _19610_/CLK _19610_/D vssd1 vssd1 vccd1 vccd1 _19610_/Q sky130_fd_sc_hd__dfxtp_1
X_16822_ _16838_/A _16822_/B _16824_/B vssd1 vssd1 vccd1 vccd1 _19580_/D sky130_fd_sc_hd__nor3_1
XANTENNA__17651__B1 _17650_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_120_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_93_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19541_ _19541_/CLK _19541_/D vssd1 vssd1 vccd1 vccd1 _19541_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09567__S0 _10518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_93_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16753_ _19555_/Q _19554_/Q _16753_/C vssd1 vssd1 vccd1 vccd1 _16754_/D sky130_fd_sc_hd__and3_1
XANTENNA__13416__B _18253_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13965_ _14537_/A vssd1 vssd1 vccd1 vccd1 _13965_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_62_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15704_ _14614_/X _19199_/Q _15704_/S vssd1 vssd1 vccd1 vccd1 _15705_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12916_ _16752_/B _12701_/X _12915_/X _12707_/X vssd1 vssd1 vccd1 vccd1 _12916_/X
+ sky130_fd_sc_hd__a211o_1
X_19472_ _19610_/CLK _19472_/D vssd1 vssd1 vccd1 vccd1 _19472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16684_ _16689_/C _16689_/D _16675_/X vssd1 vssd1 vccd1 vccd1 _16684_/Y sky130_fd_sc_hd__a21oi_1
X_13896_ _14576_/A vssd1 vssd1 vccd1 vccd1 _13896_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_73_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18423_ _19306_/CLK _18423_/D vssd1 vssd1 vccd1 vccd1 _18423_/Q sky130_fd_sc_hd__dfxtp_1
X_15635_ _19738_/Q _16024_/S _13430_/B vssd1 vssd1 vccd1 vccd1 _15635_/X sky130_fd_sc_hd__a21o_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _19741_/Q vssd1 vssd1 vccd1 vccd1 _15998_/A sky130_fd_sc_hd__buf_2
XFILLER_34_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18354_ _19235_/CLK _18354_/D vssd1 vssd1 vccd1 vccd1 _18354_/Q sky130_fd_sc_hd__dfxtp_1
X_15566_ _18270_/Q _15566_/B vssd1 vssd1 vccd1 vccd1 _15566_/X sky130_fd_sc_hd__or2_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ _19704_/Q vssd1 vssd1 vccd1 vccd1 _12975_/A sky130_fd_sc_hd__inv_2
XFILLER_148_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17305_ _17305_/A _17305_/B vssd1 vssd1 vccd1 vccd1 _17396_/B sky130_fd_sc_hd__nor2_2
XANTENNA__15717__A0 _13522_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14517_ _18163_/A vssd1 vssd1 vccd1 vccd1 _16833_/A sky130_fd_sc_hd__buf_4
XFILLER_159_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ _11729_/A _11729_/B vssd1 vssd1 vccd1 vccd1 _11788_/A sky130_fd_sc_hd__and2_2
X_18285_ _19300_/CLK _18285_/D vssd1 vssd1 vccd1 vccd1 _18285_/Q sky130_fd_sc_hd__dfxtp_1
X_15497_ _15496_/X _19144_/Q _15517_/S vssd1 vssd1 vccd1 vccd1 _15498_/A sky130_fd_sc_hd__mux2_1
X_17236_ _17231_/X _17234_/Y _17367_/S vssd1 vssd1 vccd1 vccd1 _17236_/X sky130_fd_sc_hd__mux2_1
X_14448_ _13837_/X _18710_/Q _14456_/S vssd1 vssd1 vccd1 vccd1 _14449_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_156_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_155_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10791__A _11331_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17167_ _17121_/A _17121_/B _11574_/B _17124_/B _11508_/A vssd1 vssd1 vccd1 vccd1
+ _17167_/X sky130_fd_sc_hd__o221a_1
XFILLER_156_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14379_ _14379_/A vssd1 vssd1 vccd1 vccd1 _18679_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_155_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_127_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11754__A1 _19396_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16118_ _16114_/X _15588_/X _16117_/Y vssd1 vssd1 vccd1 vccd1 _16118_/X sky130_fd_sc_hd__a21o_1
XFILLER_142_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_143_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17098_ _19695_/Q hold5/A _17098_/S vssd1 vssd1 vccd1 vccd1 _17099_/A sky130_fd_sc_hd__mux2_1
XFILLER_103_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15793__S _15793_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_131_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16049_ _16048_/X _19338_/Q _16053_/S vssd1 vssd1 vccd1 vccd1 _16050_/A sky130_fd_sc_hd__mux2_1
XFILLER_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_111_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19808_ _19845_/CLK _19808_/D vssd1 vssd1 vccd1 vccd1 _19808_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__10730__S _11297_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__A0 _13854_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_96_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09558__S0 _10518_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19739_ _19780_/CLK _19739_/D vssd1 vssd1 vccd1 vccd1 _19739_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__18198__B2 _12482_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10031__A _10031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_65_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_92_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09423_ _11048_/A vssd1 vssd1 vccd1 vccd1 _10951_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__09820__A _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_80_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15541__B hold13/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15033__S _15045_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ input70/X vssd1 vssd1 vccd1 vccd1 _17102_/A sky130_fd_sc_hd__inv_2
XFILLER_40_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_139_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10245__A1 _09844_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15968__S _15970_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _09261_/Y _09271_/X _09280_/X _09284_/X vssd1 vssd1 vccd1 vccd1 _09285_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_21_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16653__A _16666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10796__A2 _10782_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_166_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16920__A2 _12230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_147_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13488__S _13492_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_147_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15269__A _15315_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_134_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_133_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_109_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_133_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_162_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_134_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_121_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10060_ _10060_/A vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__buf_2
XFILLER_125_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_102_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_130_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14112__S _14118_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16828__A _18136_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_141_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18189__B2 _19846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13951__S _13963_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_10962_ _18487_/Q _18982_/Q _10962_/S vssd1 vssd1 vccd1 vccd1 _10963_/A sky130_fd_sc_hd__mux2_1
XFILLER_84_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13750_ _13274_/X _18442_/Q _13758_/S vssd1 vssd1 vccd1 vccd1 _13751_/A sky130_fd_sc_hd__mux2_1
X_12701_ _13055_/A vssd1 vssd1 vccd1 vccd1 _12701_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_10893_ _10889_/A _10890_/X _10892_/X _10883_/X vssd1 vssd1 vccd1 vccd1 _10893_/X
+ sky130_fd_sc_hd__o211a_1
X_13681_ _13681_/A vssd1 vssd1 vccd1 vccd1 _18411_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15420_ _19117_/Q _15041_/X _15422_/S vssd1 vssd1 vccd1 vccd1 _15421_/A sky130_fd_sc_hd__mux2_1
XFILLER_71_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12632_ _13418_/A _12716_/S _14518_/B _18234_/A vssd1 vssd1 vccd1 vccd1 _16921_/S
+ sky130_fd_sc_hd__a31oi_4
XFILLER_70_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12563_ _19605_/Q _12560_/X _12562_/X _19473_/Q vssd1 vssd1 vccd1 vccd1 _13132_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15351_ _15351_/A vssd1 vssd1 vccd1 vccd1 _19086_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14302_ _13837_/X _18646_/Q _14310_/S vssd1 vssd1 vccd1 vccd1 _14303_/A sky130_fd_sc_hd__mux2_1
X_11514_ _17145_/A _17145_/B _17112_/A _17145_/D _17183_/B vssd1 vssd1 vccd1 vccd1
+ _11514_/X sky130_fd_sc_hd__a41o_1
X_18070_ _18070_/A vssd1 vssd1 vccd1 vccd1 _19803_/D sky130_fd_sc_hd__clkbuf_1
X_12494_ _12494_/A _12522_/A _12605_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _12519_/B
+ sky130_fd_sc_hd__or4b_2
X_15282_ _15282_/A vssd1 vssd1 vccd1 vccd1 _19055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16282__B _16282_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17021_ _18097_/A vssd1 vssd1 vccd1 vccd1 _17021_/X sky130_fd_sc_hd__buf_2
XFILLER_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14233_ _14255_/A vssd1 vssd1 vccd1 vccd1 _14242_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_109_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11445_ _11445_/A _12465_/B vssd1 vssd1 vccd1 vccd1 _11446_/B sky130_fd_sc_hd__nand2_1
XFILLER_171_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_125_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_165_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_125_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_171_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_124_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_14164_ _14164_/A vssd1 vssd1 vccd1 vccd1 _18593_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_153_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ _10138_/A _11375_/X _09732_/A vssd1 vssd1 vccd1 vccd1 _11376_/X sky130_fd_sc_hd__a21o_1
XFILLER_166_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_124_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10944__C1 _10943_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_140_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_113_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10327_ _09866_/A _10324_/X _10326_/X _09857_/A vssd1 vssd1 vccd1 vccd1 _10327_/X
+ sky130_fd_sc_hd__o211a_1
X_13115_ _13306_/A _19723_/Q vssd1 vssd1 vccd1 vccd1 _13115_/X sky130_fd_sc_hd__or2_1
X_14095_ _14095_/A vssd1 vssd1 vccd1 vccd1 _18563_/D sky130_fd_sc_hd__clkbuf_1
X_18972_ _19388_/CLK _18972_/D vssd1 vssd1 vccd1 vccd1 _18972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_106_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__A _09905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17571_/A _17309_/Y _17477_/X _17922_/X vssd1 vssd1 vccd1 vccd1 _17923_/X
+ sky130_fd_sc_hd__o211a_1
X_13046_ _11538_/X _13044_/X _13045_/X vssd1 vssd1 vccd1 vccd1 _15038_/A sky130_fd_sc_hd__o21a_4
X_10258_ _09667_/A _10245_/X _10257_/X _09758_/A _19727_/Q vssd1 vssd1 vccd1 vccd1
+ _10303_/A sky130_fd_sc_hd__a32o_4
XFILLER_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_121_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17854_ _17856_/A _17856_/B vssd1 vssd1 vccd1 vccd1 _17854_/Y sky130_fd_sc_hd__nand2_1
X_10189_ _18598_/Q _18869_/Q _19093_/Q _18837_/Q _09854_/X _09871_/A vssd1 vssd1 vccd1
+ vccd1 _10189_/X sky130_fd_sc_hd__mux4_1
XFILLER_121_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10172__B1 _09823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16805_ _19575_/Q _16802_/B _16804_/Y vssd1 vssd1 vccd1 vccd1 _19575_/D sky130_fd_sc_hd__o21a_1
X_17785_ _10398_/Y _17652_/X _17784_/X vssd1 vssd1 vccd1 vccd1 _19725_/D sky130_fd_sc_hd__a21oi_1
XFILLER_82_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09343__C _19843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14997_ _15101_/A vssd1 vssd1 vccd1 vccd1 _14998_/B sky130_fd_sc_hd__clkinv_2
XFILLER_82_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16738__A _16752_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_75_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_94_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19524_ _19524_/CLK _19524_/D vssd1 vssd1 vccd1 vccd1 _19524_/Q sky130_fd_sc_hd__dfxtp_1
X_16736_ _19555_/Q _16736_/B _16736_/C vssd1 vssd1 vccd1 vccd1 _16741_/C sky130_fd_sc_hd__and3_1
XFILLER_93_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13948_ _15317_/A _15854_/B vssd1 vssd1 vccd1 vccd1 _14030_/A sky130_fd_sc_hd__nor2_2
XFILLER_19_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_93_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09640__A _10073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11672__A0 _11618_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19455_ _19524_/CLK _19455_/D vssd1 vssd1 vccd1 vccd1 _19455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16667_ _19531_/Q _16672_/D _16666_/Y vssd1 vssd1 vccd1 vccd1 _19531_/D sky130_fd_sc_hd__o21a_1
XFILLER_34_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13879_ _13879_/A vssd1 vssd1 vccd1 vccd1 _18492_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__10786__A _11321_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18406_ _19287_/CLK _18406_/D vssd1 vssd1 vccd1 vccd1 _18406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15618_ _15618_/A vssd1 vssd1 vccd1 vccd1 _19165_/D sky130_fd_sc_hd__clkbuf_1
X_19386_ _19386_/CLK _19386_/D vssd1 vssd1 vccd1 vccd1 _19386_/Q sky130_fd_sc_hd__dfxtp_1
X_16598_ _19513_/Q _16598_/B vssd1 vssd1 vccd1 vccd1 _16604_/C sky130_fd_sc_hd__and2_1
XFILLER_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18337_ _19314_/CLK _18337_/D vssd1 vssd1 vccd1 vccd1 _18337_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14692__S _14698_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15549_ _15549_/A vssd1 vssd1 vccd1 vccd1 _15549_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_148_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11975__A1 _11969_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18268_ _19162_/CLK _18268_/D vssd1 vssd1 vccd1 vccd1 _18268_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_147_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_149_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17219_ _17219_/A vssd1 vssd1 vccd1 vccd1 _17779_/B sky130_fd_sc_hd__buf_2
XANTENNA__15089__A _15089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18199_ _18231_/A _18199_/B vssd1 vssd1 vccd1 vccd1 _18200_/A sky130_fd_sc_hd__and2_1
XANTENNA__12506__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__A _12422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_144_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_128_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_115_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_115_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_104_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12225__B _12225_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_115_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_171_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_131_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15817__A _15839_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17863__B1 _17862_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_143_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ _19731_/Q vssd1 vssd1 vccd1 vccd1 _09972_/Y sky130_fd_sc_hd__inv_2
XFILLER_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10389__S1 _10263_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14867__S _14871_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15929__A0 _13509_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09406_ _09982_/A vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__buf_2
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13404__B2 hold21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15698__S _15704_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ _18146_/A _18144_/A vssd1 vssd1 vccd1 vccd1 _11522_/C sky130_fd_sc_hd__or2_1
XANTENNA__17146__A2 _17140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_138_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13800__A _13822_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09268_ _19826_/Q _19825_/Q _12522_/A _11803_/A vssd1 vssd1 vccd1 vccd1 _12584_/A
+ sky130_fd_sc_hd__or4b_4
XFILLER_138_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_153_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_153_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14107__S _14107_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_119_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ _19851_/Q vssd1 vssd1 vccd1 vccd1 _18109_/A sky130_fd_sc_hd__clkinv_2
XFILLER_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11230_ _11024_/A _11229_/X _11022_/A vssd1 vssd1 vccd1 vccd1 _11230_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_134_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_134_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _19301_/Q _18713_/Q _18750_/Q _18324_/Q _09496_/A _11030_/X vssd1 vssd1 vccd1
+ vccd1 _11161_/X sky130_fd_sc_hd__mux4_1
XFILLER_150_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10112_ _18504_/Q _18999_/Q _10112_/S vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_150_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11974__B _12134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11092_ _11085_/Y _11087_/Y _11089_/Y _11091_/Y _11044_/A vssd1 vssd1 vccd1 vccd1
+ _11092_/X sky130_fd_sc_hd__o221a_1
XANTENNA__12143__A1 _11351_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14920_ _18906_/Q _14033_/X _14926_/S vssd1 vssd1 vccd1 vccd1 _14921_/A sky130_fd_sc_hd__mux2_1
X_10043_ _19325_/Q _18737_/Q _18774_/Q _18348_/Q _09981_/S _09708_/A vssd1 vssd1 vccd1
+ vccd1 _10043_/X sky130_fd_sc_hd__mux4_1
XFILLER_103_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_103_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_152_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input25_A io_dbus_rdata[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14851_ _14851_/A vssd1 vssd1 vccd1 vccd1 _18875_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__14777__S _14781_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11990__A _12011_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13802_ _13802_/A vssd1 vssd1 vccd1 vccd1 _18464_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ _17831_/A vssd1 vssd1 vccd1 vccd1 _17570_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14782_ _14782_/A vssd1 vssd1 vccd1 vccd1 _18845_/D sky130_fd_sc_hd__clkbuf_1
X_11994_ _19644_/Q _19643_/Q _11994_/C vssd1 vssd1 vccd1 vccd1 _12044_/C sky130_fd_sc_hd__and3_1
XFILLER_16_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16521_ _16541_/A _16521_/B _16521_/C vssd1 vssd1 vccd1 vccd1 _19488_/D sky130_fd_sc_hd__nor3_1
X_13733_ _13733_/A vssd1 vssd1 vccd1 vccd1 _18434_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__09942__S0 _09840_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10945_ _18583_/Q _18854_/Q _19078_/Q _18822_/Q _11049_/S _10937_/A vssd1 vssd1 vccd1
+ vccd1 _10945_/X sky130_fd_sc_hd__mux4_1
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_19240_ _19306_/CLK _19240_/D vssd1 vssd1 vccd1 vccd1 _19240_/Q sky130_fd_sc_hd__dfxtp_1
X_16452_ _16485_/A _16452_/B _16452_/C vssd1 vssd1 vccd1 vccd1 _19467_/D sky130_fd_sc_hd__nor3_1
X_13664_ _13171_/X _18404_/Q _13664_/S vssd1 vssd1 vccd1 vccd1 _13665_/A sky130_fd_sc_hd__mux2_1
X_10876_ _09393_/A _10873_/X _11064_/A vssd1 vssd1 vccd1 vccd1 _10876_/X sky130_fd_sc_hd__a21o_1
X_15403_ _19109_/Q _15015_/X _15411_/S vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__mux2_1
X_12615_ _13400_/A _18254_/Q vssd1 vssd1 vccd1 vccd1 _12615_/Y sky130_fd_sc_hd__nand2_1
X_19171_ _19235_/CLK _19171_/D vssd1 vssd1 vccd1 vccd1 _19171_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11406__B1 _09823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16383_ _19443_/Q _16381_/B _16382_/Y vssd1 vssd1 vccd1 vccd1 _19443_/D sky130_fd_sc_hd__o21a_1
XANTENNA__13946__A2 _16622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16293__A _18079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13595_ _15079_/A vssd1 vssd1 vccd1 vccd1 _13595_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_129_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_169_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_18122_ _18122_/A _18135_/B vssd1 vssd1 vccd1 vccd1 _18122_/X sky130_fd_sc_hd__or2_1
X_15334_ _15334_/A vssd1 vssd1 vccd1 vccd1 _19078_/D sky130_fd_sc_hd__clkbuf_1
X_12546_ _15613_/A vssd1 vssd1 vccd1 vccd1 _12713_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_157_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_leaf_150_clock_A clkbuf_4_10_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18053_ _19796_/Q _19417_/Q _18061_/S vssd1 vssd1 vccd1 vccd1 _18054_/A sky130_fd_sc_hd__mux2_1
X_15265_ _14547_/X _19048_/Q _15267_/S vssd1 vssd1 vccd1 vccd1 _15266_/A sky130_fd_sc_hd__mux2_1
XFILLER_126_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12477_ _12480_/A _12477_/B vssd1 vssd1 vccd1 vccd1 _12477_/Y sky130_fd_sc_hd__nor2_1
XFILLER_126_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17004_ _12689_/X _16997_/X _17003_/X _16995_/X vssd1 vssd1 vccd1 vccd1 _19654_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_output93_A _11644_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ _18616_/Q _13972_/X _14220_/S vssd1 vssd1 vccd1 vccd1 _14217_/A sky130_fd_sc_hd__mux2_1
XANTENNA__10068__S0 _10017_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11428_ _11428_/A _11428_/B vssd1 vssd1 vccd1 vccd1 _11428_/X sky130_fd_sc_hd__and2_1
XFILLER_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ _15196_/A vssd1 vssd1 vccd1 vccd1 _19017_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_125_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10917__C1 _09553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12382__A1 _11418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_152_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_113_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14147_ _18586_/Q _13978_/X _14147_/S vssd1 vssd1 vccd1 vccd1 _14148_/A sky130_fd_sc_hd__mux2_1
X_11359_ _11435_/A _11437_/A _11435_/C _10182_/A _11358_/Y vssd1 vssd1 vccd1 vccd1
+ _11431_/C sky130_fd_sc_hd__a311o_1
XANTENNA__14659__A0 _14541_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_112_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15320__A1 _14996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ _14078_/A vssd1 vssd1 vccd1 vccd1 _18555_/D sky130_fd_sc_hd__clkbuf_1
X_18955_ _18987_/CLK _18955_/D vssd1 vssd1 vccd1 vccd1 _18955_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17906_ _17907_/B _17906_/B vssd1 vssd1 vccd1 vccd1 _17910_/B sky130_fd_sc_hd__nand2_1
X_13029_ _19750_/Q vssd1 vssd1 vccd1 vccd1 _16055_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18886_ _19367_/CLK _18886_/D vssd1 vssd1 vccd1 vccd1 _18886_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12685__A2 _12507_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11488__A3 _11492_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_94_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17837_ _17626_/X _17834_/X _17836_/Y _17532_/A vssd1 vssd1 vccd1 vccd1 _17837_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14687__S _14687_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16281__C1 _16280_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17768_ _17215_/X _17768_/B vssd1 vssd1 vccd1 vccd1 _17768_/X sky130_fd_sc_hd__and2b_1
XFILLER_81_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_75_clock_A clkbuf_4_6_0_clock/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__A2 _12433_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_82_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16719_ _16724_/C _16724_/D _16718_/X vssd1 vssd1 vccd1 vccd1 _16719_/Y sky130_fd_sc_hd__a21oi_1
X_19507_ _19540_/CLK _19507_/D vssd1 vssd1 vccd1 vccd1 _19507_/Q sky130_fd_sc_hd__dfxtp_1
X_17699_ _17478_/X _17692_/Y _17698_/X _17422_/A vssd1 vssd1 vccd1 vccd1 _17699_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_23_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10543__S1 _09590_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19438_ _19583_/CLK _19438_/D vssd1 vssd1 vccd1 vccd1 _19438_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_148_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19369_ _19369_/CLK _19369_/D vssd1 vssd1 vccd1 vccd1 _19369_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__14716__A _14772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15311__S _15311_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09122_ _09166_/A vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_148_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10620__B2 _19719_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11140__A _11254_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_151_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_117_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_144_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_116_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_104_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_117_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_116_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_143_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ _18633_/Q _18968_/Q _09955_/S vssd1 vssd1 vccd1 vccd1 _09956_/B sky130_fd_sc_hd__mux2_1
XFILLER_104_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13322__B1 _13321_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15981__S _15981_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_103_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_131_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_106_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_09886_ _09886_/A vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__buf_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17064__A1 _15550_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10687__A1 _09820_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_85_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13514__B _18091_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10730_ _18491_/Q _18986_/Q _11297_/S vssd1 vssd1 vccd1 vccd1 _10730_/X sky130_fd_sc_hd__mux2_1
X_10661_ _18460_/Q _19051_/Q _19213_/Q _18428_/Q _10660_/X _09707_/A vssd1 vssd1 vccd1
+ vccd1 _10661_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12400_ _17305_/A vssd1 vssd1 vccd1 vccd1 _17387_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_51_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13380_ _16520_/B _13260_/X _13261_/X _16321_/B _13379_/X vssd1 vssd1 vccd1 vccd1
+ _13380_/X sky130_fd_sc_hd__a221o_4
XFILLER_139_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_167_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__11969__B _11969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10592_ _10585_/A _10591_/X _10074_/X vssd1 vssd1 vccd1 vccd1 _10592_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_166_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_167_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_12331_ _17312_/A _17867_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12332_/B sky130_fd_sc_hd__a21oi_2
XFILLER_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_108_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15050_ _15050_/A vssd1 vssd1 vccd1 vccd1 _18959_/D sky130_fd_sc_hd__clkbuf_1
X_12262_ _12242_/B _12240_/A _17305_/A vssd1 vssd1 vccd1 vccd1 _12263_/B sky130_fd_sc_hd__a21o_1
XFILLER_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_135_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14001_ _14573_/A vssd1 vssd1 vccd1 vccd1 _14001_/X sky130_fd_sc_hd__clkbuf_2
X_11213_ _11007_/X _11206_/X _11208_/X _11212_/X _09464_/A vssd1 vssd1 vccd1 vccd1
+ _11213_/X sky130_fd_sc_hd__a311o_1
XFILLER_122_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12193_ _19792_/Q _11354_/A _12404_/S vssd1 vssd1 vccd1 vccd1 _12195_/A sky130_fd_sc_hd__mux2_4
X_11144_ _10807_/A _11141_/X _11143_/X _11134_/X vssd1 vssd1 vccd1 vccd1 _11144_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_123_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10470__S0 _10260_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput74 _11968_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[12] sky130_fd_sc_hd__buf_2
XFILLER_68_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput85 _12225_/B vssd1 vssd1 vccd1 vccd1 io_dbus_addr[22] sky130_fd_sc_hd__buf_2
XFILLER_163_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput96 _11683_/X vssd1 vssd1 vccd1 vccd1 io_dbus_addr[3] sky130_fd_sc_hd__buf_2
XANTENNA__11196__S _11196_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18740_ _19296_/CLK _18740_/D vssd1 vssd1 vccd1 vccd1 _18740_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_89_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15952_ _15952_/A vssd1 vssd1 vccd1 vccd1 _19308_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11075_ _11075_/A _11074_/X vssd1 vssd1 vccd1 vccd1 _11075_/X sky130_fd_sc_hd__or2b_1
XANTENNA__10127__B1 _09823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17055__A1 _12651_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14903_ _14903_/A vssd1 vssd1 vccd1 vccd1 _18898_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10026_ _09485_/A _10014_/Y _10020_/X _10025_/Y _09811_/A vssd1 vssd1 vccd1 vccd1
+ _10026_/X sky130_fd_sc_hd__o311a_4
XFILLER_102_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18671_ _19385_/CLK _18671_/D vssd1 vssd1 vccd1 vccd1 _18671_/Q sky130_fd_sc_hd__dfxtp_1
X_15883_ _19278_/Q _14560_/A _15887_/S vssd1 vssd1 vccd1 vccd1 _15884_/A sky130_fd_sc_hd__mux2_1
XFILLER_76_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17622_ _17622_/A vssd1 vssd1 vccd1 vccd1 _17622_/Y sky130_fd_sc_hd__clkinv_2
X_14834_ _14845_/A vssd1 vssd1 vccd1 vccd1 _14843_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__13705__A _13762_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11627__B1 _11600_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17553_ _17576_/S _17369_/X _17552_/Y _17550_/S vssd1 vssd1 vccd1 vccd1 _17553_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09296__A1 _19627_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14765_ _14765_/A vssd1 vssd1 vccd1 vccd1 _18837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09296__B2 _19628_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11977_ _12020_/A _12460_/A _11976_/Y vssd1 vssd1 vccd1 vccd1 _12025_/C sky130_fd_sc_hd__a21oi_1
XFILLER_17_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_16504_ _16524_/A _16504_/B vssd1 vssd1 vccd1 vccd1 _16504_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ _13762_/S vssd1 vssd1 vccd1 vccd1 _13725_/S sky130_fd_sc_hd__clkbuf_4
X_17484_ _17479_/X _17700_/A _17483_/X vssd1 vssd1 vccd1 vccd1 _17484_/Y sky130_fd_sc_hd__a21oi_2
X_10928_ _10961_/A _10927_/X _10915_/X vssd1 vssd1 vccd1 vccd1 _10928_/Y sky130_fd_sc_hd__o21ai_1
X_14696_ _14595_/X _18807_/Q _14698_/S vssd1 vssd1 vccd1 vccd1 _14697_/A sky130_fd_sc_hd__mux2_1
XFILLER_44_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19223_ _19223_/CLK _19223_/D vssd1 vssd1 vccd1 vccd1 _19223_/Q sky130_fd_sc_hd__dfxtp_1
X_16435_ _16435_/A vssd1 vssd1 vccd1 vccd1 _16440_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ _13038_/X _18396_/Q _13653_/S vssd1 vssd1 vccd1 vccd1 _13648_/A sky130_fd_sc_hd__mux2_1
XFILLER_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10859_ _10855_/A _10853_/Y _10855_/Y _10977_/A vssd1 vssd1 vccd1 vccd1 _10859_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_72_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16227__S _16235_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_158_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19154_ _19688_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 _19154_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16366_ _16390_/A _16371_/C vssd1 vssd1 vccd1 vccd1 _16366_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11879__B _19401_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ _13578_/A vssd1 vssd1 vccd1 vccd1 _18372_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_158_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_158_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18105_ _19817_/Q _18086_/X _18104_/Y _18097_/X vssd1 vssd1 vccd1 vccd1 _19817_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_173_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_158_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15317_ _15317_/A _15317_/B vssd1 vssd1 vccd1 vccd1 _15374_/A sky130_fd_sc_hd__nor2_2
X_12529_ _12529_/A vssd1 vssd1 vccd1 vccd1 _12601_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_19085_ _19085_/CLK _19085_/D vssd1 vssd1 vccd1 vccd1 _19085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_117_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16297_ _19416_/Q _16278_/X _12278_/X _16269_/X vssd1 vssd1 vccd1 vccd1 _19416_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_117_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_172_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_145_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18036_ _19789_/Q _12126_/A _18038_/S vssd1 vssd1 vccd1 vccd1 _18037_/A sky130_fd_sc_hd__mux2_1
X_15248_ _14519_/X _19040_/Q _15256_/S vssd1 vssd1 vccd1 vccd1 _15249_/A sky130_fd_sc_hd__mux2_1
XFILLER_173_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_172_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_132_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17818__B1 _17817_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_153_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14271__A _18172_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_126_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_15179_ _15179_/A vssd1 vssd1 vccd1 vccd1 _19009_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_141_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_98_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_114_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_99_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12107__A1 _19409_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_87_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_141_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09740_ _09740_/A vssd1 vssd1 vccd1 vccd1 _09740_/X sky130_fd_sc_hd__buf_2
XANTENNA__10118__B1 _09823_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18938_ _19386_/CLK _18938_/D vssd1 vssd1 vccd1 vccd1 _18938_/Q sky130_fd_sc_hd__dfxtp_1
.ends

