VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO WBM_DBus
  CLASS BLOCK ;
  FOREIGN WBM_DBus ;
  ORIGIN 0.000 0.000 ;
  SIZE 180.000 BY 180.000 ;
  PIN io_dbus_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_dbus_addr[0]
  PIN io_dbus_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_dbus_addr[10]
  PIN io_dbus_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 176.000 58.330 180.000 ;
    END
  END io_dbus_addr[11]
  PIN io_dbus_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 23.840 180.000 24.440 ;
    END
  END io_dbus_addr[12]
  PIN io_dbus_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_dbus_addr[13]
  PIN io_dbus_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 176.000 77.650 180.000 ;
    END
  END io_dbus_addr[14]
  PIN io_dbus_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_dbus_addr[15]
  PIN io_dbus_addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 51.040 180.000 51.640 ;
    END
  END io_dbus_addr[16]
  PIN io_dbus_addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END io_dbus_addr[17]
  PIN io_dbus_addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END io_dbus_addr[18]
  PIN io_dbus_addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_dbus_addr[19]
  PIN io_dbus_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 132.640 180.000 133.240 ;
    END
  END io_dbus_addr[1]
  PIN io_dbus_addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END io_dbus_addr[20]
  PIN io_dbus_addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_dbus_addr[21]
  PIN io_dbus_addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_dbus_addr[22]
  PIN io_dbus_addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 17.040 180.000 17.640 ;
    END
  END io_dbus_addr[23]
  PIN io_dbus_addr[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 176.000 64.770 180.000 ;
    END
  END io_dbus_addr[24]
  PIN io_dbus_addr[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END io_dbus_addr[25]
  PIN io_dbus_addr[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END io_dbus_addr[26]
  PIN io_dbus_addr[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 176.000 16.470 180.000 ;
    END
  END io_dbus_addr[27]
  PIN io_dbus_addr[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 176.000 109.850 180.000 ;
    END
  END io_dbus_addr[28]
  PIN io_dbus_addr[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END io_dbus_addr[29]
  PIN io_dbus_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END io_dbus_addr[2]
  PIN io_dbus_addr[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END io_dbus_addr[30]
  PIN io_dbus_addr[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 176.000 100.190 180.000 ;
    END
  END io_dbus_addr[31]
  PIN io_dbus_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 129.240 180.000 129.840 ;
    END
  END io_dbus_addr[3]
  PIN io_dbus_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_dbus_addr[4]
  PIN io_dbus_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_dbus_addr[5]
  PIN io_dbus_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 156.440 180.000 157.040 ;
    END
  END io_dbus_addr[6]
  PIN io_dbus_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END io_dbus_addr[7]
  PIN io_dbus_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 176.000 51.890 180.000 ;
    END
  END io_dbus_addr[8]
  PIN io_dbus_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 176.000 151.710 180.000 ;
    END
  END io_dbus_addr[9]
  PIN io_dbus_ld_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 119.040 180.000 119.640 ;
    END
  END io_dbus_ld_type[0]
  PIN io_dbus_ld_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 173.440 180.000 174.040 ;
    END
  END io_dbus_ld_type[1]
  PIN io_dbus_ld_type[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 176.000 13.250 180.000 ;
    END
  END io_dbus_ld_type[2]
  PIN io_dbus_rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 91.840 180.000 92.440 ;
    END
  END io_dbus_rd_en
  PIN io_dbus_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 159.840 180.000 160.440 ;
    END
  END io_dbus_rdata[0]
  PIN io_dbus_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 57.840 180.000 58.440 ;
    END
  END io_dbus_rdata[10]
  PIN io_dbus_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END io_dbus_rdata[11]
  PIN io_dbus_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END io_dbus_rdata[12]
  PIN io_dbus_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 176.000 90.530 180.000 ;
    END
  END io_dbus_rdata[13]
  PIN io_dbus_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END io_dbus_rdata[14]
  PIN io_dbus_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_dbus_rdata[15]
  PIN io_dbus_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_dbus_rdata[16]
  PIN io_dbus_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END io_dbus_rdata[17]
  PIN io_dbus_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 176.000 93.750 180.000 ;
    END
  END io_dbus_rdata[18]
  PIN io_dbus_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 170.040 180.000 170.640 ;
    END
  END io_dbus_rdata[19]
  PIN io_dbus_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_dbus_rdata[1]
  PIN io_dbus_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 176.000 161.370 180.000 ;
    END
  END io_dbus_rdata[20]
  PIN io_dbus_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 176.000 148.490 180.000 ;
    END
  END io_dbus_rdata[21]
  PIN io_dbus_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 176.000 135.610 180.000 ;
    END
  END io_dbus_rdata[22]
  PIN io_dbus_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_dbus_rdata[23]
  PIN io_dbus_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 74.840 180.000 75.440 ;
    END
  END io_dbus_rdata[24]
  PIN io_dbus_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_dbus_rdata[25]
  PIN io_dbus_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END io_dbus_rdata[26]
  PIN io_dbus_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END io_dbus_rdata[27]
  PIN io_dbus_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_dbus_rdata[28]
  PIN io_dbus_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 176.000 32.570 180.000 ;
    END
  END io_dbus_rdata[29]
  PIN io_dbus_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 176.000 67.990 180.000 ;
    END
  END io_dbus_rdata[2]
  PIN io_dbus_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END io_dbus_rdata[30]
  PIN io_dbus_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 139.440 180.000 140.040 ;
    END
  END io_dbus_rdata[31]
  PIN io_dbus_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END io_dbus_rdata[3]
  PIN io_dbus_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END io_dbus_rdata[4]
  PIN io_dbus_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 44.240 180.000 44.840 ;
    END
  END io_dbus_rdata[5]
  PIN io_dbus_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 88.440 180.000 89.040 ;
    END
  END io_dbus_rdata[6]
  PIN io_dbus_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END io_dbus_rdata[7]
  PIN io_dbus_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 20.440 180.000 21.040 ;
    END
  END io_dbus_rdata[8]
  PIN io_dbus_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_dbus_rdata[9]
  PIN io_dbus_st_type[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 176.000 158.150 180.000 ;
    END
  END io_dbus_st_type[0]
  PIN io_dbus_st_type[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 176.000 26.130 180.000 ;
    END
  END io_dbus_st_type[1]
  PIN io_dbus_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 176.000 48.670 180.000 ;
    END
  END io_dbus_valid
  PIN io_dbus_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 40.840 180.000 41.440 ;
    END
  END io_dbus_wdata[0]
  PIN io_dbus_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END io_dbus_wdata[10]
  PIN io_dbus_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END io_dbus_wdata[11]
  PIN io_dbus_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 176.000 142.050 180.000 ;
    END
  END io_dbus_wdata[12]
  PIN io_dbus_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 146.240 180.000 146.840 ;
    END
  END io_dbus_wdata[13]
  PIN io_dbus_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END io_dbus_wdata[14]
  PIN io_dbus_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_dbus_wdata[15]
  PIN io_dbus_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 176.000 45.450 180.000 ;
    END
  END io_dbus_wdata[16]
  PIN io_dbus_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 176.000 154.930 180.000 ;
    END
  END io_dbus_wdata[17]
  PIN io_dbus_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 95.240 180.000 95.840 ;
    END
  END io_dbus_wdata[18]
  PIN io_dbus_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_dbus_wdata[19]
  PIN io_dbus_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 176.000 119.510 180.000 ;
    END
  END io_dbus_wdata[1]
  PIN io_dbus_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 105.440 180.000 106.040 ;
    END
  END io_dbus_wdata[20]
  PIN io_dbus_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_dbus_wdata[21]
  PIN io_dbus_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 176.000 3.590 180.000 ;
    END
  END io_dbus_wdata[22]
  PIN io_dbus_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END io_dbus_wdata[23]
  PIN io_dbus_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END io_dbus_wdata[24]
  PIN io_dbus_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_dbus_wdata[25]
  PIN io_dbus_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 176.000 167.810 180.000 ;
    END
  END io_dbus_wdata[26]
  PIN io_dbus_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 176.000 55.110 180.000 ;
    END
  END io_dbus_wdata[27]
  PIN io_dbus_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END io_dbus_wdata[28]
  PIN io_dbus_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END io_dbus_wdata[29]
  PIN io_dbus_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 176.000 132.390 180.000 ;
    END
  END io_dbus_wdata[2]
  PIN io_dbus_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 6.840 180.000 7.440 ;
    END
  END io_dbus_wdata[30]
  PIN io_dbus_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END io_dbus_wdata[31]
  PIN io_dbus_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 3.440 180.000 4.040 ;
    END
  END io_dbus_wdata[3]
  PIN io_dbus_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_dbus_wdata[4]
  PIN io_dbus_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_dbus_wdata[5]
  PIN io_dbus_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 98.640 180.000 99.240 ;
    END
  END io_dbus_wdata[6]
  PIN io_dbus_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END io_dbus_wdata[7]
  PIN io_dbus_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_dbus_wdata[8]
  PIN io_dbus_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 176.000 106.630 180.000 ;
    END
  END io_dbus_wdata[9]
  PIN io_dbus_wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END io_dbus_wr_en
  PIN io_wbm_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 176.840 180.000 177.440 ;
    END
  END io_wbm_ack_i
  PIN io_wbm_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END io_wbm_data_i[0]
  PIN io_wbm_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_wbm_data_i[10]
  PIN io_wbm_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 153.040 180.000 153.640 ;
    END
  END io_wbm_data_i[11]
  PIN io_wbm_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 176.000 0.370 180.000 ;
    END
  END io_wbm_data_i[12]
  PIN io_wbm_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 68.040 180.000 68.640 ;
    END
  END io_wbm_data_i[13]
  PIN io_wbm_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END io_wbm_data_i[14]
  PIN io_wbm_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 102.040 180.000 102.640 ;
    END
  END io_wbm_data_i[15]
  PIN io_wbm_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END io_wbm_data_i[16]
  PIN io_wbm_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 176.000 22.910 180.000 ;
    END
  END io_wbm_data_i[17]
  PIN io_wbm_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 112.240 180.000 112.840 ;
    END
  END io_wbm_data_i[18]
  PIN io_wbm_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END io_wbm_data_i[19]
  PIN io_wbm_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END io_wbm_data_i[1]
  PIN io_wbm_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 176.000 71.210 180.000 ;
    END
  END io_wbm_data_i[20]
  PIN io_wbm_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_wbm_data_i[21]
  PIN io_wbm_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_wbm_data_i[22]
  PIN io_wbm_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 176.000 174.250 180.000 ;
    END
  END io_wbm_data_i[23]
  PIN io_wbm_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 71.440 180.000 72.040 ;
    END
  END io_wbm_data_i[24]
  PIN io_wbm_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 176.000 74.430 180.000 ;
    END
  END io_wbm_data_i[25]
  PIN io_wbm_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 176.000 103.410 180.000 ;
    END
  END io_wbm_data_i[26]
  PIN io_wbm_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 176.000 96.970 180.000 ;
    END
  END io_wbm_data_i[27]
  PIN io_wbm_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END io_wbm_data_i[28]
  PIN io_wbm_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END io_wbm_data_i[29]
  PIN io_wbm_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 30.640 180.000 31.240 ;
    END
  END io_wbm_data_i[2]
  PIN io_wbm_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END io_wbm_data_i[30]
  PIN io_wbm_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 149.640 180.000 150.240 ;
    END
  END io_wbm_data_i[31]
  PIN io_wbm_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 176.000 39.010 180.000 ;
    END
  END io_wbm_data_i[3]
  PIN io_wbm_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 176.000 116.290 180.000 ;
    END
  END io_wbm_data_i[4]
  PIN io_wbm_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_wbm_data_i[5]
  PIN io_wbm_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 47.640 180.000 48.240 ;
    END
  END io_wbm_data_i[6]
  PIN io_wbm_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_wbm_data_i[7]
  PIN io_wbm_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 176.000 42.230 180.000 ;
    END
  END io_wbm_data_i[8]
  PIN io_wbm_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 78.240 180.000 78.840 ;
    END
  END io_wbm_data_i[9]
  PIN io_wbm_m2s_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 10.240 180.000 10.840 ;
    END
  END io_wbm_m2s_addr[0]
  PIN io_wbm_m2s_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_wbm_m2s_addr[10]
  PIN io_wbm_m2s_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 142.840 180.000 143.440 ;
    END
  END io_wbm_m2s_addr[11]
  PIN io_wbm_m2s_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_wbm_m2s_addr[12]
  PIN io_wbm_m2s_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_wbm_m2s_addr[13]
  PIN io_wbm_m2s_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 61.240 180.000 61.840 ;
    END
  END io_wbm_m2s_addr[14]
  PIN io_wbm_m2s_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END io_wbm_m2s_addr[15]
  PIN io_wbm_m2s_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 13.640 180.000 14.240 ;
    END
  END io_wbm_m2s_addr[1]
  PIN io_wbm_m2s_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 176.000 6.810 180.000 ;
    END
  END io_wbm_m2s_addr[2]
  PIN io_wbm_m2s_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END io_wbm_m2s_addr[3]
  PIN io_wbm_m2s_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_wbm_m2s_addr[4]
  PIN io_wbm_m2s_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END io_wbm_m2s_addr[5]
  PIN io_wbm_m2s_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 37.440 180.000 38.040 ;
    END
  END io_wbm_m2s_addr[6]
  PIN io_wbm_m2s_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 166.640 180.000 167.240 ;
    END
  END io_wbm_m2s_addr[7]
  PIN io_wbm_m2s_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 115.640 180.000 116.240 ;
    END
  END io_wbm_m2s_addr[8]
  PIN io_wbm_m2s_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END io_wbm_m2s_addr[9]
  PIN io_wbm_m2s_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_wbm_m2s_data[0]
  PIN io_wbm_m2s_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 64.640 180.000 65.240 ;
    END
  END io_wbm_m2s_data[10]
  PIN io_wbm_m2s_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END io_wbm_m2s_data[11]
  PIN io_wbm_m2s_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 125.840 180.000 126.440 ;
    END
  END io_wbm_m2s_data[12]
  PIN io_wbm_m2s_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 176.000 177.470 180.000 ;
    END
  END io_wbm_m2s_data[13]
  PIN io_wbm_m2s_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_wbm_m2s_data[14]
  PIN io_wbm_m2s_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 176.000 171.030 180.000 ;
    END
  END io_wbm_m2s_data[15]
  PIN io_wbm_m2s_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_wbm_m2s_data[16]
  PIN io_wbm_m2s_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_wbm_m2s_data[17]
  PIN io_wbm_m2s_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END io_wbm_m2s_data[18]
  PIN io_wbm_m2s_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_wbm_m2s_data[19]
  PIN io_wbm_m2s_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END io_wbm_m2s_data[1]
  PIN io_wbm_m2s_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_wbm_m2s_data[20]
  PIN io_wbm_m2s_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 176.000 19.690 180.000 ;
    END
  END io_wbm_m2s_data[21]
  PIN io_wbm_m2s_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 176.000 84.090 180.000 ;
    END
  END io_wbm_m2s_data[22]
  PIN io_wbm_m2s_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_wbm_m2s_data[23]
  PIN io_wbm_m2s_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_wbm_m2s_data[24]
  PIN io_wbm_m2s_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END io_wbm_m2s_data[25]
  PIN io_wbm_m2s_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 176.000 122.730 180.000 ;
    END
  END io_wbm_m2s_data[26]
  PIN io_wbm_m2s_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 176.000 80.870 180.000 ;
    END
  END io_wbm_m2s_data[27]
  PIN io_wbm_m2s_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END io_wbm_m2s_data[28]
  PIN io_wbm_m2s_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 176.000 145.270 180.000 ;
    END
  END io_wbm_m2s_data[29]
  PIN io_wbm_m2s_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 34.040 180.000 34.640 ;
    END
  END io_wbm_m2s_data[2]
  PIN io_wbm_m2s_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_wbm_m2s_data[30]
  PIN io_wbm_m2s_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END io_wbm_m2s_data[31]
  PIN io_wbm_m2s_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END io_wbm_m2s_data[3]
  PIN io_wbm_m2s_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END io_wbm_m2s_data[4]
  PIN io_wbm_m2s_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END io_wbm_m2s_data[5]
  PIN io_wbm_m2s_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 122.440 180.000 123.040 ;
    END
  END io_wbm_m2s_data[6]
  PIN io_wbm_m2s_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END io_wbm_m2s_data[7]
  PIN io_wbm_m2s_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 176.000 129.170 180.000 ;
    END
  END io_wbm_m2s_data[8]
  PIN io_wbm_m2s_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 176.000 125.950 180.000 ;
    END
  END io_wbm_m2s_data[9]
  PIN io_wbm_m2s_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_wbm_m2s_sel[0]
  PIN io_wbm_m2s_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 176.000 29.350 180.000 ;
    END
  END io_wbm_m2s_sel[1]
  PIN io_wbm_m2s_sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END io_wbm_m2s_sel[2]
  PIN io_wbm_m2s_sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END io_wbm_m2s_sel[3]
  PIN io_wbm_m2s_stb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_wbm_m2s_stb
  PIN io_wbm_m2s_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.000 85.040 180.000 85.640 ;
    END
  END io_wbm_m2s_we
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 32.880 10.640 34.480 168.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.200 10.640 90.800 168.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 145.520 10.640 147.120 168.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 61.040 10.640 62.640 168.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 117.360 10.640 118.960 168.880 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 174.340 168.725 ;
      LAYER met1 ;
        RECT 0.070 8.880 177.490 169.960 ;
      LAYER met2 ;
        RECT 0.650 175.720 3.030 177.325 ;
        RECT 3.870 175.720 6.250 177.325 ;
        RECT 7.090 175.720 12.690 177.325 ;
        RECT 13.530 175.720 15.910 177.325 ;
        RECT 16.750 175.720 19.130 177.325 ;
        RECT 19.970 175.720 22.350 177.325 ;
        RECT 23.190 175.720 25.570 177.325 ;
        RECT 26.410 175.720 28.790 177.325 ;
        RECT 29.630 175.720 32.010 177.325 ;
        RECT 32.850 175.720 38.450 177.325 ;
        RECT 39.290 175.720 41.670 177.325 ;
        RECT 42.510 175.720 44.890 177.325 ;
        RECT 45.730 175.720 48.110 177.325 ;
        RECT 48.950 175.720 51.330 177.325 ;
        RECT 52.170 175.720 54.550 177.325 ;
        RECT 55.390 175.720 57.770 177.325 ;
        RECT 58.610 175.720 64.210 177.325 ;
        RECT 65.050 175.720 67.430 177.325 ;
        RECT 68.270 175.720 70.650 177.325 ;
        RECT 71.490 175.720 73.870 177.325 ;
        RECT 74.710 175.720 77.090 177.325 ;
        RECT 77.930 175.720 80.310 177.325 ;
        RECT 81.150 175.720 83.530 177.325 ;
        RECT 84.370 175.720 89.970 177.325 ;
        RECT 90.810 175.720 93.190 177.325 ;
        RECT 94.030 175.720 96.410 177.325 ;
        RECT 97.250 175.720 99.630 177.325 ;
        RECT 100.470 175.720 102.850 177.325 ;
        RECT 103.690 175.720 106.070 177.325 ;
        RECT 106.910 175.720 109.290 177.325 ;
        RECT 110.130 175.720 115.730 177.325 ;
        RECT 116.570 175.720 118.950 177.325 ;
        RECT 119.790 175.720 122.170 177.325 ;
        RECT 123.010 175.720 125.390 177.325 ;
        RECT 126.230 175.720 128.610 177.325 ;
        RECT 129.450 175.720 131.830 177.325 ;
        RECT 132.670 175.720 135.050 177.325 ;
        RECT 135.890 175.720 141.490 177.325 ;
        RECT 142.330 175.720 144.710 177.325 ;
        RECT 145.550 175.720 147.930 177.325 ;
        RECT 148.770 175.720 151.150 177.325 ;
        RECT 151.990 175.720 154.370 177.325 ;
        RECT 155.210 175.720 157.590 177.325 ;
        RECT 158.430 175.720 160.810 177.325 ;
        RECT 161.650 175.720 167.250 177.325 ;
        RECT 168.090 175.720 170.470 177.325 ;
        RECT 171.310 175.720 173.690 177.325 ;
        RECT 174.530 175.720 176.910 177.325 ;
        RECT 0.100 4.280 177.460 175.720 ;
        RECT 0.650 3.555 3.030 4.280 ;
        RECT 3.870 3.555 6.250 4.280 ;
        RECT 7.090 3.555 9.470 4.280 ;
        RECT 10.310 3.555 12.690 4.280 ;
        RECT 13.530 3.555 15.910 4.280 ;
        RECT 16.750 3.555 19.130 4.280 ;
        RECT 19.970 3.555 22.350 4.280 ;
        RECT 23.190 3.555 28.790 4.280 ;
        RECT 29.630 3.555 32.010 4.280 ;
        RECT 32.850 3.555 35.230 4.280 ;
        RECT 36.070 3.555 38.450 4.280 ;
        RECT 39.290 3.555 41.670 4.280 ;
        RECT 42.510 3.555 44.890 4.280 ;
        RECT 45.730 3.555 48.110 4.280 ;
        RECT 48.950 3.555 54.550 4.280 ;
        RECT 55.390 3.555 57.770 4.280 ;
        RECT 58.610 3.555 60.990 4.280 ;
        RECT 61.830 3.555 64.210 4.280 ;
        RECT 65.050 3.555 67.430 4.280 ;
        RECT 68.270 3.555 70.650 4.280 ;
        RECT 71.490 3.555 73.870 4.280 ;
        RECT 74.710 3.555 80.310 4.280 ;
        RECT 81.150 3.555 83.530 4.280 ;
        RECT 84.370 3.555 86.750 4.280 ;
        RECT 87.590 3.555 89.970 4.280 ;
        RECT 90.810 3.555 93.190 4.280 ;
        RECT 94.030 3.555 96.410 4.280 ;
        RECT 97.250 3.555 99.630 4.280 ;
        RECT 100.470 3.555 106.070 4.280 ;
        RECT 106.910 3.555 109.290 4.280 ;
        RECT 110.130 3.555 112.510 4.280 ;
        RECT 113.350 3.555 115.730 4.280 ;
        RECT 116.570 3.555 118.950 4.280 ;
        RECT 119.790 3.555 122.170 4.280 ;
        RECT 123.010 3.555 125.390 4.280 ;
        RECT 126.230 3.555 131.830 4.280 ;
        RECT 132.670 3.555 135.050 4.280 ;
        RECT 135.890 3.555 138.270 4.280 ;
        RECT 139.110 3.555 141.490 4.280 ;
        RECT 142.330 3.555 144.710 4.280 ;
        RECT 145.550 3.555 147.930 4.280 ;
        RECT 148.770 3.555 151.150 4.280 ;
        RECT 151.990 3.555 157.590 4.280 ;
        RECT 158.430 3.555 160.810 4.280 ;
        RECT 161.650 3.555 164.030 4.280 ;
        RECT 164.870 3.555 167.250 4.280 ;
        RECT 168.090 3.555 170.470 4.280 ;
        RECT 171.310 3.555 173.690 4.280 ;
        RECT 174.530 3.555 176.910 4.280 ;
      LAYER met3 ;
        RECT 4.400 176.440 175.600 177.305 ;
        RECT 4.000 174.440 176.000 176.440 ;
        RECT 4.400 173.040 175.600 174.440 ;
        RECT 4.000 171.040 176.000 173.040 ;
        RECT 4.400 169.640 175.600 171.040 ;
        RECT 4.000 167.640 176.000 169.640 ;
        RECT 4.400 166.240 175.600 167.640 ;
        RECT 4.000 160.840 176.000 166.240 ;
        RECT 4.400 159.440 175.600 160.840 ;
        RECT 4.000 157.440 176.000 159.440 ;
        RECT 4.400 156.040 175.600 157.440 ;
        RECT 4.000 154.040 176.000 156.040 ;
        RECT 4.400 152.640 175.600 154.040 ;
        RECT 4.000 150.640 176.000 152.640 ;
        RECT 4.400 149.240 175.600 150.640 ;
        RECT 4.000 147.240 176.000 149.240 ;
        RECT 4.400 145.840 175.600 147.240 ;
        RECT 4.000 143.840 176.000 145.840 ;
        RECT 4.400 142.440 175.600 143.840 ;
        RECT 4.000 140.440 176.000 142.440 ;
        RECT 4.400 139.040 175.600 140.440 ;
        RECT 4.000 133.640 176.000 139.040 ;
        RECT 4.400 132.240 175.600 133.640 ;
        RECT 4.000 130.240 176.000 132.240 ;
        RECT 4.400 128.840 175.600 130.240 ;
        RECT 4.000 126.840 176.000 128.840 ;
        RECT 4.400 125.440 175.600 126.840 ;
        RECT 4.000 123.440 176.000 125.440 ;
        RECT 4.400 122.040 175.600 123.440 ;
        RECT 4.000 120.040 176.000 122.040 ;
        RECT 4.400 118.640 175.600 120.040 ;
        RECT 4.000 116.640 176.000 118.640 ;
        RECT 4.400 115.240 175.600 116.640 ;
        RECT 4.000 113.240 176.000 115.240 ;
        RECT 4.400 111.840 175.600 113.240 ;
        RECT 4.000 106.440 176.000 111.840 ;
        RECT 4.400 105.040 175.600 106.440 ;
        RECT 4.000 103.040 176.000 105.040 ;
        RECT 4.400 101.640 175.600 103.040 ;
        RECT 4.000 99.640 176.000 101.640 ;
        RECT 4.400 98.240 175.600 99.640 ;
        RECT 4.000 96.240 176.000 98.240 ;
        RECT 4.400 94.840 175.600 96.240 ;
        RECT 4.000 92.840 176.000 94.840 ;
        RECT 4.400 91.440 175.600 92.840 ;
        RECT 4.000 89.440 176.000 91.440 ;
        RECT 4.400 88.040 175.600 89.440 ;
        RECT 4.000 86.040 176.000 88.040 ;
        RECT 4.400 84.640 175.600 86.040 ;
        RECT 4.000 79.240 176.000 84.640 ;
        RECT 4.400 77.840 175.600 79.240 ;
        RECT 4.000 75.840 176.000 77.840 ;
        RECT 4.400 74.440 175.600 75.840 ;
        RECT 4.000 72.440 176.000 74.440 ;
        RECT 4.400 71.040 175.600 72.440 ;
        RECT 4.000 69.040 176.000 71.040 ;
        RECT 4.400 67.640 175.600 69.040 ;
        RECT 4.000 65.640 176.000 67.640 ;
        RECT 4.400 64.240 175.600 65.640 ;
        RECT 4.000 62.240 176.000 64.240 ;
        RECT 4.400 60.840 175.600 62.240 ;
        RECT 4.000 58.840 176.000 60.840 ;
        RECT 4.400 57.440 175.600 58.840 ;
        RECT 4.000 52.040 176.000 57.440 ;
        RECT 4.400 50.640 175.600 52.040 ;
        RECT 4.000 48.640 176.000 50.640 ;
        RECT 4.400 47.240 175.600 48.640 ;
        RECT 4.000 45.240 176.000 47.240 ;
        RECT 4.400 43.840 175.600 45.240 ;
        RECT 4.000 41.840 176.000 43.840 ;
        RECT 4.400 40.440 175.600 41.840 ;
        RECT 4.000 38.440 176.000 40.440 ;
        RECT 4.400 37.040 175.600 38.440 ;
        RECT 4.000 35.040 176.000 37.040 ;
        RECT 4.400 33.640 175.600 35.040 ;
        RECT 4.000 31.640 176.000 33.640 ;
        RECT 4.400 30.240 175.600 31.640 ;
        RECT 4.000 24.840 176.000 30.240 ;
        RECT 4.400 23.440 175.600 24.840 ;
        RECT 4.000 21.440 176.000 23.440 ;
        RECT 4.400 20.040 175.600 21.440 ;
        RECT 4.000 18.040 176.000 20.040 ;
        RECT 4.400 16.640 175.600 18.040 ;
        RECT 4.000 14.640 176.000 16.640 ;
        RECT 4.400 13.240 175.600 14.640 ;
        RECT 4.000 11.240 176.000 13.240 ;
        RECT 4.400 9.840 175.600 11.240 ;
        RECT 4.000 7.840 176.000 9.840 ;
        RECT 4.400 6.440 175.600 7.840 ;
        RECT 4.000 4.440 176.000 6.440 ;
        RECT 4.400 3.575 175.600 4.440 ;
  END
END WBM_DBus
END LIBRARY

