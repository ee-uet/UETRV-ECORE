magic
tech sky130A
magscale 1 2
timestamp 1647842912
<< obsli1 >>
rect 1104 2159 218868 217617
<< obsm1 >>
rect 1104 2128 218868 217796
<< metal2 >>
rect 1122 219200 1178 220000
rect 3422 219200 3478 220000
rect 5722 219200 5778 220000
rect 8022 219200 8078 220000
rect 10322 219200 10378 220000
rect 12622 219200 12678 220000
rect 15014 219200 15070 220000
rect 17314 219200 17370 220000
rect 19614 219200 19670 220000
rect 21914 219200 21970 220000
rect 24214 219200 24270 220000
rect 26514 219200 26570 220000
rect 28906 219200 28962 220000
rect 31206 219200 31262 220000
rect 33506 219200 33562 220000
rect 35806 219200 35862 220000
rect 38106 219200 38162 220000
rect 40406 219200 40462 220000
rect 42798 219200 42854 220000
rect 45098 219200 45154 220000
rect 47398 219200 47454 220000
rect 49698 219200 49754 220000
rect 51998 219200 52054 220000
rect 54298 219200 54354 220000
rect 56690 219200 56746 220000
rect 58990 219200 59046 220000
rect 61290 219200 61346 220000
rect 63590 219200 63646 220000
rect 65890 219200 65946 220000
rect 68190 219200 68246 220000
rect 70582 219200 70638 220000
rect 72882 219200 72938 220000
rect 75182 219200 75238 220000
rect 77482 219200 77538 220000
rect 79782 219200 79838 220000
rect 82082 219200 82138 220000
rect 84474 219200 84530 220000
rect 86774 219200 86830 220000
rect 89074 219200 89130 220000
rect 91374 219200 91430 220000
rect 93674 219200 93730 220000
rect 95974 219200 96030 220000
rect 98366 219200 98422 220000
rect 100666 219200 100722 220000
rect 102966 219200 103022 220000
rect 105266 219200 105322 220000
rect 107566 219200 107622 220000
rect 109866 219200 109922 220000
rect 112258 219200 112314 220000
rect 114558 219200 114614 220000
rect 116858 219200 116914 220000
rect 119158 219200 119214 220000
rect 121458 219200 121514 220000
rect 123758 219200 123814 220000
rect 126150 219200 126206 220000
rect 128450 219200 128506 220000
rect 130750 219200 130806 220000
rect 133050 219200 133106 220000
rect 135350 219200 135406 220000
rect 137650 219200 137706 220000
rect 140042 219200 140098 220000
rect 142342 219200 142398 220000
rect 144642 219200 144698 220000
rect 146942 219200 146998 220000
rect 149242 219200 149298 220000
rect 151542 219200 151598 220000
rect 153934 219200 153990 220000
rect 156234 219200 156290 220000
rect 158534 219200 158590 220000
rect 160834 219200 160890 220000
rect 163134 219200 163190 220000
rect 165434 219200 165490 220000
rect 167826 219200 167882 220000
rect 170126 219200 170182 220000
rect 172426 219200 172482 220000
rect 174726 219200 174782 220000
rect 177026 219200 177082 220000
rect 179326 219200 179382 220000
rect 181718 219200 181774 220000
rect 184018 219200 184074 220000
rect 186318 219200 186374 220000
rect 188618 219200 188674 220000
rect 190918 219200 190974 220000
rect 193218 219200 193274 220000
rect 195610 219200 195666 220000
rect 197910 219200 197966 220000
rect 200210 219200 200266 220000
rect 202510 219200 202566 220000
rect 204810 219200 204866 220000
rect 207110 219200 207166 220000
rect 209502 219200 209558 220000
rect 211802 219200 211858 220000
rect 214102 219200 214158 220000
rect 216402 219200 216458 220000
rect 218702 219200 218758 220000
rect 5446 0 5502 800
rect 16394 0 16450 800
rect 27434 0 27490 800
rect 38382 0 38438 800
rect 49422 0 49478 800
rect 60370 0 60426 800
rect 71410 0 71466 800
rect 82358 0 82414 800
rect 93398 0 93454 800
rect 104346 0 104402 800
rect 115386 0 115442 800
rect 126426 0 126482 800
rect 137374 0 137430 800
rect 148414 0 148470 800
rect 159362 0 159418 800
rect 170402 0 170458 800
rect 181350 0 181406 800
rect 192390 0 192446 800
rect 203338 0 203394 800
rect 214378 0 214434 800
<< obsm2 >>
rect 1234 219144 3366 219473
rect 3534 219144 5666 219473
rect 5834 219144 7966 219473
rect 8134 219144 10266 219473
rect 10434 219144 12566 219473
rect 12734 219144 14958 219473
rect 15126 219144 17258 219473
rect 17426 219144 19558 219473
rect 19726 219144 21858 219473
rect 22026 219144 24158 219473
rect 24326 219144 26458 219473
rect 26626 219144 28850 219473
rect 29018 219144 31150 219473
rect 31318 219144 33450 219473
rect 33618 219144 35750 219473
rect 35918 219144 38050 219473
rect 38218 219144 40350 219473
rect 40518 219144 42742 219473
rect 42910 219144 45042 219473
rect 45210 219144 47342 219473
rect 47510 219144 49642 219473
rect 49810 219144 51942 219473
rect 52110 219144 54242 219473
rect 54410 219144 56634 219473
rect 56802 219144 58934 219473
rect 59102 219144 61234 219473
rect 61402 219144 63534 219473
rect 63702 219144 65834 219473
rect 66002 219144 68134 219473
rect 68302 219144 70526 219473
rect 70694 219144 72826 219473
rect 72994 219144 75126 219473
rect 75294 219144 77426 219473
rect 77594 219144 79726 219473
rect 79894 219144 82026 219473
rect 82194 219144 84418 219473
rect 84586 219144 86718 219473
rect 86886 219144 89018 219473
rect 89186 219144 91318 219473
rect 91486 219144 93618 219473
rect 93786 219144 95918 219473
rect 96086 219144 98310 219473
rect 98478 219144 100610 219473
rect 100778 219144 102910 219473
rect 103078 219144 105210 219473
rect 105378 219144 107510 219473
rect 107678 219144 109810 219473
rect 109978 219144 112202 219473
rect 112370 219144 114502 219473
rect 114670 219144 116802 219473
rect 116970 219144 119102 219473
rect 119270 219144 121402 219473
rect 121570 219144 123702 219473
rect 123870 219144 126094 219473
rect 126262 219144 128394 219473
rect 128562 219144 130694 219473
rect 130862 219144 132994 219473
rect 133162 219144 135294 219473
rect 135462 219144 137594 219473
rect 137762 219144 139986 219473
rect 140154 219144 142286 219473
rect 142454 219144 144586 219473
rect 144754 219144 146886 219473
rect 147054 219144 149186 219473
rect 149354 219144 151486 219473
rect 151654 219144 153878 219473
rect 154046 219144 156178 219473
rect 156346 219144 158478 219473
rect 158646 219144 160778 219473
rect 160946 219144 163078 219473
rect 163246 219144 165378 219473
rect 165546 219144 167770 219473
rect 167938 219144 170070 219473
rect 170238 219144 172370 219473
rect 172538 219144 174670 219473
rect 174838 219144 176970 219473
rect 177138 219144 179270 219473
rect 179438 219144 181662 219473
rect 181830 219144 183962 219473
rect 184130 219144 186262 219473
rect 186430 219144 188562 219473
rect 188730 219144 190862 219473
rect 191030 219144 193162 219473
rect 193330 219144 195554 219473
rect 195722 219144 197854 219473
rect 198022 219144 200154 219473
rect 200322 219144 202454 219473
rect 202622 219144 204754 219473
rect 204922 219144 207054 219473
rect 207222 219144 209446 219473
rect 209614 219144 211746 219473
rect 211914 219144 214046 219473
rect 214214 219144 216346 219473
rect 216514 219144 218646 219473
rect 1124 856 218756 219144
rect 1124 575 5390 856
rect 5558 575 16338 856
rect 16506 575 27378 856
rect 27546 575 38326 856
rect 38494 575 49366 856
rect 49534 575 60314 856
rect 60482 575 71354 856
rect 71522 575 82302 856
rect 82470 575 93342 856
rect 93510 575 104290 856
rect 104458 575 115330 856
rect 115498 575 126370 856
rect 126538 575 137318 856
rect 137486 575 148358 856
rect 148526 575 159306 856
rect 159474 575 170346 856
rect 170514 575 181294 856
rect 181462 575 192334 856
rect 192502 575 203282 856
rect 203450 575 214322 856
rect 214490 575 218756 856
<< metal3 >>
rect 0 219376 800 219496
rect 219200 218968 220000 219088
rect 0 218152 800 218272
rect 0 217064 800 217184
rect 219200 217064 220000 217184
rect 0 215840 800 215960
rect 219200 215160 220000 215280
rect 0 214752 800 214872
rect 0 213528 800 213648
rect 219200 213256 220000 213376
rect 0 212440 800 212560
rect 0 211216 800 211336
rect 219200 211352 220000 211472
rect 0 209992 800 210112
rect 219200 209448 220000 209568
rect 0 208904 800 209024
rect 0 207680 800 207800
rect 219200 207544 220000 207664
rect 0 206592 800 206712
rect 219200 205640 220000 205760
rect 0 205368 800 205488
rect 0 204280 800 204400
rect 219200 203736 220000 203856
rect 0 203056 800 203176
rect 0 201968 800 202088
rect 219200 201832 220000 201952
rect 0 200744 800 200864
rect 219200 199928 220000 200048
rect 0 199520 800 199640
rect 0 198432 800 198552
rect 219200 198024 220000 198144
rect 0 197208 800 197328
rect 0 196120 800 196240
rect 219200 196120 220000 196240
rect 0 194896 800 195016
rect 219200 194216 220000 194336
rect 0 193808 800 193928
rect 0 192584 800 192704
rect 219200 192312 220000 192432
rect 0 191360 800 191480
rect 0 190272 800 190392
rect 219200 190408 220000 190528
rect 0 189048 800 189168
rect 219200 188504 220000 188624
rect 0 187960 800 188080
rect 0 186736 800 186856
rect 219200 186600 220000 186720
rect 0 185648 800 185768
rect 219200 184696 220000 184816
rect 0 184424 800 184544
rect 0 183336 800 183456
rect 219200 182928 220000 183048
rect 0 182112 800 182232
rect 0 180888 800 181008
rect 219200 181024 220000 181144
rect 0 179800 800 179920
rect 219200 179120 220000 179240
rect 0 178576 800 178696
rect 0 177488 800 177608
rect 219200 177216 220000 177336
rect 0 176264 800 176384
rect 0 175176 800 175296
rect 219200 175312 220000 175432
rect 0 173952 800 174072
rect 219200 173408 220000 173528
rect 0 172864 800 172984
rect 0 171640 800 171760
rect 219200 171504 220000 171624
rect 0 170416 800 170536
rect 219200 169600 220000 169720
rect 0 169328 800 169448
rect 0 168104 800 168224
rect 219200 167696 220000 167816
rect 0 167016 800 167136
rect 0 165792 800 165912
rect 219200 165792 220000 165912
rect 0 164704 800 164824
rect 219200 163888 220000 164008
rect 0 163480 800 163600
rect 0 162256 800 162376
rect 219200 161984 220000 162104
rect 0 161168 800 161288
rect 0 159944 800 160064
rect 219200 160080 220000 160200
rect 0 158856 800 158976
rect 219200 158176 220000 158296
rect 0 157632 800 157752
rect 0 156544 800 156664
rect 219200 156272 220000 156392
rect 0 155320 800 155440
rect 0 154232 800 154352
rect 219200 154368 220000 154488
rect 0 153008 800 153128
rect 219200 152464 220000 152584
rect 0 151784 800 151904
rect 0 150696 800 150816
rect 219200 150560 220000 150680
rect 0 149472 800 149592
rect 219200 148656 220000 148776
rect 0 148384 800 148504
rect 0 147160 800 147280
rect 219200 146888 220000 147008
rect 0 146072 800 146192
rect 0 144848 800 144968
rect 219200 144984 220000 145104
rect 0 143624 800 143744
rect 219200 143080 220000 143200
rect 0 142536 800 142656
rect 0 141312 800 141432
rect 219200 141176 220000 141296
rect 0 140224 800 140344
rect 219200 139272 220000 139392
rect 0 139000 800 139120
rect 0 137912 800 138032
rect 219200 137368 220000 137488
rect 0 136688 800 136808
rect 0 135600 800 135720
rect 219200 135464 220000 135584
rect 0 134376 800 134496
rect 219200 133560 220000 133680
rect 0 133152 800 133272
rect 0 132064 800 132184
rect 219200 131656 220000 131776
rect 0 130840 800 130960
rect 0 129752 800 129872
rect 219200 129752 220000 129872
rect 0 128528 800 128648
rect 219200 127848 220000 127968
rect 0 127440 800 127560
rect 0 126216 800 126336
rect 219200 125944 220000 126064
rect 0 125128 800 125248
rect 0 123904 800 124024
rect 219200 124040 220000 124160
rect 0 122680 800 122800
rect 219200 122136 220000 122256
rect 0 121592 800 121712
rect 0 120368 800 120488
rect 219200 120232 220000 120352
rect 0 119280 800 119400
rect 219200 118328 220000 118448
rect 0 118056 800 118176
rect 0 116968 800 117088
rect 219200 116424 220000 116544
rect 0 115744 800 115864
rect 0 114520 800 114640
rect 219200 114520 220000 114640
rect 0 113432 800 113552
rect 219200 112616 220000 112736
rect 0 112208 800 112328
rect 0 111120 800 111240
rect 219200 110848 220000 110968
rect 0 109896 800 110016
rect 0 108808 800 108928
rect 219200 108944 220000 109064
rect 0 107584 800 107704
rect 219200 107040 220000 107160
rect 0 106496 800 106616
rect 0 105272 800 105392
rect 219200 105136 220000 105256
rect 0 104048 800 104168
rect 219200 103232 220000 103352
rect 0 102960 800 103080
rect 0 101736 800 101856
rect 219200 101328 220000 101448
rect 0 100648 800 100768
rect 0 99424 800 99544
rect 219200 99424 220000 99544
rect 0 98336 800 98456
rect 219200 97520 220000 97640
rect 0 97112 800 97232
rect 0 95888 800 96008
rect 219200 95616 220000 95736
rect 0 94800 800 94920
rect 0 93576 800 93696
rect 219200 93712 220000 93832
rect 0 92488 800 92608
rect 219200 91808 220000 91928
rect 0 91264 800 91384
rect 0 90176 800 90296
rect 219200 89904 220000 90024
rect 0 88952 800 89072
rect 0 87864 800 87984
rect 219200 88000 220000 88120
rect 0 86640 800 86760
rect 219200 86096 220000 86216
rect 0 85416 800 85536
rect 0 84328 800 84448
rect 219200 84192 220000 84312
rect 0 83104 800 83224
rect 219200 82288 220000 82408
rect 0 82016 800 82136
rect 0 80792 800 80912
rect 219200 80384 220000 80504
rect 0 79704 800 79824
rect 0 78480 800 78600
rect 219200 78480 220000 78600
rect 0 77392 800 77512
rect 219200 76576 220000 76696
rect 0 76168 800 76288
rect 0 74944 800 75064
rect 219200 74672 220000 74792
rect 0 73856 800 73976
rect 219200 72904 220000 73024
rect 0 72632 800 72752
rect 0 71544 800 71664
rect 219200 71000 220000 71120
rect 0 70320 800 70440
rect 0 69232 800 69352
rect 219200 69096 220000 69216
rect 0 68008 800 68128
rect 219200 67192 220000 67312
rect 0 66784 800 66904
rect 0 65696 800 65816
rect 219200 65288 220000 65408
rect 0 64472 800 64592
rect 0 63384 800 63504
rect 219200 63384 220000 63504
rect 0 62160 800 62280
rect 219200 61480 220000 61600
rect 0 61072 800 61192
rect 0 59848 800 59968
rect 219200 59576 220000 59696
rect 0 58760 800 58880
rect 0 57536 800 57656
rect 219200 57672 220000 57792
rect 0 56312 800 56432
rect 219200 55768 220000 55888
rect 0 55224 800 55344
rect 0 54000 800 54120
rect 219200 53864 220000 53984
rect 0 52912 800 53032
rect 219200 51960 220000 52080
rect 0 51688 800 51808
rect 0 50600 800 50720
rect 219200 50056 220000 50176
rect 0 49376 800 49496
rect 0 48152 800 48272
rect 219200 48152 220000 48272
rect 0 47064 800 47184
rect 219200 46248 220000 46368
rect 0 45840 800 45960
rect 0 44752 800 44872
rect 219200 44344 220000 44464
rect 0 43528 800 43648
rect 0 42440 800 42560
rect 219200 42440 220000 42560
rect 0 41216 800 41336
rect 219200 40536 220000 40656
rect 0 40128 800 40248
rect 0 38904 800 39024
rect 219200 38632 220000 38752
rect 0 37680 800 37800
rect 219200 36864 220000 36984
rect 0 36592 800 36712
rect 0 35368 800 35488
rect 219200 34960 220000 35080
rect 0 34280 800 34400
rect 0 33056 800 33176
rect 219200 33056 220000 33176
rect 0 31968 800 32088
rect 219200 31152 220000 31272
rect 0 30744 800 30864
rect 0 29656 800 29776
rect 219200 29248 220000 29368
rect 0 28432 800 28552
rect 0 27208 800 27328
rect 219200 27344 220000 27464
rect 0 26120 800 26240
rect 219200 25440 220000 25560
rect 0 24896 800 25016
rect 0 23808 800 23928
rect 219200 23536 220000 23656
rect 0 22584 800 22704
rect 0 21496 800 21616
rect 219200 21632 220000 21752
rect 0 20272 800 20392
rect 219200 19728 220000 19848
rect 0 19048 800 19168
rect 0 17960 800 18080
rect 219200 17824 220000 17944
rect 0 16736 800 16856
rect 219200 15920 220000 16040
rect 0 15648 800 15768
rect 0 14424 800 14544
rect 219200 14016 220000 14136
rect 0 13336 800 13456
rect 0 12112 800 12232
rect 219200 12112 220000 12232
rect 0 11024 800 11144
rect 219200 10208 220000 10328
rect 0 9800 800 9920
rect 0 8576 800 8696
rect 219200 8304 220000 8424
rect 0 7488 800 7608
rect 0 6264 800 6384
rect 219200 6400 220000 6520
rect 0 5176 800 5296
rect 219200 4496 220000 4616
rect 0 3952 800 4072
rect 0 2864 800 2984
rect 219200 2592 220000 2712
rect 0 1640 800 1760
rect 219200 824 220000 944
rect 0 552 800 672
<< obsm3 >>
rect 880 219296 219200 219469
rect 800 219168 219200 219296
rect 800 218888 219120 219168
rect 800 218352 219200 218888
rect 880 218072 219200 218352
rect 800 217264 219200 218072
rect 880 216984 219120 217264
rect 800 216040 219200 216984
rect 880 215760 219200 216040
rect 800 215360 219200 215760
rect 800 215080 219120 215360
rect 800 214952 219200 215080
rect 880 214672 219200 214952
rect 800 213728 219200 214672
rect 880 213456 219200 213728
rect 880 213448 219120 213456
rect 800 213176 219120 213448
rect 800 212640 219200 213176
rect 880 212360 219200 212640
rect 800 211552 219200 212360
rect 800 211416 219120 211552
rect 880 211272 219120 211416
rect 880 211136 219200 211272
rect 800 210192 219200 211136
rect 880 209912 219200 210192
rect 800 209648 219200 209912
rect 800 209368 219120 209648
rect 800 209104 219200 209368
rect 880 208824 219200 209104
rect 800 207880 219200 208824
rect 880 207744 219200 207880
rect 880 207600 219120 207744
rect 800 207464 219120 207600
rect 800 206792 219200 207464
rect 880 206512 219200 206792
rect 800 205840 219200 206512
rect 800 205568 219120 205840
rect 880 205560 219120 205568
rect 880 205288 219200 205560
rect 800 204480 219200 205288
rect 880 204200 219200 204480
rect 800 203936 219200 204200
rect 800 203656 219120 203936
rect 800 203256 219200 203656
rect 880 202976 219200 203256
rect 800 202168 219200 202976
rect 880 202032 219200 202168
rect 880 201888 219120 202032
rect 800 201752 219120 201888
rect 800 200944 219200 201752
rect 880 200664 219200 200944
rect 800 200128 219200 200664
rect 800 199848 219120 200128
rect 800 199720 219200 199848
rect 880 199440 219200 199720
rect 800 198632 219200 199440
rect 880 198352 219200 198632
rect 800 198224 219200 198352
rect 800 197944 219120 198224
rect 800 197408 219200 197944
rect 880 197128 219200 197408
rect 800 196320 219200 197128
rect 880 196040 219120 196320
rect 800 195096 219200 196040
rect 880 194816 219200 195096
rect 800 194416 219200 194816
rect 800 194136 219120 194416
rect 800 194008 219200 194136
rect 880 193728 219200 194008
rect 800 192784 219200 193728
rect 880 192512 219200 192784
rect 880 192504 219120 192512
rect 800 192232 219120 192504
rect 800 191560 219200 192232
rect 880 191280 219200 191560
rect 800 190608 219200 191280
rect 800 190472 219120 190608
rect 880 190328 219120 190472
rect 880 190192 219200 190328
rect 800 189248 219200 190192
rect 880 188968 219200 189248
rect 800 188704 219200 188968
rect 800 188424 219120 188704
rect 800 188160 219200 188424
rect 880 187880 219200 188160
rect 800 186936 219200 187880
rect 880 186800 219200 186936
rect 880 186656 219120 186800
rect 800 186520 219120 186656
rect 800 185848 219200 186520
rect 880 185568 219200 185848
rect 800 184896 219200 185568
rect 800 184624 219120 184896
rect 880 184616 219120 184624
rect 880 184344 219200 184616
rect 800 183536 219200 184344
rect 880 183256 219200 183536
rect 800 183128 219200 183256
rect 800 182848 219120 183128
rect 800 182312 219200 182848
rect 880 182032 219200 182312
rect 800 181224 219200 182032
rect 800 181088 219120 181224
rect 880 180944 219120 181088
rect 880 180808 219200 180944
rect 800 180000 219200 180808
rect 880 179720 219200 180000
rect 800 179320 219200 179720
rect 800 179040 219120 179320
rect 800 178776 219200 179040
rect 880 178496 219200 178776
rect 800 177688 219200 178496
rect 880 177416 219200 177688
rect 880 177408 219120 177416
rect 800 177136 219120 177408
rect 800 176464 219200 177136
rect 880 176184 219200 176464
rect 800 175512 219200 176184
rect 800 175376 219120 175512
rect 880 175232 219120 175376
rect 880 175096 219200 175232
rect 800 174152 219200 175096
rect 880 173872 219200 174152
rect 800 173608 219200 173872
rect 800 173328 219120 173608
rect 800 173064 219200 173328
rect 880 172784 219200 173064
rect 800 171840 219200 172784
rect 880 171704 219200 171840
rect 880 171560 219120 171704
rect 800 171424 219120 171560
rect 800 170616 219200 171424
rect 880 170336 219200 170616
rect 800 169800 219200 170336
rect 800 169528 219120 169800
rect 880 169520 219120 169528
rect 880 169248 219200 169520
rect 800 168304 219200 169248
rect 880 168024 219200 168304
rect 800 167896 219200 168024
rect 800 167616 219120 167896
rect 800 167216 219200 167616
rect 880 166936 219200 167216
rect 800 165992 219200 166936
rect 880 165712 219120 165992
rect 800 164904 219200 165712
rect 880 164624 219200 164904
rect 800 164088 219200 164624
rect 800 163808 219120 164088
rect 800 163680 219200 163808
rect 880 163400 219200 163680
rect 800 162456 219200 163400
rect 880 162184 219200 162456
rect 880 162176 219120 162184
rect 800 161904 219120 162176
rect 800 161368 219200 161904
rect 880 161088 219200 161368
rect 800 160280 219200 161088
rect 800 160144 219120 160280
rect 880 160000 219120 160144
rect 880 159864 219200 160000
rect 800 159056 219200 159864
rect 880 158776 219200 159056
rect 800 158376 219200 158776
rect 800 158096 219120 158376
rect 800 157832 219200 158096
rect 880 157552 219200 157832
rect 800 156744 219200 157552
rect 880 156472 219200 156744
rect 880 156464 219120 156472
rect 800 156192 219120 156464
rect 800 155520 219200 156192
rect 880 155240 219200 155520
rect 800 154568 219200 155240
rect 800 154432 219120 154568
rect 880 154288 219120 154432
rect 880 154152 219200 154288
rect 800 153208 219200 154152
rect 880 152928 219200 153208
rect 800 152664 219200 152928
rect 800 152384 219120 152664
rect 800 151984 219200 152384
rect 880 151704 219200 151984
rect 800 150896 219200 151704
rect 880 150760 219200 150896
rect 880 150616 219120 150760
rect 800 150480 219120 150616
rect 800 149672 219200 150480
rect 880 149392 219200 149672
rect 800 148856 219200 149392
rect 800 148584 219120 148856
rect 880 148576 219120 148584
rect 880 148304 219200 148576
rect 800 147360 219200 148304
rect 880 147088 219200 147360
rect 880 147080 219120 147088
rect 800 146808 219120 147080
rect 800 146272 219200 146808
rect 880 145992 219200 146272
rect 800 145184 219200 145992
rect 800 145048 219120 145184
rect 880 144904 219120 145048
rect 880 144768 219200 144904
rect 800 143824 219200 144768
rect 880 143544 219200 143824
rect 800 143280 219200 143544
rect 800 143000 219120 143280
rect 800 142736 219200 143000
rect 880 142456 219200 142736
rect 800 141512 219200 142456
rect 880 141376 219200 141512
rect 880 141232 219120 141376
rect 800 141096 219120 141232
rect 800 140424 219200 141096
rect 880 140144 219200 140424
rect 800 139472 219200 140144
rect 800 139200 219120 139472
rect 880 139192 219120 139200
rect 880 138920 219200 139192
rect 800 138112 219200 138920
rect 880 137832 219200 138112
rect 800 137568 219200 137832
rect 800 137288 219120 137568
rect 800 136888 219200 137288
rect 880 136608 219200 136888
rect 800 135800 219200 136608
rect 880 135664 219200 135800
rect 880 135520 219120 135664
rect 800 135384 219120 135520
rect 800 134576 219200 135384
rect 880 134296 219200 134576
rect 800 133760 219200 134296
rect 800 133480 219120 133760
rect 800 133352 219200 133480
rect 880 133072 219200 133352
rect 800 132264 219200 133072
rect 880 131984 219200 132264
rect 800 131856 219200 131984
rect 800 131576 219120 131856
rect 800 131040 219200 131576
rect 880 130760 219200 131040
rect 800 129952 219200 130760
rect 880 129672 219120 129952
rect 800 128728 219200 129672
rect 880 128448 219200 128728
rect 800 128048 219200 128448
rect 800 127768 219120 128048
rect 800 127640 219200 127768
rect 880 127360 219200 127640
rect 800 126416 219200 127360
rect 880 126144 219200 126416
rect 880 126136 219120 126144
rect 800 125864 219120 126136
rect 800 125328 219200 125864
rect 880 125048 219200 125328
rect 800 124240 219200 125048
rect 800 124104 219120 124240
rect 880 123960 219120 124104
rect 880 123824 219200 123960
rect 800 122880 219200 123824
rect 880 122600 219200 122880
rect 800 122336 219200 122600
rect 800 122056 219120 122336
rect 800 121792 219200 122056
rect 880 121512 219200 121792
rect 800 120568 219200 121512
rect 880 120432 219200 120568
rect 880 120288 219120 120432
rect 800 120152 219120 120288
rect 800 119480 219200 120152
rect 880 119200 219200 119480
rect 800 118528 219200 119200
rect 800 118256 219120 118528
rect 880 118248 219120 118256
rect 880 117976 219200 118248
rect 800 117168 219200 117976
rect 880 116888 219200 117168
rect 800 116624 219200 116888
rect 800 116344 219120 116624
rect 800 115944 219200 116344
rect 880 115664 219200 115944
rect 800 114720 219200 115664
rect 880 114440 219120 114720
rect 800 113632 219200 114440
rect 880 113352 219200 113632
rect 800 112816 219200 113352
rect 800 112536 219120 112816
rect 800 112408 219200 112536
rect 880 112128 219200 112408
rect 800 111320 219200 112128
rect 880 111048 219200 111320
rect 880 111040 219120 111048
rect 800 110768 219120 111040
rect 800 110096 219200 110768
rect 880 109816 219200 110096
rect 800 109144 219200 109816
rect 800 109008 219120 109144
rect 880 108864 219120 109008
rect 880 108728 219200 108864
rect 800 107784 219200 108728
rect 880 107504 219200 107784
rect 800 107240 219200 107504
rect 800 106960 219120 107240
rect 800 106696 219200 106960
rect 880 106416 219200 106696
rect 800 105472 219200 106416
rect 880 105336 219200 105472
rect 880 105192 219120 105336
rect 800 105056 219120 105192
rect 800 104248 219200 105056
rect 880 103968 219200 104248
rect 800 103432 219200 103968
rect 800 103160 219120 103432
rect 880 103152 219120 103160
rect 880 102880 219200 103152
rect 800 101936 219200 102880
rect 880 101656 219200 101936
rect 800 101528 219200 101656
rect 800 101248 219120 101528
rect 800 100848 219200 101248
rect 880 100568 219200 100848
rect 800 99624 219200 100568
rect 880 99344 219120 99624
rect 800 98536 219200 99344
rect 880 98256 219200 98536
rect 800 97720 219200 98256
rect 800 97440 219120 97720
rect 800 97312 219200 97440
rect 880 97032 219200 97312
rect 800 96088 219200 97032
rect 880 95816 219200 96088
rect 880 95808 219120 95816
rect 800 95536 219120 95808
rect 800 95000 219200 95536
rect 880 94720 219200 95000
rect 800 93912 219200 94720
rect 800 93776 219120 93912
rect 880 93632 219120 93776
rect 880 93496 219200 93632
rect 800 92688 219200 93496
rect 880 92408 219200 92688
rect 800 92008 219200 92408
rect 800 91728 219120 92008
rect 800 91464 219200 91728
rect 880 91184 219200 91464
rect 800 90376 219200 91184
rect 880 90104 219200 90376
rect 880 90096 219120 90104
rect 800 89824 219120 90096
rect 800 89152 219200 89824
rect 880 88872 219200 89152
rect 800 88200 219200 88872
rect 800 88064 219120 88200
rect 880 87920 219120 88064
rect 880 87784 219200 87920
rect 800 86840 219200 87784
rect 880 86560 219200 86840
rect 800 86296 219200 86560
rect 800 86016 219120 86296
rect 800 85616 219200 86016
rect 880 85336 219200 85616
rect 800 84528 219200 85336
rect 880 84392 219200 84528
rect 880 84248 219120 84392
rect 800 84112 219120 84248
rect 800 83304 219200 84112
rect 880 83024 219200 83304
rect 800 82488 219200 83024
rect 800 82216 219120 82488
rect 880 82208 219120 82216
rect 880 81936 219200 82208
rect 800 80992 219200 81936
rect 880 80712 219200 80992
rect 800 80584 219200 80712
rect 800 80304 219120 80584
rect 800 79904 219200 80304
rect 880 79624 219200 79904
rect 800 78680 219200 79624
rect 880 78400 219120 78680
rect 800 77592 219200 78400
rect 880 77312 219200 77592
rect 800 76776 219200 77312
rect 800 76496 219120 76776
rect 800 76368 219200 76496
rect 880 76088 219200 76368
rect 800 75144 219200 76088
rect 880 74872 219200 75144
rect 880 74864 219120 74872
rect 800 74592 219120 74864
rect 800 74056 219200 74592
rect 880 73776 219200 74056
rect 800 73104 219200 73776
rect 800 72832 219120 73104
rect 880 72824 219120 72832
rect 880 72552 219200 72824
rect 800 71744 219200 72552
rect 880 71464 219200 71744
rect 800 71200 219200 71464
rect 800 70920 219120 71200
rect 800 70520 219200 70920
rect 880 70240 219200 70520
rect 800 69432 219200 70240
rect 880 69296 219200 69432
rect 880 69152 219120 69296
rect 800 69016 219120 69152
rect 800 68208 219200 69016
rect 880 67928 219200 68208
rect 800 67392 219200 67928
rect 800 67112 219120 67392
rect 800 66984 219200 67112
rect 880 66704 219200 66984
rect 800 65896 219200 66704
rect 880 65616 219200 65896
rect 800 65488 219200 65616
rect 800 65208 219120 65488
rect 800 64672 219200 65208
rect 880 64392 219200 64672
rect 800 63584 219200 64392
rect 880 63304 219120 63584
rect 800 62360 219200 63304
rect 880 62080 219200 62360
rect 800 61680 219200 62080
rect 800 61400 219120 61680
rect 800 61272 219200 61400
rect 880 60992 219200 61272
rect 800 60048 219200 60992
rect 880 59776 219200 60048
rect 880 59768 219120 59776
rect 800 59496 219120 59768
rect 800 58960 219200 59496
rect 880 58680 219200 58960
rect 800 57872 219200 58680
rect 800 57736 219120 57872
rect 880 57592 219120 57736
rect 880 57456 219200 57592
rect 800 56512 219200 57456
rect 880 56232 219200 56512
rect 800 55968 219200 56232
rect 800 55688 219120 55968
rect 800 55424 219200 55688
rect 880 55144 219200 55424
rect 800 54200 219200 55144
rect 880 54064 219200 54200
rect 880 53920 219120 54064
rect 800 53784 219120 53920
rect 800 53112 219200 53784
rect 880 52832 219200 53112
rect 800 52160 219200 52832
rect 800 51888 219120 52160
rect 880 51880 219120 51888
rect 880 51608 219200 51880
rect 800 50800 219200 51608
rect 880 50520 219200 50800
rect 800 50256 219200 50520
rect 800 49976 219120 50256
rect 800 49576 219200 49976
rect 880 49296 219200 49576
rect 800 48352 219200 49296
rect 880 48072 219120 48352
rect 800 47264 219200 48072
rect 880 46984 219200 47264
rect 800 46448 219200 46984
rect 800 46168 219120 46448
rect 800 46040 219200 46168
rect 880 45760 219200 46040
rect 800 44952 219200 45760
rect 880 44672 219200 44952
rect 800 44544 219200 44672
rect 800 44264 219120 44544
rect 800 43728 219200 44264
rect 880 43448 219200 43728
rect 800 42640 219200 43448
rect 880 42360 219120 42640
rect 800 41416 219200 42360
rect 880 41136 219200 41416
rect 800 40736 219200 41136
rect 800 40456 219120 40736
rect 800 40328 219200 40456
rect 880 40048 219200 40328
rect 800 39104 219200 40048
rect 880 38832 219200 39104
rect 880 38824 219120 38832
rect 800 38552 219120 38824
rect 800 37880 219200 38552
rect 880 37600 219200 37880
rect 800 37064 219200 37600
rect 800 36792 219120 37064
rect 880 36784 219120 36792
rect 880 36512 219200 36784
rect 800 35568 219200 36512
rect 880 35288 219200 35568
rect 800 35160 219200 35288
rect 800 34880 219120 35160
rect 800 34480 219200 34880
rect 880 34200 219200 34480
rect 800 33256 219200 34200
rect 880 32976 219120 33256
rect 800 32168 219200 32976
rect 880 31888 219200 32168
rect 800 31352 219200 31888
rect 800 31072 219120 31352
rect 800 30944 219200 31072
rect 880 30664 219200 30944
rect 800 29856 219200 30664
rect 880 29576 219200 29856
rect 800 29448 219200 29576
rect 800 29168 219120 29448
rect 800 28632 219200 29168
rect 880 28352 219200 28632
rect 800 27544 219200 28352
rect 800 27408 219120 27544
rect 880 27264 219120 27408
rect 880 27128 219200 27264
rect 800 26320 219200 27128
rect 880 26040 219200 26320
rect 800 25640 219200 26040
rect 800 25360 219120 25640
rect 800 25096 219200 25360
rect 880 24816 219200 25096
rect 800 24008 219200 24816
rect 880 23736 219200 24008
rect 880 23728 219120 23736
rect 800 23456 219120 23728
rect 800 22784 219200 23456
rect 880 22504 219200 22784
rect 800 21832 219200 22504
rect 800 21696 219120 21832
rect 880 21552 219120 21696
rect 880 21416 219200 21552
rect 800 20472 219200 21416
rect 880 20192 219200 20472
rect 800 19928 219200 20192
rect 800 19648 219120 19928
rect 800 19248 219200 19648
rect 880 18968 219200 19248
rect 800 18160 219200 18968
rect 880 18024 219200 18160
rect 880 17880 219120 18024
rect 800 17744 219120 17880
rect 800 16936 219200 17744
rect 880 16656 219200 16936
rect 800 16120 219200 16656
rect 800 15848 219120 16120
rect 880 15840 219120 15848
rect 880 15568 219200 15840
rect 800 14624 219200 15568
rect 880 14344 219200 14624
rect 800 14216 219200 14344
rect 800 13936 219120 14216
rect 800 13536 219200 13936
rect 880 13256 219200 13536
rect 800 12312 219200 13256
rect 880 12032 219120 12312
rect 800 11224 219200 12032
rect 880 10944 219200 11224
rect 800 10408 219200 10944
rect 800 10128 219120 10408
rect 800 10000 219200 10128
rect 880 9720 219200 10000
rect 800 8776 219200 9720
rect 880 8504 219200 8776
rect 880 8496 219120 8504
rect 800 8224 219120 8496
rect 800 7688 219200 8224
rect 880 7408 219200 7688
rect 800 6600 219200 7408
rect 800 6464 219120 6600
rect 880 6320 219120 6464
rect 880 6184 219200 6320
rect 800 5376 219200 6184
rect 880 5096 219200 5376
rect 800 4696 219200 5096
rect 800 4416 219120 4696
rect 800 4152 219200 4416
rect 880 3872 219200 4152
rect 800 3064 219200 3872
rect 880 2792 219200 3064
rect 880 2784 219120 2792
rect 800 2512 219120 2784
rect 800 1840 219200 2512
rect 880 1560 219200 1840
rect 800 1024 219200 1560
rect 800 752 219120 1024
rect 880 744 219120 752
rect 880 579 219200 744
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
rect 50288 2128 50608 217648
rect 65648 2128 65968 217648
rect 81008 2128 81328 217648
rect 96368 2128 96688 217648
rect 111728 2128 112048 217648
rect 127088 2128 127408 217648
rect 142448 2128 142768 217648
rect 157808 2128 158128 217648
rect 173168 2128 173488 217648
rect 188528 2128 188848 217648
rect 203888 2128 204208 217648
<< obsm4 >>
rect 2083 2483 4128 217293
rect 4608 2483 19488 217293
rect 19968 2483 34848 217293
rect 35328 2483 50208 217293
rect 50688 2483 65568 217293
rect 66048 2483 80928 217293
rect 81408 2483 96288 217293
rect 96768 2483 111648 217293
rect 112128 2483 127008 217293
rect 127488 2483 142368 217293
rect 142848 2483 157728 217293
rect 158208 2483 173088 217293
rect 173568 2483 188448 217293
rect 188928 2483 203808 217293
rect 204288 2483 217797 217293
<< labels >>
rlabel metal2 s 5446 0 5502 800 6 clock
port 1 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 io_dbus_addr[0]
port 2 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 io_dbus_addr[10]
port 3 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 io_dbus_addr[11]
port 4 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 io_dbus_addr[12]
port 5 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 io_dbus_addr[13]
port 6 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 io_dbus_addr[14]
port 7 nsew signal input
rlabel metal3 s 0 62160 800 62280 6 io_dbus_addr[15]
port 8 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 io_dbus_addr[16]
port 9 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 io_dbus_addr[17]
port 10 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 io_dbus_addr[18]
port 11 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 io_dbus_addr[19]
port 12 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 io_dbus_addr[1]
port 13 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 io_dbus_addr[20]
port 14 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 io_dbus_addr[21]
port 15 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 io_dbus_addr[22]
port 16 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 io_dbus_addr[23]
port 17 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 io_dbus_addr[24]
port 18 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 io_dbus_addr[25]
port 19 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 io_dbus_addr[26]
port 20 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 io_dbus_addr[27]
port 21 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 io_dbus_addr[28]
port 22 nsew signal input
rlabel metal3 s 0 111120 800 111240 6 io_dbus_addr[29]
port 23 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 io_dbus_addr[2]
port 24 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 io_dbus_addr[30]
port 25 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 io_dbus_addr[31]
port 26 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 io_dbus_addr[3]
port 27 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 io_dbus_addr[4]
port 28 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 io_dbus_addr[5]
port 29 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 io_dbus_addr[6]
port 30 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 io_dbus_addr[7]
port 31 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 io_dbus_addr[8]
port 32 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 io_dbus_addr[9]
port 33 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 io_dbus_ld_type[0]
port 34 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 io_dbus_ld_type[1]
port 35 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 io_dbus_ld_type[2]
port 36 nsew signal input
rlabel metal3 s 0 552 800 672 6 io_dbus_rd_en
port 37 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 io_dbus_rdata[0]
port 38 nsew signal output
rlabel metal3 s 0 45840 800 45960 6 io_dbus_rdata[10]
port 39 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 io_dbus_rdata[11]
port 40 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 io_dbus_rdata[12]
port 41 nsew signal output
rlabel metal3 s 0 56312 800 56432 6 io_dbus_rdata[13]
port 42 nsew signal output
rlabel metal3 s 0 59848 800 59968 6 io_dbus_rdata[14]
port 43 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 io_dbus_rdata[15]
port 44 nsew signal output
rlabel metal3 s 0 66784 800 66904 6 io_dbus_rdata[16]
port 45 nsew signal output
rlabel metal3 s 0 70320 800 70440 6 io_dbus_rdata[17]
port 46 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 io_dbus_rdata[18]
port 47 nsew signal output
rlabel metal3 s 0 77392 800 77512 6 io_dbus_rdata[19]
port 48 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 io_dbus_rdata[1]
port 49 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 io_dbus_rdata[20]
port 50 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 io_dbus_rdata[21]
port 51 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 io_dbus_rdata[22]
port 52 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 io_dbus_rdata[23]
port 53 nsew signal output
rlabel metal3 s 0 94800 800 94920 6 io_dbus_rdata[24]
port 54 nsew signal output
rlabel metal3 s 0 98336 800 98456 6 io_dbus_rdata[25]
port 55 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 io_dbus_rdata[26]
port 56 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 io_dbus_rdata[27]
port 57 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 io_dbus_rdata[28]
port 58 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 io_dbus_rdata[29]
port 59 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 io_dbus_rdata[2]
port 60 nsew signal output
rlabel metal3 s 0 115744 800 115864 6 io_dbus_rdata[30]
port 61 nsew signal output
rlabel metal3 s 0 119280 800 119400 6 io_dbus_rdata[31]
port 62 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 io_dbus_rdata[3]
port 63 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 io_dbus_rdata[4]
port 64 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 io_dbus_rdata[5]
port 65 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_dbus_rdata[6]
port 66 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_dbus_rdata[7]
port 67 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 io_dbus_rdata[8]
port 68 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 io_dbus_rdata[9]
port 69 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 io_dbus_st_type[0]
port 70 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 io_dbus_st_type[1]
port 71 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 io_dbus_valid
port 72 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 io_dbus_wdata[0]
port 73 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 io_dbus_wdata[10]
port 74 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 io_dbus_wdata[11]
port 75 nsew signal input
rlabel metal3 s 0 54000 800 54120 6 io_dbus_wdata[12]
port 76 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 io_dbus_wdata[13]
port 77 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 io_dbus_wdata[14]
port 78 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 io_dbus_wdata[15]
port 79 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 io_dbus_wdata[16]
port 80 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 io_dbus_wdata[17]
port 81 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 io_dbus_wdata[18]
port 82 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 io_dbus_wdata[19]
port 83 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 io_dbus_wdata[1]
port 84 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 io_dbus_wdata[20]
port 85 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 io_dbus_wdata[21]
port 86 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 io_dbus_wdata[22]
port 87 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 io_dbus_wdata[23]
port 88 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 io_dbus_wdata[24]
port 89 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 io_dbus_wdata[25]
port 90 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 io_dbus_wdata[26]
port 91 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 io_dbus_wdata[27]
port 92 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 io_dbus_wdata[28]
port 93 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 io_dbus_wdata[29]
port 94 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 io_dbus_wdata[2]
port 95 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 io_dbus_wdata[30]
port 96 nsew signal input
rlabel metal3 s 0 120368 800 120488 6 io_dbus_wdata[31]
port 97 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 io_dbus_wdata[3]
port 98 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 io_dbus_wdata[4]
port 99 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 io_dbus_wdata[5]
port 100 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 io_dbus_wdata[6]
port 101 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 io_dbus_wdata[7]
port 102 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 io_dbus_wdata[8]
port 103 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 io_dbus_wdata[9]
port 104 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 io_dbus_wr_en
port 105 nsew signal input
rlabel metal2 s 5722 219200 5778 220000 6 io_dmem_io_addr[0]
port 106 nsew signal output
rlabel metal2 s 15014 219200 15070 220000 6 io_dmem_io_addr[1]
port 107 nsew signal output
rlabel metal2 s 24214 219200 24270 220000 6 io_dmem_io_addr[2]
port 108 nsew signal output
rlabel metal2 s 33506 219200 33562 220000 6 io_dmem_io_addr[3]
port 109 nsew signal output
rlabel metal2 s 42798 219200 42854 220000 6 io_dmem_io_addr[4]
port 110 nsew signal output
rlabel metal2 s 49698 219200 49754 220000 6 io_dmem_io_addr[5]
port 111 nsew signal output
rlabel metal2 s 56690 219200 56746 220000 6 io_dmem_io_addr[6]
port 112 nsew signal output
rlabel metal2 s 63590 219200 63646 220000 6 io_dmem_io_addr[7]
port 113 nsew signal output
rlabel metal2 s 1122 219200 1178 220000 6 io_dmem_io_cs
port 114 nsew signal output
rlabel metal2 s 8022 219200 8078 220000 6 io_dmem_io_rdata[0]
port 115 nsew signal input
rlabel metal2 s 79782 219200 79838 220000 6 io_dmem_io_rdata[10]
port 116 nsew signal input
rlabel metal2 s 84474 219200 84530 220000 6 io_dmem_io_rdata[11]
port 117 nsew signal input
rlabel metal2 s 89074 219200 89130 220000 6 io_dmem_io_rdata[12]
port 118 nsew signal input
rlabel metal2 s 93674 219200 93730 220000 6 io_dmem_io_rdata[13]
port 119 nsew signal input
rlabel metal2 s 98366 219200 98422 220000 6 io_dmem_io_rdata[14]
port 120 nsew signal input
rlabel metal2 s 102966 219200 103022 220000 6 io_dmem_io_rdata[15]
port 121 nsew signal input
rlabel metal2 s 107566 219200 107622 220000 6 io_dmem_io_rdata[16]
port 122 nsew signal input
rlabel metal2 s 112258 219200 112314 220000 6 io_dmem_io_rdata[17]
port 123 nsew signal input
rlabel metal2 s 116858 219200 116914 220000 6 io_dmem_io_rdata[18]
port 124 nsew signal input
rlabel metal2 s 121458 219200 121514 220000 6 io_dmem_io_rdata[19]
port 125 nsew signal input
rlabel metal2 s 17314 219200 17370 220000 6 io_dmem_io_rdata[1]
port 126 nsew signal input
rlabel metal2 s 126150 219200 126206 220000 6 io_dmem_io_rdata[20]
port 127 nsew signal input
rlabel metal2 s 130750 219200 130806 220000 6 io_dmem_io_rdata[21]
port 128 nsew signal input
rlabel metal2 s 135350 219200 135406 220000 6 io_dmem_io_rdata[22]
port 129 nsew signal input
rlabel metal2 s 140042 219200 140098 220000 6 io_dmem_io_rdata[23]
port 130 nsew signal input
rlabel metal2 s 144642 219200 144698 220000 6 io_dmem_io_rdata[24]
port 131 nsew signal input
rlabel metal2 s 149242 219200 149298 220000 6 io_dmem_io_rdata[25]
port 132 nsew signal input
rlabel metal2 s 153934 219200 153990 220000 6 io_dmem_io_rdata[26]
port 133 nsew signal input
rlabel metal2 s 158534 219200 158590 220000 6 io_dmem_io_rdata[27]
port 134 nsew signal input
rlabel metal2 s 163134 219200 163190 220000 6 io_dmem_io_rdata[28]
port 135 nsew signal input
rlabel metal2 s 167826 219200 167882 220000 6 io_dmem_io_rdata[29]
port 136 nsew signal input
rlabel metal2 s 26514 219200 26570 220000 6 io_dmem_io_rdata[2]
port 137 nsew signal input
rlabel metal2 s 172426 219200 172482 220000 6 io_dmem_io_rdata[30]
port 138 nsew signal input
rlabel metal2 s 177026 219200 177082 220000 6 io_dmem_io_rdata[31]
port 139 nsew signal input
rlabel metal2 s 35806 219200 35862 220000 6 io_dmem_io_rdata[3]
port 140 nsew signal input
rlabel metal2 s 45098 219200 45154 220000 6 io_dmem_io_rdata[4]
port 141 nsew signal input
rlabel metal2 s 51998 219200 52054 220000 6 io_dmem_io_rdata[5]
port 142 nsew signal input
rlabel metal2 s 58990 219200 59046 220000 6 io_dmem_io_rdata[6]
port 143 nsew signal input
rlabel metal2 s 65890 219200 65946 220000 6 io_dmem_io_rdata[7]
port 144 nsew signal input
rlabel metal2 s 70582 219200 70638 220000 6 io_dmem_io_rdata[8]
port 145 nsew signal input
rlabel metal2 s 75182 219200 75238 220000 6 io_dmem_io_rdata[9]
port 146 nsew signal input
rlabel metal2 s 10322 219200 10378 220000 6 io_dmem_io_st_type[0]
port 147 nsew signal output
rlabel metal2 s 19614 219200 19670 220000 6 io_dmem_io_st_type[1]
port 148 nsew signal output
rlabel metal2 s 28906 219200 28962 220000 6 io_dmem_io_st_type[2]
port 149 nsew signal output
rlabel metal2 s 38106 219200 38162 220000 6 io_dmem_io_st_type[3]
port 150 nsew signal output
rlabel metal2 s 12622 219200 12678 220000 6 io_dmem_io_wdata[0]
port 151 nsew signal output
rlabel metal2 s 82082 219200 82138 220000 6 io_dmem_io_wdata[10]
port 152 nsew signal output
rlabel metal2 s 86774 219200 86830 220000 6 io_dmem_io_wdata[11]
port 153 nsew signal output
rlabel metal2 s 91374 219200 91430 220000 6 io_dmem_io_wdata[12]
port 154 nsew signal output
rlabel metal2 s 95974 219200 96030 220000 6 io_dmem_io_wdata[13]
port 155 nsew signal output
rlabel metal2 s 100666 219200 100722 220000 6 io_dmem_io_wdata[14]
port 156 nsew signal output
rlabel metal2 s 105266 219200 105322 220000 6 io_dmem_io_wdata[15]
port 157 nsew signal output
rlabel metal2 s 109866 219200 109922 220000 6 io_dmem_io_wdata[16]
port 158 nsew signal output
rlabel metal2 s 114558 219200 114614 220000 6 io_dmem_io_wdata[17]
port 159 nsew signal output
rlabel metal2 s 119158 219200 119214 220000 6 io_dmem_io_wdata[18]
port 160 nsew signal output
rlabel metal2 s 123758 219200 123814 220000 6 io_dmem_io_wdata[19]
port 161 nsew signal output
rlabel metal2 s 21914 219200 21970 220000 6 io_dmem_io_wdata[1]
port 162 nsew signal output
rlabel metal2 s 128450 219200 128506 220000 6 io_dmem_io_wdata[20]
port 163 nsew signal output
rlabel metal2 s 133050 219200 133106 220000 6 io_dmem_io_wdata[21]
port 164 nsew signal output
rlabel metal2 s 137650 219200 137706 220000 6 io_dmem_io_wdata[22]
port 165 nsew signal output
rlabel metal2 s 142342 219200 142398 220000 6 io_dmem_io_wdata[23]
port 166 nsew signal output
rlabel metal2 s 146942 219200 146998 220000 6 io_dmem_io_wdata[24]
port 167 nsew signal output
rlabel metal2 s 151542 219200 151598 220000 6 io_dmem_io_wdata[25]
port 168 nsew signal output
rlabel metal2 s 156234 219200 156290 220000 6 io_dmem_io_wdata[26]
port 169 nsew signal output
rlabel metal2 s 160834 219200 160890 220000 6 io_dmem_io_wdata[27]
port 170 nsew signal output
rlabel metal2 s 165434 219200 165490 220000 6 io_dmem_io_wdata[28]
port 171 nsew signal output
rlabel metal2 s 170126 219200 170182 220000 6 io_dmem_io_wdata[29]
port 172 nsew signal output
rlabel metal2 s 31206 219200 31262 220000 6 io_dmem_io_wdata[2]
port 173 nsew signal output
rlabel metal2 s 174726 219200 174782 220000 6 io_dmem_io_wdata[30]
port 174 nsew signal output
rlabel metal2 s 179326 219200 179382 220000 6 io_dmem_io_wdata[31]
port 175 nsew signal output
rlabel metal2 s 40406 219200 40462 220000 6 io_dmem_io_wdata[3]
port 176 nsew signal output
rlabel metal2 s 47398 219200 47454 220000 6 io_dmem_io_wdata[4]
port 177 nsew signal output
rlabel metal2 s 54298 219200 54354 220000 6 io_dmem_io_wdata[5]
port 178 nsew signal output
rlabel metal2 s 61290 219200 61346 220000 6 io_dmem_io_wdata[6]
port 179 nsew signal output
rlabel metal2 s 68190 219200 68246 220000 6 io_dmem_io_wdata[7]
port 180 nsew signal output
rlabel metal2 s 72882 219200 72938 220000 6 io_dmem_io_wdata[8]
port 181 nsew signal output
rlabel metal2 s 77482 219200 77538 220000 6 io_dmem_io_wdata[9]
port 182 nsew signal output
rlabel metal2 s 3422 219200 3478 220000 6 io_dmem_io_wr_en
port 183 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 io_ibus_addr[0]
port 184 nsew signal input
rlabel metal3 s 0 146072 800 146192 6 io_ibus_addr[10]
port 185 nsew signal input
rlabel metal3 s 0 148384 800 148504 6 io_ibus_addr[11]
port 186 nsew signal input
rlabel metal3 s 0 150696 800 150816 6 io_ibus_addr[12]
port 187 nsew signal input
rlabel metal3 s 0 153008 800 153128 6 io_ibus_addr[13]
port 188 nsew signal input
rlabel metal3 s 0 155320 800 155440 6 io_ibus_addr[14]
port 189 nsew signal input
rlabel metal3 s 0 157632 800 157752 6 io_ibus_addr[15]
port 190 nsew signal input
rlabel metal3 s 0 159944 800 160064 6 io_ibus_addr[16]
port 191 nsew signal input
rlabel metal3 s 0 162256 800 162376 6 io_ibus_addr[17]
port 192 nsew signal input
rlabel metal3 s 0 164704 800 164824 6 io_ibus_addr[18]
port 193 nsew signal input
rlabel metal3 s 0 167016 800 167136 6 io_ibus_addr[19]
port 194 nsew signal input
rlabel metal3 s 0 125128 800 125248 6 io_ibus_addr[1]
port 195 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 io_ibus_addr[20]
port 196 nsew signal input
rlabel metal3 s 0 171640 800 171760 6 io_ibus_addr[21]
port 197 nsew signal input
rlabel metal3 s 0 173952 800 174072 6 io_ibus_addr[22]
port 198 nsew signal input
rlabel metal3 s 0 176264 800 176384 6 io_ibus_addr[23]
port 199 nsew signal input
rlabel metal3 s 0 178576 800 178696 6 io_ibus_addr[24]
port 200 nsew signal input
rlabel metal3 s 0 180888 800 181008 6 io_ibus_addr[25]
port 201 nsew signal input
rlabel metal3 s 0 183336 800 183456 6 io_ibus_addr[26]
port 202 nsew signal input
rlabel metal3 s 0 185648 800 185768 6 io_ibus_addr[27]
port 203 nsew signal input
rlabel metal3 s 0 187960 800 188080 6 io_ibus_addr[28]
port 204 nsew signal input
rlabel metal3 s 0 190272 800 190392 6 io_ibus_addr[29]
port 205 nsew signal input
rlabel metal3 s 0 127440 800 127560 6 io_ibus_addr[2]
port 206 nsew signal input
rlabel metal3 s 0 192584 800 192704 6 io_ibus_addr[30]
port 207 nsew signal input
rlabel metal3 s 0 194896 800 195016 6 io_ibus_addr[31]
port 208 nsew signal input
rlabel metal3 s 0 129752 800 129872 6 io_ibus_addr[3]
port 209 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 io_ibus_addr[4]
port 210 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 io_ibus_addr[5]
port 211 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 io_ibus_addr[6]
port 212 nsew signal input
rlabel metal3 s 0 139000 800 139120 6 io_ibus_addr[7]
port 213 nsew signal input
rlabel metal3 s 0 141312 800 141432 6 io_ibus_addr[8]
port 214 nsew signal input
rlabel metal3 s 0 143624 800 143744 6 io_ibus_addr[9]
port 215 nsew signal input
rlabel metal3 s 0 123904 800 124024 6 io_ibus_inst[0]
port 216 nsew signal output
rlabel metal3 s 0 147160 800 147280 6 io_ibus_inst[10]
port 217 nsew signal output
rlabel metal3 s 0 149472 800 149592 6 io_ibus_inst[11]
port 218 nsew signal output
rlabel metal3 s 0 151784 800 151904 6 io_ibus_inst[12]
port 219 nsew signal output
rlabel metal3 s 0 154232 800 154352 6 io_ibus_inst[13]
port 220 nsew signal output
rlabel metal3 s 0 156544 800 156664 6 io_ibus_inst[14]
port 221 nsew signal output
rlabel metal3 s 0 158856 800 158976 6 io_ibus_inst[15]
port 222 nsew signal output
rlabel metal3 s 0 161168 800 161288 6 io_ibus_inst[16]
port 223 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 io_ibus_inst[17]
port 224 nsew signal output
rlabel metal3 s 0 165792 800 165912 6 io_ibus_inst[18]
port 225 nsew signal output
rlabel metal3 s 0 168104 800 168224 6 io_ibus_inst[19]
port 226 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 io_ibus_inst[1]
port 227 nsew signal output
rlabel metal3 s 0 170416 800 170536 6 io_ibus_inst[20]
port 228 nsew signal output
rlabel metal3 s 0 172864 800 172984 6 io_ibus_inst[21]
port 229 nsew signal output
rlabel metal3 s 0 175176 800 175296 6 io_ibus_inst[22]
port 230 nsew signal output
rlabel metal3 s 0 177488 800 177608 6 io_ibus_inst[23]
port 231 nsew signal output
rlabel metal3 s 0 179800 800 179920 6 io_ibus_inst[24]
port 232 nsew signal output
rlabel metal3 s 0 182112 800 182232 6 io_ibus_inst[25]
port 233 nsew signal output
rlabel metal3 s 0 184424 800 184544 6 io_ibus_inst[26]
port 234 nsew signal output
rlabel metal3 s 0 186736 800 186856 6 io_ibus_inst[27]
port 235 nsew signal output
rlabel metal3 s 0 189048 800 189168 6 io_ibus_inst[28]
port 236 nsew signal output
rlabel metal3 s 0 191360 800 191480 6 io_ibus_inst[29]
port 237 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 io_ibus_inst[2]
port 238 nsew signal output
rlabel metal3 s 0 193808 800 193928 6 io_ibus_inst[30]
port 239 nsew signal output
rlabel metal3 s 0 196120 800 196240 6 io_ibus_inst[31]
port 240 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 io_ibus_inst[3]
port 241 nsew signal output
rlabel metal3 s 0 133152 800 133272 6 io_ibus_inst[4]
port 242 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 io_ibus_inst[5]
port 243 nsew signal output
rlabel metal3 s 0 137912 800 138032 6 io_ibus_inst[6]
port 244 nsew signal output
rlabel metal3 s 0 140224 800 140344 6 io_ibus_inst[7]
port 245 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 io_ibus_inst[8]
port 246 nsew signal output
rlabel metal3 s 0 144848 800 144968 6 io_ibus_inst[9]
port 247 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 io_ibus_valid
port 248 nsew signal output
rlabel metal3 s 219200 175312 220000 175432 6 io_imem_io_addr[0]
port 249 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 io_imem_io_addr[1]
port 250 nsew signal output
rlabel metal2 s 184018 219200 184074 220000 6 io_imem_io_addr[2]
port 251 nsew signal output
rlabel metal3 s 0 201968 800 202088 6 io_imem_io_addr[3]
port 252 nsew signal output
rlabel metal3 s 219200 179120 220000 179240 6 io_imem_io_addr[4]
port 253 nsew signal output
rlabel metal3 s 219200 182928 220000 183048 6 io_imem_io_addr[5]
port 254 nsew signal output
rlabel metal3 s 219200 186600 220000 186720 6 io_imem_io_addr[6]
port 255 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 io_imem_io_addr[7]
port 256 nsew signal output
rlabel metal2 s 115386 0 115442 800 6 io_imem_io_addr[8]
port 257 nsew signal output
rlabel metal2 s 181718 219200 181774 220000 6 io_imem_io_cs
port 258 nsew signal output
rlabel metal2 s 60370 0 60426 800 6 io_imem_io_rdata[0]
port 259 nsew signal input
rlabel metal3 s 219200 194216 220000 194336 6 io_imem_io_rdata[10]
port 260 nsew signal input
rlabel metal3 s 219200 196120 220000 196240 6 io_imem_io_rdata[11]
port 261 nsew signal input
rlabel metal3 s 219200 198024 220000 198144 6 io_imem_io_rdata[12]
port 262 nsew signal input
rlabel metal3 s 0 208904 800 209024 6 io_imem_io_rdata[13]
port 263 nsew signal input
rlabel metal3 s 0 209992 800 210112 6 io_imem_io_rdata[14]
port 264 nsew signal input
rlabel metal3 s 219200 201832 220000 201952 6 io_imem_io_rdata[15]
port 265 nsew signal input
rlabel metal2 s 137374 0 137430 800 6 io_imem_io_rdata[16]
port 266 nsew signal input
rlabel metal3 s 219200 203736 220000 203856 6 io_imem_io_rdata[17]
port 267 nsew signal input
rlabel metal3 s 0 212440 800 212560 6 io_imem_io_rdata[18]
port 268 nsew signal input
rlabel metal3 s 0 213528 800 213648 6 io_imem_io_rdata[19]
port 269 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 io_imem_io_rdata[1]
port 270 nsew signal input
rlabel metal3 s 0 214752 800 214872 6 io_imem_io_rdata[20]
port 271 nsew signal input
rlabel metal2 s 204810 219200 204866 220000 6 io_imem_io_rdata[21]
port 272 nsew signal input
rlabel metal3 s 0 217064 800 217184 6 io_imem_io_rdata[22]
port 273 nsew signal input
rlabel metal3 s 0 218152 800 218272 6 io_imem_io_rdata[23]
port 274 nsew signal input
rlabel metal2 s 207110 219200 207166 220000 6 io_imem_io_rdata[24]
port 275 nsew signal input
rlabel metal2 s 192390 0 192446 800 6 io_imem_io_rdata[25]
port 276 nsew signal input
rlabel metal3 s 219200 211352 220000 211472 6 io_imem_io_rdata[26]
port 277 nsew signal input
rlabel metal2 s 203338 0 203394 800 6 io_imem_io_rdata[27]
port 278 nsew signal input
rlabel metal2 s 211802 219200 211858 220000 6 io_imem_io_rdata[28]
port 279 nsew signal input
rlabel metal3 s 0 219376 800 219496 6 io_imem_io_rdata[29]
port 280 nsew signal input
rlabel metal2 s 186318 219200 186374 220000 6 io_imem_io_rdata[2]
port 281 nsew signal input
rlabel metal2 s 214102 219200 214158 220000 6 io_imem_io_rdata[30]
port 282 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 io_imem_io_rdata[31]
port 283 nsew signal input
rlabel metal3 s 219200 177216 220000 177336 6 io_imem_io_rdata[3]
port 284 nsew signal input
rlabel metal3 s 219200 181024 220000 181144 6 io_imem_io_rdata[4]
port 285 nsew signal input
rlabel metal3 s 219200 184696 220000 184816 6 io_imem_io_rdata[5]
port 286 nsew signal input
rlabel metal3 s 0 203056 800 203176 6 io_imem_io_rdata[6]
port 287 nsew signal input
rlabel metal3 s 0 204280 800 204400 6 io_imem_io_rdata[7]
port 288 nsew signal input
rlabel metal2 s 197910 219200 197966 220000 6 io_imem_io_rdata[8]
port 289 nsew signal input
rlabel metal3 s 0 205368 800 205488 6 io_imem_io_rdata[9]
port 290 nsew signal input
rlabel metal3 s 0 199520 800 199640 6 io_imem_io_wdata[0]
port 291 nsew signal output
rlabel metal3 s 0 206592 800 206712 6 io_imem_io_wdata[10]
port 292 nsew signal output
rlabel metal2 s 200210 219200 200266 220000 6 io_imem_io_wdata[11]
port 293 nsew signal output
rlabel metal3 s 0 207680 800 207800 6 io_imem_io_wdata[12]
port 294 nsew signal output
rlabel metal3 s 219200 199928 220000 200048 6 io_imem_io_wdata[13]
port 295 nsew signal output
rlabel metal3 s 0 211216 800 211336 6 io_imem_io_wdata[14]
port 296 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 io_imem_io_wdata[15]
port 297 nsew signal output
rlabel metal2 s 202510 219200 202566 220000 6 io_imem_io_wdata[16]
port 298 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 io_imem_io_wdata[17]
port 299 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 io_imem_io_wdata[18]
port 300 nsew signal output
rlabel metal2 s 170402 0 170458 800 6 io_imem_io_wdata[19]
port 301 nsew signal output
rlabel metal3 s 0 200744 800 200864 6 io_imem_io_wdata[1]
port 302 nsew signal output
rlabel metal3 s 0 215840 800 215960 6 io_imem_io_wdata[20]
port 303 nsew signal output
rlabel metal3 s 219200 205640 220000 205760 6 io_imem_io_wdata[21]
port 304 nsew signal output
rlabel metal2 s 181350 0 181406 800 6 io_imem_io_wdata[22]
port 305 nsew signal output
rlabel metal3 s 219200 207544 220000 207664 6 io_imem_io_wdata[23]
port 306 nsew signal output
rlabel metal2 s 209502 219200 209558 220000 6 io_imem_io_wdata[24]
port 307 nsew signal output
rlabel metal3 s 219200 209448 220000 209568 6 io_imem_io_wdata[25]
port 308 nsew signal output
rlabel metal3 s 219200 213256 220000 213376 6 io_imem_io_wdata[26]
port 309 nsew signal output
rlabel metal3 s 219200 215160 220000 215280 6 io_imem_io_wdata[27]
port 310 nsew signal output
rlabel metal3 s 219200 217064 220000 217184 6 io_imem_io_wdata[28]
port 311 nsew signal output
rlabel metal3 s 219200 218968 220000 219088 6 io_imem_io_wdata[29]
port 312 nsew signal output
rlabel metal2 s 188618 219200 188674 220000 6 io_imem_io_wdata[2]
port 313 nsew signal output
rlabel metal2 s 216402 219200 216458 220000 6 io_imem_io_wdata[30]
port 314 nsew signal output
rlabel metal2 s 218702 219200 218758 220000 6 io_imem_io_wdata[31]
port 315 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 io_imem_io_wdata[3]
port 316 nsew signal output
rlabel metal2 s 190918 219200 190974 220000 6 io_imem_io_wdata[4]
port 317 nsew signal output
rlabel metal2 s 193218 219200 193274 220000 6 io_imem_io_wdata[5]
port 318 nsew signal output
rlabel metal3 s 219200 188504 220000 188624 6 io_imem_io_wdata[6]
port 319 nsew signal output
rlabel metal2 s 195610 219200 195666 220000 6 io_imem_io_wdata[7]
port 320 nsew signal output
rlabel metal3 s 219200 190408 220000 190528 6 io_imem_io_wdata[8]
port 321 nsew signal output
rlabel metal3 s 219200 192312 220000 192432 6 io_imem_io_wdata[9]
port 322 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 io_imem_io_wr_en
port 323 nsew signal output
rlabel metal3 s 219200 824 220000 944 6 io_motor_ack_i
port 324 nsew signal input
rlabel metal3 s 219200 2592 220000 2712 6 io_motor_addr_sel
port 325 nsew signal output
rlabel metal3 s 219200 4496 220000 4616 6 io_motor_data_i[0]
port 326 nsew signal input
rlabel metal3 s 219200 23536 220000 23656 6 io_motor_data_i[10]
port 327 nsew signal input
rlabel metal3 s 219200 25440 220000 25560 6 io_motor_data_i[11]
port 328 nsew signal input
rlabel metal3 s 219200 27344 220000 27464 6 io_motor_data_i[12]
port 329 nsew signal input
rlabel metal3 s 219200 29248 220000 29368 6 io_motor_data_i[13]
port 330 nsew signal input
rlabel metal3 s 219200 31152 220000 31272 6 io_motor_data_i[14]
port 331 nsew signal input
rlabel metal3 s 219200 33056 220000 33176 6 io_motor_data_i[15]
port 332 nsew signal input
rlabel metal3 s 219200 34960 220000 35080 6 io_motor_data_i[16]
port 333 nsew signal input
rlabel metal3 s 219200 36864 220000 36984 6 io_motor_data_i[17]
port 334 nsew signal input
rlabel metal3 s 219200 38632 220000 38752 6 io_motor_data_i[18]
port 335 nsew signal input
rlabel metal3 s 219200 40536 220000 40656 6 io_motor_data_i[19]
port 336 nsew signal input
rlabel metal3 s 219200 6400 220000 6520 6 io_motor_data_i[1]
port 337 nsew signal input
rlabel metal3 s 219200 42440 220000 42560 6 io_motor_data_i[20]
port 338 nsew signal input
rlabel metal3 s 219200 44344 220000 44464 6 io_motor_data_i[21]
port 339 nsew signal input
rlabel metal3 s 219200 46248 220000 46368 6 io_motor_data_i[22]
port 340 nsew signal input
rlabel metal3 s 219200 48152 220000 48272 6 io_motor_data_i[23]
port 341 nsew signal input
rlabel metal3 s 219200 50056 220000 50176 6 io_motor_data_i[24]
port 342 nsew signal input
rlabel metal3 s 219200 51960 220000 52080 6 io_motor_data_i[25]
port 343 nsew signal input
rlabel metal3 s 219200 53864 220000 53984 6 io_motor_data_i[26]
port 344 nsew signal input
rlabel metal3 s 219200 55768 220000 55888 6 io_motor_data_i[27]
port 345 nsew signal input
rlabel metal3 s 219200 57672 220000 57792 6 io_motor_data_i[28]
port 346 nsew signal input
rlabel metal3 s 219200 59576 220000 59696 6 io_motor_data_i[29]
port 347 nsew signal input
rlabel metal3 s 219200 8304 220000 8424 6 io_motor_data_i[2]
port 348 nsew signal input
rlabel metal3 s 219200 61480 220000 61600 6 io_motor_data_i[30]
port 349 nsew signal input
rlabel metal3 s 219200 63384 220000 63504 6 io_motor_data_i[31]
port 350 nsew signal input
rlabel metal3 s 219200 10208 220000 10328 6 io_motor_data_i[3]
port 351 nsew signal input
rlabel metal3 s 219200 12112 220000 12232 6 io_motor_data_i[4]
port 352 nsew signal input
rlabel metal3 s 219200 14016 220000 14136 6 io_motor_data_i[5]
port 353 nsew signal input
rlabel metal3 s 219200 15920 220000 16040 6 io_motor_data_i[6]
port 354 nsew signal input
rlabel metal3 s 219200 17824 220000 17944 6 io_motor_data_i[7]
port 355 nsew signal input
rlabel metal3 s 219200 19728 220000 19848 6 io_motor_data_i[8]
port 356 nsew signal input
rlabel metal3 s 219200 21632 220000 21752 6 io_motor_data_i[9]
port 357 nsew signal input
rlabel metal3 s 219200 167696 220000 167816 6 io_spi_clk
port 358 nsew signal output
rlabel metal3 s 219200 169600 220000 169720 6 io_spi_cs
port 359 nsew signal output
rlabel metal3 s 0 197208 800 197328 6 io_spi_irq
port 360 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 io_spi_miso
port 361 nsew signal input
rlabel metal3 s 219200 171504 220000 171624 6 io_spi_mosi
port 362 nsew signal output
rlabel metal3 s 0 198432 800 198552 6 io_uart_irq
port 363 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 io_uart_rx
port 364 nsew signal input
rlabel metal3 s 219200 173408 220000 173528 6 io_uart_tx
port 365 nsew signal output
rlabel metal3 s 219200 69096 220000 69216 6 io_wbm_m2s_addr[0]
port 366 nsew signal output
rlabel metal3 s 219200 114520 220000 114640 6 io_wbm_m2s_addr[10]
port 367 nsew signal output
rlabel metal3 s 219200 118328 220000 118448 6 io_wbm_m2s_addr[11]
port 368 nsew signal output
rlabel metal3 s 219200 122136 220000 122256 6 io_wbm_m2s_addr[12]
port 369 nsew signal output
rlabel metal3 s 219200 125944 220000 126064 6 io_wbm_m2s_addr[13]
port 370 nsew signal output
rlabel metal3 s 219200 129752 220000 129872 6 io_wbm_m2s_addr[14]
port 371 nsew signal output
rlabel metal3 s 219200 133560 220000 133680 6 io_wbm_m2s_addr[15]
port 372 nsew signal output
rlabel metal3 s 219200 74672 220000 74792 6 io_wbm_m2s_addr[1]
port 373 nsew signal output
rlabel metal3 s 219200 80384 220000 80504 6 io_wbm_m2s_addr[2]
port 374 nsew signal output
rlabel metal3 s 219200 86096 220000 86216 6 io_wbm_m2s_addr[3]
port 375 nsew signal output
rlabel metal3 s 219200 91808 220000 91928 6 io_wbm_m2s_addr[4]
port 376 nsew signal output
rlabel metal3 s 219200 95616 220000 95736 6 io_wbm_m2s_addr[5]
port 377 nsew signal output
rlabel metal3 s 219200 99424 220000 99544 6 io_wbm_m2s_addr[6]
port 378 nsew signal output
rlabel metal3 s 219200 103232 220000 103352 6 io_wbm_m2s_addr[7]
port 379 nsew signal output
rlabel metal3 s 219200 107040 220000 107160 6 io_wbm_m2s_addr[8]
port 380 nsew signal output
rlabel metal3 s 219200 110848 220000 110968 6 io_wbm_m2s_addr[9]
port 381 nsew signal output
rlabel metal3 s 219200 71000 220000 71120 6 io_wbm_m2s_data[0]
port 382 nsew signal output
rlabel metal3 s 219200 116424 220000 116544 6 io_wbm_m2s_data[10]
port 383 nsew signal output
rlabel metal3 s 219200 120232 220000 120352 6 io_wbm_m2s_data[11]
port 384 nsew signal output
rlabel metal3 s 219200 124040 220000 124160 6 io_wbm_m2s_data[12]
port 385 nsew signal output
rlabel metal3 s 219200 127848 220000 127968 6 io_wbm_m2s_data[13]
port 386 nsew signal output
rlabel metal3 s 219200 131656 220000 131776 6 io_wbm_m2s_data[14]
port 387 nsew signal output
rlabel metal3 s 219200 135464 220000 135584 6 io_wbm_m2s_data[15]
port 388 nsew signal output
rlabel metal3 s 219200 137368 220000 137488 6 io_wbm_m2s_data[16]
port 389 nsew signal output
rlabel metal3 s 219200 139272 220000 139392 6 io_wbm_m2s_data[17]
port 390 nsew signal output
rlabel metal3 s 219200 141176 220000 141296 6 io_wbm_m2s_data[18]
port 391 nsew signal output
rlabel metal3 s 219200 143080 220000 143200 6 io_wbm_m2s_data[19]
port 392 nsew signal output
rlabel metal3 s 219200 76576 220000 76696 6 io_wbm_m2s_data[1]
port 393 nsew signal output
rlabel metal3 s 219200 144984 220000 145104 6 io_wbm_m2s_data[20]
port 394 nsew signal output
rlabel metal3 s 219200 146888 220000 147008 6 io_wbm_m2s_data[21]
port 395 nsew signal output
rlabel metal3 s 219200 148656 220000 148776 6 io_wbm_m2s_data[22]
port 396 nsew signal output
rlabel metal3 s 219200 150560 220000 150680 6 io_wbm_m2s_data[23]
port 397 nsew signal output
rlabel metal3 s 219200 152464 220000 152584 6 io_wbm_m2s_data[24]
port 398 nsew signal output
rlabel metal3 s 219200 154368 220000 154488 6 io_wbm_m2s_data[25]
port 399 nsew signal output
rlabel metal3 s 219200 156272 220000 156392 6 io_wbm_m2s_data[26]
port 400 nsew signal output
rlabel metal3 s 219200 158176 220000 158296 6 io_wbm_m2s_data[27]
port 401 nsew signal output
rlabel metal3 s 219200 160080 220000 160200 6 io_wbm_m2s_data[28]
port 402 nsew signal output
rlabel metal3 s 219200 161984 220000 162104 6 io_wbm_m2s_data[29]
port 403 nsew signal output
rlabel metal3 s 219200 82288 220000 82408 6 io_wbm_m2s_data[2]
port 404 nsew signal output
rlabel metal3 s 219200 163888 220000 164008 6 io_wbm_m2s_data[30]
port 405 nsew signal output
rlabel metal3 s 219200 165792 220000 165912 6 io_wbm_m2s_data[31]
port 406 nsew signal output
rlabel metal3 s 219200 88000 220000 88120 6 io_wbm_m2s_data[3]
port 407 nsew signal output
rlabel metal3 s 219200 93712 220000 93832 6 io_wbm_m2s_data[4]
port 408 nsew signal output
rlabel metal3 s 219200 97520 220000 97640 6 io_wbm_m2s_data[5]
port 409 nsew signal output
rlabel metal3 s 219200 101328 220000 101448 6 io_wbm_m2s_data[6]
port 410 nsew signal output
rlabel metal3 s 219200 105136 220000 105256 6 io_wbm_m2s_data[7]
port 411 nsew signal output
rlabel metal3 s 219200 108944 220000 109064 6 io_wbm_m2s_data[8]
port 412 nsew signal output
rlabel metal3 s 219200 112616 220000 112736 6 io_wbm_m2s_data[9]
port 413 nsew signal output
rlabel metal3 s 219200 72904 220000 73024 6 io_wbm_m2s_sel[0]
port 414 nsew signal output
rlabel metal3 s 219200 78480 220000 78600 6 io_wbm_m2s_sel[1]
port 415 nsew signal output
rlabel metal3 s 219200 84192 220000 84312 6 io_wbm_m2s_sel[2]
port 416 nsew signal output
rlabel metal3 s 219200 89904 220000 90024 6 io_wbm_m2s_sel[3]
port 417 nsew signal output
rlabel metal3 s 219200 65288 220000 65408 6 io_wbm_m2s_stb
port 418 nsew signal output
rlabel metal3 s 219200 67192 220000 67312 6 io_wbm_m2s_we
port 419 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 reset
port 420 nsew signal input
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 421 nsew power input
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 421 nsew power input
rlabel metal4 s 65648 2128 65968 217648 6 vccd1
port 421 nsew power input
rlabel metal4 s 96368 2128 96688 217648 6 vccd1
port 421 nsew power input
rlabel metal4 s 127088 2128 127408 217648 6 vccd1
port 421 nsew power input
rlabel metal4 s 157808 2128 158128 217648 6 vccd1
port 421 nsew power input
rlabel metal4 s 188528 2128 188848 217648 6 vccd1
port 421 nsew power input
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 422 nsew ground input
rlabel metal4 s 50288 2128 50608 217648 6 vssd1
port 422 nsew ground input
rlabel metal4 s 81008 2128 81328 217648 6 vssd1
port 422 nsew ground input
rlabel metal4 s 111728 2128 112048 217648 6 vssd1
port 422 nsew ground input
rlabel metal4 s 142448 2128 142768 217648 6 vssd1
port 422 nsew ground input
rlabel metal4 s 173168 2128 173488 217648 6 vssd1
port 422 nsew ground input
rlabel metal4 s 203888 2128 204208 217648 6 vssd1
port 422 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 220000 220000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18604204
string GDS_FILE /home/em/mpw/UETRV-ECORE/openlane/Wishbone_InterConnect/runs/Wishbone_InterConnect/results/finishing/WB_InterConnect.magic.gds
string GDS_START 865950
<< end >>

