VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Motor_Top
  CLASS BLOCK ;
  FOREIGN Motor_Top ;
  ORIGIN 0.000 0.000 ;
  SIZE 400.000 BY 400.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END clock
  PIN io_ba_match
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END io_ba_match
  PIN io_motor_irq
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 8.200 400.000 8.800 ;
    END
  END io_motor_irq
  PIN io_pwm_high
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 396.000 9.110 400.000 ;
    END
  END io_pwm_high
  PIN io_pwm_low
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 396.000 27.050 400.000 ;
    END
  END io_pwm_low
  PIN io_qei_ch_a
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 25.200 400.000 25.800 ;
    END
  END io_qei_ch_a
  PIN io_qei_ch_b
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END io_qei_ch_b
  PIN io_wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 42.880 400.000 43.480 ;
    END
  END io_wbs_ack_o
  PIN io_wbs_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END io_wbs_data_o[0]
  PIN io_wbs_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 396.000 190.810 400.000 ;
    END
  END io_wbs_data_o[10]
  PIN io_wbs_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 199.280 400.000 199.880 ;
    END
  END io_wbs_data_o[11]
  PIN io_wbs_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END io_wbs_data_o[12]
  PIN io_wbs_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END io_wbs_data_o[13]
  PIN io_wbs_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_wbs_data_o[14]
  PIN io_wbs_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 233.960 400.000 234.560 ;
    END
  END io_wbs_data_o[15]
  PIN io_wbs_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 396.000 227.150 400.000 ;
    END
  END io_wbs_data_o[16]
  PIN io_wbs_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END io_wbs_data_o[17]
  PIN io_wbs_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END io_wbs_data_o[18]
  PIN io_wbs_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.210 396.000 263.490 400.000 ;
    END
  END io_wbs_data_o[19]
  PIN io_wbs_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END io_wbs_data_o[1]
  PIN io_wbs_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 268.640 400.000 269.240 ;
    END
  END io_wbs_data_o[20]
  PIN io_wbs_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END io_wbs_data_o[21]
  PIN io_wbs_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 396.000 299.830 400.000 ;
    END
  END io_wbs_data_o[22]
  PIN io_wbs_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END io_wbs_data_o[23]
  PIN io_wbs_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 321.000 400.000 321.600 ;
    END
  END io_wbs_data_o[24]
  PIN io_wbs_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 396.000 336.170 400.000 ;
    END
  END io_wbs_data_o[25]
  PIN io_wbs_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END io_wbs_data_o[26]
  PIN io_wbs_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 338.000 400.000 338.600 ;
    END
  END io_wbs_data_o[27]
  PIN io_wbs_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 355.680 400.000 356.280 ;
    END
  END io_wbs_data_o[28]
  PIN io_wbs_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END io_wbs_data_o[29]
  PIN io_wbs_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 59.880 400.000 60.480 ;
    END
  END io_wbs_data_o[2]
  PIN io_wbs_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END io_wbs_data_o[30]
  PIN io_wbs_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 396.000 390.910 400.000 ;
    END
  END io_wbs_data_o[31]
  PIN io_wbs_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END io_wbs_data_o[3]
  PIN io_wbs_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END io_wbs_data_o[4]
  PIN io_wbs_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 396.000 63.390 400.000 ;
    END
  END io_wbs_data_o[5]
  PIN io_wbs_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 112.240 400.000 112.840 ;
    END
  END io_wbs_data_o[6]
  PIN io_wbs_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END io_wbs_data_o[7]
  PIN io_wbs_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END io_wbs_data_o[8]
  PIN io_wbs_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 129.240 400.000 129.840 ;
    END
  END io_wbs_data_o[9]
  PIN io_wbs_m2s_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END io_wbs_m2s_addr[0]
  PIN io_wbs_m2s_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END io_wbs_m2s_addr[10]
  PIN io_wbs_m2s_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 216.280 400.000 216.880 ;
    END
  END io_wbs_m2s_addr[11]
  PIN io_wbs_m2s_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END io_wbs_m2s_addr[12]
  PIN io_wbs_m2s_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 396.000 209.210 400.000 ;
    END
  END io_wbs_m2s_addr[13]
  PIN io_wbs_m2s_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END io_wbs_m2s_addr[14]
  PIN io_wbs_m2s_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END io_wbs_m2s_addr[15]
  PIN io_wbs_m2s_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END io_wbs_m2s_addr[1]
  PIN io_wbs_m2s_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END io_wbs_m2s_addr[2]
  PIN io_wbs_m2s_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END io_wbs_m2s_addr[3]
  PIN io_wbs_m2s_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END io_wbs_m2s_addr[4]
  PIN io_wbs_m2s_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 396.000 81.790 400.000 ;
    END
  END io_wbs_m2s_addr[5]
  PIN io_wbs_m2s_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 396.000 118.130 400.000 ;
    END
  END io_wbs_m2s_addr[6]
  PIN io_wbs_m2s_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END io_wbs_m2s_addr[7]
  PIN io_wbs_m2s_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 396.000 154.470 400.000 ;
    END
  END io_wbs_m2s_addr[8]
  PIN io_wbs_m2s_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 146.920 400.000 147.520 ;
    END
  END io_wbs_m2s_addr[9]
  PIN io_wbs_m2s_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END io_wbs_m2s_data[0]
  PIN io_wbs_m2s_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 181.600 400.000 182.200 ;
    END
  END io_wbs_m2s_data[10]
  PIN io_wbs_m2s_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END io_wbs_m2s_data[11]
  PIN io_wbs_m2s_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END io_wbs_m2s_data[12]
  PIN io_wbs_m2s_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END io_wbs_m2s_data[13]
  PIN io_wbs_m2s_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END io_wbs_m2s_data[14]
  PIN io_wbs_m2s_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 0.000 275.450 4.000 ;
    END
  END io_wbs_m2s_data[15]
  PIN io_wbs_m2s_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.880 4.000 315.480 ;
    END
  END io_wbs_m2s_data[16]
  PIN io_wbs_m2s_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 396.000 245.550 400.000 ;
    END
  END io_wbs_m2s_data[17]
  PIN io_wbs_m2s_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 250.960 400.000 251.560 ;
    END
  END io_wbs_m2s_data[18]
  PIN io_wbs_m2s_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 396.000 281.890 400.000 ;
    END
  END io_wbs_m2s_data[19]
  PIN io_wbs_m2s_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END io_wbs_m2s_data[1]
  PIN io_wbs_m2s_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 286.320 400.000 286.920 ;
    END
  END io_wbs_m2s_data[20]
  PIN io_wbs_m2s_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END io_wbs_m2s_data[21]
  PIN io_wbs_m2s_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 396.000 318.230 400.000 ;
    END
  END io_wbs_m2s_data[22]
  PIN io_wbs_m2s_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 303.320 400.000 303.920 ;
    END
  END io_wbs_m2s_data[23]
  PIN io_wbs_m2s_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END io_wbs_m2s_data[24]
  PIN io_wbs_m2s_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END io_wbs_m2s_data[25]
  PIN io_wbs_m2s_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 396.000 354.570 400.000 ;
    END
  END io_wbs_m2s_data[26]
  PIN io_wbs_m2s_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.120 4.000 361.720 ;
    END
  END io_wbs_m2s_data[27]
  PIN io_wbs_m2s_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 372.680 400.000 373.280 ;
    END
  END io_wbs_m2s_data[28]
  PIN io_wbs_m2s_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 396.000 372.510 400.000 ;
    END
  END io_wbs_m2s_data[29]
  PIN io_wbs_m2s_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END io_wbs_m2s_data[2]
  PIN io_wbs_m2s_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END io_wbs_m2s_data[30]
  PIN io_wbs_m2s_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 390.360 400.000 390.960 ;
    END
  END io_wbs_m2s_data[31]
  PIN io_wbs_m2s_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END io_wbs_m2s_data[3]
  PIN io_wbs_m2s_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 94.560 400.000 95.160 ;
    END
  END io_wbs_m2s_data[4]
  PIN io_wbs_m2s_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 396.000 99.730 400.000 ;
    END
  END io_wbs_m2s_data[5]
  PIN io_wbs_m2s_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END io_wbs_m2s_data[6]
  PIN io_wbs_m2s_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 396.000 136.070 400.000 ;
    END
  END io_wbs_m2s_data[7]
  PIN io_wbs_m2s_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 396.000 172.410 400.000 ;
    END
  END io_wbs_m2s_data[8]
  PIN io_wbs_m2s_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 164.600 400.000 165.200 ;
    END
  END io_wbs_m2s_data[9]
  PIN io_wbs_m2s_sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END io_wbs_m2s_sel[0]
  PIN io_wbs_m2s_sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 396.000 45.450 400.000 ;
    END
  END io_wbs_m2s_sel[1]
  PIN io_wbs_m2s_sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END io_wbs_m2s_sel[2]
  PIN io_wbs_m2s_sel[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 396.000 77.560 400.000 78.160 ;
    END
  END io_wbs_m2s_sel[3]
  PIN io_wbs_m2s_stb
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END io_wbs_m2s_stb
  PIN io_wbs_m2s_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END io_wbs_m2s_we
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 389.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 389.200 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 394.220 389.045 ;
      LAYER met1 ;
        RECT 5.520 9.900 394.220 389.200 ;
      LAYER met2 ;
        RECT 6.990 395.720 8.550 396.000 ;
        RECT 9.390 395.720 26.490 396.000 ;
        RECT 27.330 395.720 44.890 396.000 ;
        RECT 45.730 395.720 62.830 396.000 ;
        RECT 63.670 395.720 81.230 396.000 ;
        RECT 82.070 395.720 99.170 396.000 ;
        RECT 100.010 395.720 117.570 396.000 ;
        RECT 118.410 395.720 135.510 396.000 ;
        RECT 136.350 395.720 153.910 396.000 ;
        RECT 154.750 395.720 171.850 396.000 ;
        RECT 172.690 395.720 190.250 396.000 ;
        RECT 191.090 395.720 208.650 396.000 ;
        RECT 209.490 395.720 226.590 396.000 ;
        RECT 227.430 395.720 244.990 396.000 ;
        RECT 245.830 395.720 262.930 396.000 ;
        RECT 263.770 395.720 281.330 396.000 ;
        RECT 282.170 395.720 299.270 396.000 ;
        RECT 300.110 395.720 317.670 396.000 ;
        RECT 318.510 395.720 335.610 396.000 ;
        RECT 336.450 395.720 354.010 396.000 ;
        RECT 354.850 395.720 371.950 396.000 ;
        RECT 372.790 395.720 390.350 396.000 ;
        RECT 391.190 395.720 391.830 396.000 ;
        RECT 6.990 4.280 391.830 395.720 ;
        RECT 6.990 3.670 8.090 4.280 ;
        RECT 8.930 3.670 24.650 4.280 ;
        RECT 25.490 3.670 41.210 4.280 ;
        RECT 42.050 3.670 57.770 4.280 ;
        RECT 58.610 3.670 74.790 4.280 ;
        RECT 75.630 3.670 91.350 4.280 ;
        RECT 92.190 3.670 107.910 4.280 ;
        RECT 108.750 3.670 124.470 4.280 ;
        RECT 125.310 3.670 141.490 4.280 ;
        RECT 142.330 3.670 158.050 4.280 ;
        RECT 158.890 3.670 174.610 4.280 ;
        RECT 175.450 3.670 191.170 4.280 ;
        RECT 192.010 3.670 208.190 4.280 ;
        RECT 209.030 3.670 224.750 4.280 ;
        RECT 225.590 3.670 241.310 4.280 ;
        RECT 242.150 3.670 257.870 4.280 ;
        RECT 258.710 3.670 274.890 4.280 ;
        RECT 275.730 3.670 291.450 4.280 ;
        RECT 292.290 3.670 308.010 4.280 ;
        RECT 308.850 3.670 324.570 4.280 ;
        RECT 325.410 3.670 341.590 4.280 ;
        RECT 342.430 3.670 358.150 4.280 ;
        RECT 358.990 3.670 374.710 4.280 ;
        RECT 375.550 3.670 391.270 4.280 ;
      LAYER met3 ;
        RECT 4.400 391.360 396.000 392.185 ;
        RECT 4.400 391.320 395.600 391.360 ;
        RECT 4.000 389.960 395.600 391.320 ;
        RECT 4.000 377.080 396.000 389.960 ;
        RECT 4.400 375.680 396.000 377.080 ;
        RECT 4.000 373.680 396.000 375.680 ;
        RECT 4.000 372.280 395.600 373.680 ;
        RECT 4.000 362.120 396.000 372.280 ;
        RECT 4.400 360.720 396.000 362.120 ;
        RECT 4.000 356.680 396.000 360.720 ;
        RECT 4.000 355.280 395.600 356.680 ;
        RECT 4.000 346.480 396.000 355.280 ;
        RECT 4.400 345.080 396.000 346.480 ;
        RECT 4.000 339.000 396.000 345.080 ;
        RECT 4.000 337.600 395.600 339.000 ;
        RECT 4.000 330.840 396.000 337.600 ;
        RECT 4.400 329.440 396.000 330.840 ;
        RECT 4.000 322.000 396.000 329.440 ;
        RECT 4.000 320.600 395.600 322.000 ;
        RECT 4.000 315.880 396.000 320.600 ;
        RECT 4.400 314.480 396.000 315.880 ;
        RECT 4.000 304.320 396.000 314.480 ;
        RECT 4.000 302.920 395.600 304.320 ;
        RECT 4.000 300.240 396.000 302.920 ;
        RECT 4.400 298.840 396.000 300.240 ;
        RECT 4.000 287.320 396.000 298.840 ;
        RECT 4.000 285.920 395.600 287.320 ;
        RECT 4.000 285.280 396.000 285.920 ;
        RECT 4.400 283.880 396.000 285.280 ;
        RECT 4.000 269.640 396.000 283.880 ;
        RECT 4.400 268.240 395.600 269.640 ;
        RECT 4.000 254.000 396.000 268.240 ;
        RECT 4.400 252.600 396.000 254.000 ;
        RECT 4.000 251.960 396.000 252.600 ;
        RECT 4.000 250.560 395.600 251.960 ;
        RECT 4.000 239.040 396.000 250.560 ;
        RECT 4.400 237.640 396.000 239.040 ;
        RECT 4.000 234.960 396.000 237.640 ;
        RECT 4.000 233.560 395.600 234.960 ;
        RECT 4.000 223.400 396.000 233.560 ;
        RECT 4.400 222.000 396.000 223.400 ;
        RECT 4.000 217.280 396.000 222.000 ;
        RECT 4.000 215.880 395.600 217.280 ;
        RECT 4.000 208.440 396.000 215.880 ;
        RECT 4.400 207.040 396.000 208.440 ;
        RECT 4.000 200.280 396.000 207.040 ;
        RECT 4.000 198.880 395.600 200.280 ;
        RECT 4.000 192.800 396.000 198.880 ;
        RECT 4.400 191.400 396.000 192.800 ;
        RECT 4.000 182.600 396.000 191.400 ;
        RECT 4.000 181.200 395.600 182.600 ;
        RECT 4.000 177.160 396.000 181.200 ;
        RECT 4.400 175.760 396.000 177.160 ;
        RECT 4.000 165.600 396.000 175.760 ;
        RECT 4.000 164.200 395.600 165.600 ;
        RECT 4.000 162.200 396.000 164.200 ;
        RECT 4.400 160.800 396.000 162.200 ;
        RECT 4.000 147.920 396.000 160.800 ;
        RECT 4.000 146.560 395.600 147.920 ;
        RECT 4.400 146.520 395.600 146.560 ;
        RECT 4.400 145.160 396.000 146.520 ;
        RECT 4.000 130.920 396.000 145.160 ;
        RECT 4.400 130.240 396.000 130.920 ;
        RECT 4.400 129.520 395.600 130.240 ;
        RECT 4.000 128.840 395.600 129.520 ;
        RECT 4.000 115.960 396.000 128.840 ;
        RECT 4.400 114.560 396.000 115.960 ;
        RECT 4.000 113.240 396.000 114.560 ;
        RECT 4.000 111.840 395.600 113.240 ;
        RECT 4.000 100.320 396.000 111.840 ;
        RECT 4.400 98.920 396.000 100.320 ;
        RECT 4.000 95.560 396.000 98.920 ;
        RECT 4.000 94.160 395.600 95.560 ;
        RECT 4.000 85.360 396.000 94.160 ;
        RECT 4.400 83.960 396.000 85.360 ;
        RECT 4.000 78.560 396.000 83.960 ;
        RECT 4.000 77.160 395.600 78.560 ;
        RECT 4.000 69.720 396.000 77.160 ;
        RECT 4.400 68.320 396.000 69.720 ;
        RECT 4.000 60.880 396.000 68.320 ;
        RECT 4.000 59.480 395.600 60.880 ;
        RECT 4.000 54.080 396.000 59.480 ;
        RECT 4.400 52.680 396.000 54.080 ;
        RECT 4.000 43.880 396.000 52.680 ;
        RECT 4.000 42.480 395.600 43.880 ;
        RECT 4.000 39.120 396.000 42.480 ;
        RECT 4.400 37.720 396.000 39.120 ;
        RECT 4.000 26.200 396.000 37.720 ;
        RECT 4.000 24.800 395.600 26.200 ;
        RECT 4.000 23.480 396.000 24.800 ;
        RECT 4.400 22.080 396.000 23.480 ;
        RECT 4.000 9.200 396.000 22.080 ;
        RECT 4.000 8.520 395.600 9.200 ;
        RECT 4.400 7.800 395.600 8.520 ;
        RECT 4.400 7.655 396.000 7.800 ;
      LAYER met4 ;
        RECT 101.495 11.055 174.240 388.105 ;
        RECT 176.640 11.055 251.040 388.105 ;
        RECT 253.440 11.055 327.840 388.105 ;
        RECT 330.240 11.055 364.945 388.105 ;
  END
END Motor_Top
END LIBRARY

